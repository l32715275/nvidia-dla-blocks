module NV_NVDLA_BASIC_REG_single( // @[:@3.2]
  input         reset, // @[:@5.4]
  input         io_nvdla_core_clk, // @[:@6.4]
  output [31:0] io_reg_rd_data, // @[:@6.4]
  input  [11:0] io_reg_offset, // @[:@6.4]
  input  [31:0] io_reg_wr_data, // @[:@6.4]
  input         io_reg_wr_en, // @[:@6.4]
  output        io_producer, // @[:@6.4]
  input         io_consumer, // @[:@6.4]
  input  [1:0]  io_status_0, // @[:@6.4]
  input  [1:0]  io_status_1 // @[:@6.4]
);
  wire [31:0] _GEN_1; // @[NV_NVDLA_BASIC_REG_single.scala 46:43:@8.4]
  wire  _T_24; // @[NV_NVDLA_BASIC_REG_single.scala 46:43:@8.4]
  wire  _T_25; // @[NV_NVDLA_BASIC_REG_single.scala 46:66:@9.4]
  wire [31:0] _T_35; // @[Cat.scala 30:58:@14.4]
  wire [31:0] _T_41; // @[Cat.scala 30:58:@17.4]
  wire  _T_42; // @[Mux.scala 46:19:@18.4]
  wire [31:0] _T_43; // @[Mux.scala 46:16:@19.4]
  wire  _T_44; // @[Mux.scala 46:19:@20.4]
  wire  _T_46; // @[NV_NVDLA_BASIC_REG_single.scala 59:44:@23.4]
  reg  _T_49; // @[Reg.scala 19:20:@24.4]
  reg [31:0] _RAND_0;
  wire  _GEN_0; // @[Reg.scala 20:19:@25.4]
  assign _GEN_1 = {{20'd0}, io_reg_offset}; // @[NV_NVDLA_BASIC_REG_single.scala 46:43:@8.4]
  assign _T_24 = _GEN_1 == 32'h4; // @[NV_NVDLA_BASIC_REG_single.scala 46:43:@8.4]
  assign _T_25 = _T_24 & io_reg_wr_en; // @[NV_NVDLA_BASIC_REG_single.scala 46:66:@9.4]
  assign _T_35 = {15'h0,io_consumer,15'h0,io_producer}; // @[Cat.scala 30:58:@14.4]
  assign _T_41 = {14'h0,io_status_1,14'h0,io_status_0}; // @[Cat.scala 30:58:@17.4]
  assign _T_42 = 32'h0 == _GEN_1; // @[Mux.scala 46:19:@18.4]
  assign _T_43 = _T_42 ? _T_41 : 32'h0; // @[Mux.scala 46:16:@19.4]
  assign _T_44 = 32'h4 == _GEN_1; // @[Mux.scala 46:19:@20.4]
  assign _T_46 = io_reg_wr_data[0]; // @[NV_NVDLA_BASIC_REG_single.scala 59:44:@23.4]
  assign _GEN_0 = _T_25 ? _T_46 : _T_49; // @[Reg.scala 20:19:@25.4]
  assign io_reg_rd_data = _T_44 ? _T_35 : _T_43; // @[NV_NVDLA_BASIC_REG_single.scala 50:20:@22.4]
  assign io_producer = _T_49; // @[NV_NVDLA_BASIC_REG_single.scala 59:17:@28.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_49 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_49 <= 1'h0;
    end else begin
      if (_T_25) begin
        _T_49 <= _T_46;
      end
    end
  end
endmodule
module NV_NVDLA_CSC_dual_reg( // @[:@30.2]
  input         reset, // @[:@32.4]
  input         io_nvdla_core_clk, // @[:@33.4]
  output [31:0] io_reg_rd_data, // @[:@33.4]
  input  [11:0] io_reg_offset, // @[:@33.4]
  input  [31:0] io_reg_wr_data, // @[:@33.4]
  input         io_reg_wr_en, // @[:@33.4]
  output [20:0] io_field_atomics, // @[:@33.4]
  output [4:0]  io_field_data_bank, // @[:@33.4]
  output [4:0]  io_field_weight_bank, // @[:@33.4]
  output [4:0]  io_field_batches, // @[:@33.4]
  output [2:0]  io_field_conv_x_stride_ext, // @[:@33.4]
  output [2:0]  io_field_conv_y_stride_ext, // @[:@33.4]
  output [31:0] io_field_cya, // @[:@33.4]
  output        io_field_datain_format, // @[:@33.4]
  output [12:0] io_field_datain_height_ext, // @[:@33.4]
  output [12:0] io_field_datain_width_ext, // @[:@33.4]
  output [12:0] io_field_datain_channel_ext, // @[:@33.4]
  output [12:0] io_field_dataout_height, // @[:@33.4]
  output [12:0] io_field_dataout_width, // @[:@33.4]
  output [12:0] io_field_dataout_channel, // @[:@33.4]
  output [4:0]  io_field_x_dilation_ext, // @[:@33.4]
  output [4:0]  io_field_y_dilation_ext, // @[:@33.4]
  output [13:0] io_field_entries, // @[:@33.4]
  output        io_field_conv_mode, // @[:@33.4]
  output        io_field_data_reuse, // @[:@33.4]
  output [1:0]  io_field_in_precision, // @[:@33.4]
  output [1:0]  io_field_proc_precision, // @[:@33.4]
  output        io_field_skip_data_rls, // @[:@33.4]
  output        io_field_skip_weight_rls, // @[:@33.4]
  output        io_field_weight_reuse, // @[:@33.4]
  output [1:0]  io_field_y_extension, // @[:@33.4]
  output [1:0]  io_field_pra_truncate, // @[:@33.4]
  output [11:0] io_field_rls_slices, // @[:@33.4]
  output [31:0] io_field_weight_bytes, // @[:@33.4]
  output        io_field_weight_format, // @[:@33.4]
  output [4:0]  io_field_weight_height_ext, // @[:@33.4]
  output [4:0]  io_field_weight_width_ext, // @[:@33.4]
  output [12:0] io_field_weight_channel_ext, // @[:@33.4]
  output [12:0] io_field_weight_kernel, // @[:@33.4]
  output [27:0] io_field_wmb_bytes, // @[:@33.4]
  output [4:0]  io_field_pad_left, // @[:@33.4]
  output [4:0]  io_field_pad_top, // @[:@33.4]
  output [15:0] io_field_pad_value, // @[:@33.4]
  output        io_op_en_trigger, // @[:@33.4]
  input         io_op_en // @[:@33.4]
);
  wire [31:0] _GEN_37; // @[NV_NVDLA_CSC_dual_reg.scala 46:53:@35.4]
  wire  _T_94; // @[NV_NVDLA_CSC_dual_reg.scala 46:53:@35.4]
  wire  _T_95; // @[NV_NVDLA_CSC_dual_reg.scala 46:77:@36.4]
  wire  _T_97; // @[NV_NVDLA_CSC_dual_reg.scala 47:50:@37.4]
  wire  _T_98; // @[NV_NVDLA_CSC_dual_reg.scala 47:75:@38.4]
  wire  _T_100; // @[NV_NVDLA_CSC_dual_reg.scala 48:58:@39.4]
  wire  _T_101; // @[NV_NVDLA_CSC_dual_reg.scala 48:83:@40.4]
  wire  _T_103; // @[NV_NVDLA_CSC_dual_reg.scala 49:61:@41.4]
  wire  _T_104; // @[NV_NVDLA_CSC_dual_reg.scala 49:86:@42.4]
  wire  _T_106; // @[NV_NVDLA_CSC_dual_reg.scala 50:49:@43.4]
  wire  _T_107; // @[NV_NVDLA_CSC_dual_reg.scala 50:73:@44.4]
  wire  _T_109; // @[NV_NVDLA_CSC_dual_reg.scala 51:59:@45.4]
  wire  _T_110; // @[NV_NVDLA_CSC_dual_reg.scala 51:83:@46.4]
  wire  _T_112; // @[NV_NVDLA_CSC_dual_reg.scala 52:63:@47.4]
  wire  _T_113; // @[NV_NVDLA_CSC_dual_reg.scala 52:87:@48.4]
  wire  _T_115; // @[NV_NVDLA_CSC_dual_reg.scala 53:63:@49.4]
  wire  _T_116; // @[NV_NVDLA_CSC_dual_reg.scala 53:87:@50.4]
  wire  _T_118; // @[NV_NVDLA_CSC_dual_reg.scala 54:60:@51.4]
  wire  _T_119; // @[NV_NVDLA_CSC_dual_reg.scala 54:84:@52.4]
  wire  _T_121; // @[NV_NVDLA_CSC_dual_reg.scala 55:60:@53.4]
  wire  _T_122; // @[NV_NVDLA_CSC_dual_reg.scala 55:84:@54.4]
  wire  _T_124; // @[NV_NVDLA_CSC_dual_reg.scala 56:58:@55.4]
  wire  _T_125; // @[NV_NVDLA_CSC_dual_reg.scala 56:82:@56.4]
  wire  _T_127; // @[NV_NVDLA_CSC_dual_reg.scala 57:61:@57.4]
  wire  _T_128; // @[NV_NVDLA_CSC_dual_reg.scala 57:85:@58.4]
  wire  _T_130; // @[NV_NVDLA_CSC_dual_reg.scala 58:54:@59.4]
  wire  _T_131; // @[NV_NVDLA_CSC_dual_reg.scala 58:78:@60.4]
  wire  _T_133; // @[NV_NVDLA_CSC_dual_reg.scala 59:55:@61.4]
  wire  _T_136; // @[NV_NVDLA_CSC_dual_reg.scala 60:62:@63.4]
  wire  _T_137; // @[NV_NVDLA_CSC_dual_reg.scala 60:86:@64.4]
  wire  _T_139; // @[NV_NVDLA_CSC_dual_reg.scala 61:53:@65.4]
  wire  _T_140; // @[NV_NVDLA_CSC_dual_reg.scala 61:77:@66.4]
  wire  _T_142; // @[NV_NVDLA_CSC_dual_reg.scala 62:53:@67.4]
  wire  _T_143; // @[NV_NVDLA_CSC_dual_reg.scala 62:77:@68.4]
  wire  _T_145; // @[NV_NVDLA_CSC_dual_reg.scala 63:58:@69.4]
  wire  _T_146; // @[NV_NVDLA_CSC_dual_reg.scala 63:82:@70.4]
  wire  _T_148; // @[NV_NVDLA_CSC_dual_reg.scala 64:59:@71.4]
  wire  _T_149; // @[NV_NVDLA_CSC_dual_reg.scala 64:83:@72.4]
  wire  _T_151; // @[NV_NVDLA_CSC_dual_reg.scala 65:63:@73.4]
  wire  _T_152; // @[NV_NVDLA_CSC_dual_reg.scala 65:87:@74.4]
  wire  _T_154; // @[NV_NVDLA_CSC_dual_reg.scala 66:63:@75.4]
  wire  _T_155; // @[NV_NVDLA_CSC_dual_reg.scala 66:87:@76.4]
  wire  _T_157; // @[NV_NVDLA_CSC_dual_reg.scala 67:55:@77.4]
  wire  _T_158; // @[NV_NVDLA_CSC_dual_reg.scala 67:79:@78.4]
  wire  _T_160; // @[NV_NVDLA_CSC_dual_reg.scala 68:58:@79.4]
  wire  _T_161; // @[NV_NVDLA_CSC_dual_reg.scala 68:82:@80.4]
  wire  _T_163; // @[NV_NVDLA_CSC_dual_reg.scala 69:64:@81.4]
  wire  _T_164; // @[NV_NVDLA_CSC_dual_reg.scala 69:88:@82.4]
  wire [31:0] _T_168; // @[Cat.scala 30:58:@84.4]
  wire [31:0] _T_174; // @[Cat.scala 30:58:@87.4]
  wire [31:0] _T_177; // @[Cat.scala 30:58:@88.4]
  wire [31:0] _T_183; // @[Cat.scala 30:58:@91.4]
  wire [31:0] _T_187; // @[Cat.scala 30:58:@92.4]
  wire [31:0] _T_193; // @[Cat.scala 30:58:@95.4]
  wire [31:0] _T_196; // @[Cat.scala 30:58:@96.4]
  wire [31:0] _T_202; // @[Cat.scala 30:58:@99.4]
  wire [31:0] _T_205; // @[Cat.scala 30:58:@100.4]
  wire [31:0] _T_211; // @[Cat.scala 30:58:@103.4]
  wire [31:0] _T_214; // @[Cat.scala 30:58:@104.4]
  wire [16:0] _T_228; // @[Cat.scala 30:58:@110.4]
  wire [31:0] _T_235; // @[Cat.scala 30:58:@117.4]
  wire [31:0] _T_238; // @[Cat.scala 30:58:@118.4]
  wire [31:0] _T_241; // @[Cat.scala 30:58:@119.4]
  wire [31:0] _T_244; // @[Cat.scala 30:58:@120.4]
  wire [31:0] _T_247; // @[Cat.scala 30:58:@121.4]
  wire [31:0] _T_251; // @[Cat.scala 30:58:@122.4]
  wire [31:0] _T_257; // @[Cat.scala 30:58:@125.4]
  wire [31:0] _T_263; // @[Cat.scala 30:58:@128.4]
  wire [31:0] _T_266; // @[Cat.scala 30:58:@129.4]
  wire [31:0] _T_272; // @[Cat.scala 30:58:@132.4]
  wire [31:0] _T_275; // @[Cat.scala 30:58:@133.4]
  wire  _T_276; // @[Mux.scala 46:19:@134.4]
  wire [31:0] _T_277; // @[Mux.scala 46:16:@135.4]
  wire  _T_278; // @[Mux.scala 46:19:@136.4]
  wire [31:0] _T_279; // @[Mux.scala 46:16:@137.4]
  wire  _T_280; // @[Mux.scala 46:19:@138.4]
  wire [31:0] _T_281; // @[Mux.scala 46:16:@139.4]
  wire  _T_282; // @[Mux.scala 46:19:@140.4]
  wire [31:0] _T_283; // @[Mux.scala 46:16:@141.4]
  wire  _T_284; // @[Mux.scala 46:19:@142.4]
  wire [31:0] _T_285; // @[Mux.scala 46:16:@143.4]
  wire  _T_286; // @[Mux.scala 46:19:@144.4]
  wire [31:0] _T_287; // @[Mux.scala 46:16:@145.4]
  wire  _T_288; // @[Mux.scala 46:19:@146.4]
  wire [31:0] _T_289; // @[Mux.scala 46:16:@147.4]
  wire  _T_290; // @[Mux.scala 46:19:@148.4]
  wire [31:0] _T_291; // @[Mux.scala 46:16:@149.4]
  wire  _T_292; // @[Mux.scala 46:19:@150.4]
  wire [31:0] _T_293; // @[Mux.scala 46:16:@151.4]
  wire  _T_294; // @[Mux.scala 46:19:@152.4]
  wire [31:0] _T_295; // @[Mux.scala 46:16:@153.4]
  wire  _T_296; // @[Mux.scala 46:19:@154.4]
  wire [31:0] _T_297; // @[Mux.scala 46:16:@155.4]
  wire  _T_298; // @[Mux.scala 46:19:@156.4]
  wire [31:0] _T_299; // @[Mux.scala 46:16:@157.4]
  wire  _T_300; // @[Mux.scala 46:19:@158.4]
  wire [31:0] _T_301; // @[Mux.scala 46:16:@159.4]
  wire  _T_302; // @[Mux.scala 46:19:@160.4]
  wire [31:0] _T_303; // @[Mux.scala 46:16:@161.4]
  wire  _T_304; // @[Mux.scala 46:19:@162.4]
  wire [31:0] _T_305; // @[Mux.scala 46:16:@163.4]
  wire  _T_306; // @[Mux.scala 46:19:@164.4]
  wire [31:0] _T_307; // @[Mux.scala 46:16:@165.4]
  wire  _T_308; // @[Mux.scala 46:19:@166.4]
  wire [31:0] _T_309; // @[Mux.scala 46:16:@167.4]
  wire  _T_310; // @[Mux.scala 46:19:@168.4]
  wire [31:0] _T_311; // @[Mux.scala 46:16:@169.4]
  wire  _T_312; // @[Mux.scala 46:19:@170.4]
  wire [31:0] _T_313; // @[Mux.scala 46:16:@171.4]
  wire  _T_314; // @[Mux.scala 46:19:@172.4]
  wire [31:0] _T_315; // @[Mux.scala 46:16:@173.4]
  wire  _T_316; // @[Mux.scala 46:19:@174.4]
  wire [31:0] _T_317; // @[Mux.scala 46:16:@175.4]
  wire  _T_318; // @[Mux.scala 46:19:@176.4]
  wire [31:0] _T_319; // @[Mux.scala 46:16:@177.4]
  wire  _T_320; // @[Mux.scala 46:19:@178.4]
  wire [31:0] _T_321; // @[Mux.scala 46:16:@179.4]
  wire  _T_322; // @[Mux.scala 46:19:@180.4]
  wire [20:0] _T_324; // @[NV_NVDLA_CSC_dual_reg.scala 132:49:@183.4]
  reg [20:0] _T_327; // @[Reg.scala 19:20:@184.4]
  reg [31:0] _RAND_0;
  wire [20:0] _GEN_0; // @[Reg.scala 20:19:@185.4]
  wire [4:0] _T_328; // @[NV_NVDLA_CSC_dual_reg.scala 134:51:@189.4]
  reg [4:0] _T_331; // @[Reg.scala 19:20:@190.4]
  reg [31:0] _RAND_1;
  wire [4:0] _GEN_1; // @[Reg.scala 20:19:@191.4]
  wire [4:0] _T_332; // @[NV_NVDLA_CSC_dual_reg.scala 136:53:@195.4]
  reg [4:0] _T_335; // @[Reg.scala 19:20:@196.4]
  reg [31:0] _RAND_2;
  wire [4:0] _GEN_2; // @[Reg.scala 20:19:@197.4]
  reg [4:0] _T_339; // @[Reg.scala 19:20:@202.4]
  reg [31:0] _RAND_3;
  wire [4:0] _GEN_3; // @[Reg.scala 20:19:@203.4]
  wire [2:0] _T_340; // @[NV_NVDLA_CSC_dual_reg.scala 140:59:@207.4]
  reg [2:0] _T_343; // @[Reg.scala 19:20:@208.4]
  reg [31:0] _RAND_4;
  wire [2:0] _GEN_4; // @[Reg.scala 20:19:@209.4]
  wire [2:0] _T_344; // @[NV_NVDLA_CSC_dual_reg.scala 142:59:@213.4]
  reg [2:0] _T_347; // @[Reg.scala 19:20:@214.4]
  reg [31:0] _RAND_5;
  wire [2:0] _GEN_5; // @[Reg.scala 20:19:@215.4]
  reg [31:0] _T_350; // @[Reg.scala 19:20:@219.4]
  reg [31:0] _RAND_6;
  wire [31:0] _GEN_6; // @[Reg.scala 20:19:@220.4]
  wire  _T_351; // @[NV_NVDLA_CSC_dual_reg.scala 146:55:@224.4]
  reg  _T_354; // @[Reg.scala 19:20:@225.4]
  reg [31:0] _RAND_7;
  wire  _GEN_7; // @[Reg.scala 20:19:@226.4]
  wire [12:0] _T_355; // @[NV_NVDLA_CSC_dual_reg.scala 148:59:@230.4]
  reg [12:0] _T_358; // @[Reg.scala 19:20:@231.4]
  reg [31:0] _RAND_8;
  wire [12:0] _GEN_8; // @[Reg.scala 20:19:@232.4]
  wire [12:0] _T_359; // @[NV_NVDLA_CSC_dual_reg.scala 150:58:@236.4]
  reg [12:0] _T_362; // @[Reg.scala 19:20:@237.4]
  reg [31:0] _RAND_9;
  wire [12:0] _GEN_9; // @[Reg.scala 20:19:@238.4]
  reg [12:0] _T_366; // @[Reg.scala 19:20:@243.4]
  reg [31:0] _RAND_10;
  wire [12:0] _GEN_10; // @[Reg.scala 20:19:@244.4]
  reg [12:0] _T_370; // @[Reg.scala 19:20:@249.4]
  reg [31:0] _RAND_11;
  wire [12:0] _GEN_11; // @[Reg.scala 20:19:@250.4]
  reg [12:0] _T_374; // @[Reg.scala 19:20:@255.4]
  reg [31:0] _RAND_12;
  wire [12:0] _GEN_12; // @[Reg.scala 20:19:@256.4]
  reg [12:0] _T_378; // @[Reg.scala 19:20:@261.4]
  reg [31:0] _RAND_13;
  wire [12:0] _GEN_13; // @[Reg.scala 20:19:@262.4]
  reg [4:0] _T_382; // @[Reg.scala 19:20:@267.4]
  reg [31:0] _RAND_14;
  wire [4:0] _GEN_14; // @[Reg.scala 20:19:@268.4]
  reg [4:0] _T_386; // @[Reg.scala 19:20:@273.4]
  reg [31:0] _RAND_15;
  wire [4:0] _GEN_15; // @[Reg.scala 20:19:@274.4]
  wire [13:0] _T_387; // @[NV_NVDLA_CSC_dual_reg.scala 164:49:@278.4]
  reg [13:0] _T_390; // @[Reg.scala 19:20:@279.4]
  reg [31:0] _RAND_16;
  wire [13:0] _GEN_16; // @[Reg.scala 20:19:@280.4]
  reg  _T_394; // @[Reg.scala 19:20:@285.4]
  reg [31:0] _RAND_17;
  wire  _GEN_17; // @[Reg.scala 20:19:@286.4]
  wire  _T_395; // @[NV_NVDLA_CSC_dual_reg.scala 168:52:@290.4]
  reg  _T_398; // @[Reg.scala 19:20:@291.4]
  reg [31:0] _RAND_18;
  wire  _GEN_18; // @[Reg.scala 20:19:@292.4]
  wire [1:0] _T_399; // @[NV_NVDLA_CSC_dual_reg.scala 170:54:@296.4]
  reg [1:0] _T_402; // @[Reg.scala 19:20:@297.4]
  reg [31:0] _RAND_19;
  wire [1:0] _GEN_19; // @[Reg.scala 20:19:@298.4]
  wire [1:0] _T_403; // @[NV_NVDLA_CSC_dual_reg.scala 172:56:@302.4]
  reg [1:0] _T_406; // @[Reg.scala 19:20:@303.4]
  reg [31:0] _RAND_20;
  wire [1:0] _GEN_20; // @[Reg.scala 20:19:@304.4]
  wire  _T_407; // @[NV_NVDLA_CSC_dual_reg.scala 174:55:@308.4]
  reg  _T_410; // @[Reg.scala 19:20:@309.4]
  reg [31:0] _RAND_21;
  wire  _GEN_21; // @[Reg.scala 20:19:@310.4]
  wire  _T_411; // @[NV_NVDLA_CSC_dual_reg.scala 176:57:@314.4]
  reg  _T_414; // @[Reg.scala 19:20:@315.4]
  reg [31:0] _RAND_22;
  wire  _GEN_22; // @[Reg.scala 20:19:@316.4]
  wire  _T_415; // @[NV_NVDLA_CSC_dual_reg.scala 178:54:@320.4]
  reg  _T_418; // @[Reg.scala 19:20:@321.4]
  reg [31:0] _RAND_23;
  wire  _GEN_23; // @[Reg.scala 20:19:@322.4]
  wire [1:0] _T_419; // @[NV_NVDLA_CSC_dual_reg.scala 180:53:@326.4]
  reg [1:0] _T_422; // @[Reg.scala 19:20:@327.4]
  reg [31:0] _RAND_24;
  wire [1:0] _GEN_24; // @[Reg.scala 20:19:@328.4]
  reg [1:0] _T_426; // @[Reg.scala 19:20:@333.4]
  reg [31:0] _RAND_25;
  wire [1:0] _GEN_25; // @[Reg.scala 20:19:@334.4]
  wire [11:0] _T_427; // @[NV_NVDLA_CSC_dual_reg.scala 184:52:@338.4]
  reg [11:0] _T_430; // @[Reg.scala 19:20:@339.4]
  reg [31:0] _RAND_26;
  wire [11:0] _GEN_26; // @[Reg.scala 20:19:@340.4]
  reg [31:0] _T_434; // @[Reg.scala 19:20:@345.4]
  reg [31:0] _RAND_27;
  wire [31:0] _GEN_27; // @[Reg.scala 20:19:@346.4]
  reg  _T_438; // @[Reg.scala 19:20:@351.4]
  reg [31:0] _RAND_28;
  wire  _GEN_28; // @[Reg.scala 20:19:@352.4]
  reg [4:0] _T_442; // @[Reg.scala 19:20:@357.4]
  reg [31:0] _RAND_29;
  wire [4:0] _GEN_29; // @[Reg.scala 20:19:@358.4]
  reg [4:0] _T_446; // @[Reg.scala 19:20:@363.4]
  reg [31:0] _RAND_30;
  wire [4:0] _GEN_30; // @[Reg.scala 20:19:@364.4]
  reg [12:0] _T_450; // @[Reg.scala 19:20:@369.4]
  reg [31:0] _RAND_31;
  wire [12:0] _GEN_31; // @[Reg.scala 20:19:@370.4]
  reg [12:0] _T_454; // @[Reg.scala 19:20:@375.4]
  reg [31:0] _RAND_32;
  wire [12:0] _GEN_32; // @[Reg.scala 20:19:@376.4]
  wire [27:0] _T_455; // @[NV_NVDLA_CSC_dual_reg.scala 198:51:@380.4]
  reg [27:0] _T_458; // @[Reg.scala 19:20:@381.4]
  reg [31:0] _RAND_33;
  wire [27:0] _GEN_33; // @[Reg.scala 20:19:@382.4]
  reg [4:0] _T_462; // @[Reg.scala 19:20:@387.4]
  reg [31:0] _RAND_34;
  wire [4:0] _GEN_34; // @[Reg.scala 20:19:@388.4]
  reg [4:0] _T_466; // @[Reg.scala 19:20:@393.4]
  reg [31:0] _RAND_35;
  wire [4:0] _GEN_35; // @[Reg.scala 20:19:@394.4]
  wire [15:0] _T_467; // @[NV_NVDLA_CSC_dual_reg.scala 204:51:@398.4]
  reg [15:0] _T_470; // @[Reg.scala 19:20:@399.4]
  reg [31:0] _RAND_36;
  wire [15:0] _GEN_36; // @[Reg.scala 20:19:@400.4]
  assign _GEN_37 = {{20'd0}, io_reg_offset}; // @[NV_NVDLA_CSC_dual_reg.scala 46:53:@35.4]
  assign _T_94 = _GEN_37 == 32'h44; // @[NV_NVDLA_CSC_dual_reg.scala 46:53:@35.4]
  assign _T_95 = _T_94 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 46:77:@36.4]
  assign _T_97 = _GEN_37 == 32'h5c; // @[NV_NVDLA_CSC_dual_reg.scala 47:50:@37.4]
  assign _T_98 = _T_97 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 47:75:@38.4]
  assign _T_100 = _GEN_37 == 32'h1c; // @[NV_NVDLA_CSC_dual_reg.scala 48:58:@39.4]
  assign _T_101 = _T_100 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 48:83:@40.4]
  assign _T_103 = _GEN_37 == 32'h4c; // @[NV_NVDLA_CSC_dual_reg.scala 49:61:@41.4]
  assign _T_104 = _T_103 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 49:86:@42.4]
  assign _T_106 = _GEN_37 == 32'h64; // @[NV_NVDLA_CSC_dual_reg.scala 50:49:@43.4]
  assign _T_107 = _T_106 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 50:73:@44.4]
  assign _T_109 = _GEN_37 == 32'h10; // @[NV_NVDLA_CSC_dual_reg.scala 51:59:@45.4]
  assign _T_110 = _T_109 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 51:83:@46.4]
  assign _T_112 = _GEN_37 == 32'h14; // @[NV_NVDLA_CSC_dual_reg.scala 52:63:@47.4]
  assign _T_113 = _T_112 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 52:87:@48.4]
  assign _T_115 = _GEN_37 == 32'h18; // @[NV_NVDLA_CSC_dual_reg.scala 53:63:@49.4]
  assign _T_116 = _T_115 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 53:87:@50.4]
  assign _T_118 = _GEN_37 == 32'h3c; // @[NV_NVDLA_CSC_dual_reg.scala 54:60:@51.4]
  assign _T_119 = _T_118 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 54:84:@52.4]
  assign _T_121 = _GEN_37 == 32'h40; // @[NV_NVDLA_CSC_dual_reg.scala 55:60:@53.4]
  assign _T_122 = _T_121 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 55:84:@54.4]
  assign _T_124 = _GEN_37 == 32'h50; // @[NV_NVDLA_CSC_dual_reg.scala 56:58:@55.4]
  assign _T_125 = _T_124 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 56:82:@56.4]
  assign _T_127 = _GEN_37 == 32'h24; // @[NV_NVDLA_CSC_dual_reg.scala 57:61:@57.4]
  assign _T_128 = _T_127 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 57:85:@58.4]
  assign _T_130 = _GEN_37 == 32'hc; // @[NV_NVDLA_CSC_dual_reg.scala 58:54:@59.4]
  assign _T_131 = _T_130 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 58:78:@60.4]
  assign _T_133 = _GEN_37 == 32'h8; // @[NV_NVDLA_CSC_dual_reg.scala 59:55:@61.4]
  assign _T_136 = _GEN_37 == 32'h20; // @[NV_NVDLA_CSC_dual_reg.scala 60:62:@63.4]
  assign _T_137 = _T_136 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 60:86:@64.4]
  assign _T_139 = _GEN_37 == 32'h60; // @[NV_NVDLA_CSC_dual_reg.scala 61:53:@65.4]
  assign _T_140 = _T_139 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 61:77:@66.4]
  assign _T_142 = _GEN_37 == 32'h48; // @[NV_NVDLA_CSC_dual_reg.scala 62:53:@67.4]
  assign _T_143 = _T_142 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 62:77:@68.4]
  assign _T_145 = _GEN_37 == 32'h34; // @[NV_NVDLA_CSC_dual_reg.scala 63:58:@69.4]
  assign _T_146 = _T_145 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 63:82:@70.4]
  assign _T_148 = _GEN_37 == 32'h28; // @[NV_NVDLA_CSC_dual_reg.scala 64:59:@71.4]
  assign _T_149 = _T_148 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 64:83:@72.4]
  assign _T_151 = _GEN_37 == 32'h2c; // @[NV_NVDLA_CSC_dual_reg.scala 65:63:@73.4]
  assign _T_152 = _T_151 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 65:87:@74.4]
  assign _T_154 = _GEN_37 == 32'h30; // @[NV_NVDLA_CSC_dual_reg.scala 66:63:@75.4]
  assign _T_155 = _T_154 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 66:87:@76.4]
  assign _T_157 = _GEN_37 == 32'h38; // @[NV_NVDLA_CSC_dual_reg.scala 67:55:@77.4]
  assign _T_158 = _T_157 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 67:79:@78.4]
  assign _T_160 = _GEN_37 == 32'h54; // @[NV_NVDLA_CSC_dual_reg.scala 68:58:@79.4]
  assign _T_161 = _T_160 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 68:82:@80.4]
  assign _T_163 = _GEN_37 == 32'h58; // @[NV_NVDLA_CSC_dual_reg.scala 69:64:@81.4]
  assign _T_164 = _T_163 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 69:88:@82.4]
  assign _T_168 = {11'h0,io_field_atomics}; // @[Cat.scala 30:58:@84.4]
  assign _T_174 = {11'h0,io_field_weight_bank,11'h0,io_field_data_bank}; // @[Cat.scala 30:58:@87.4]
  assign _T_177 = {27'h0,io_field_batches}; // @[Cat.scala 30:58:@88.4]
  assign _T_183 = {13'h0,io_field_conv_y_stride_ext,13'h0,io_field_conv_x_stride_ext}; // @[Cat.scala 30:58:@91.4]
  assign _T_187 = {31'h0,io_field_datain_format}; // @[Cat.scala 30:58:@92.4]
  assign _T_193 = {3'h0,io_field_datain_height_ext,3'h0,io_field_datain_width_ext}; // @[Cat.scala 30:58:@95.4]
  assign _T_196 = {19'h0,io_field_datain_channel_ext}; // @[Cat.scala 30:58:@96.4]
  assign _T_202 = {3'h0,io_field_dataout_height,3'h0,io_field_dataout_width}; // @[Cat.scala 30:58:@99.4]
  assign _T_205 = {19'h0,io_field_dataout_channel}; // @[Cat.scala 30:58:@100.4]
  assign _T_211 = {11'h0,io_field_y_dilation_ext,11'h0,io_field_x_dilation_ext}; // @[Cat.scala 30:58:@103.4]
  assign _T_214 = {18'h0,io_field_entries}; // @[Cat.scala 30:58:@104.4]
  assign _T_228 = {io_field_data_reuse,2'h0,io_field_proc_precision,2'h0,io_field_in_precision,7'h0,io_field_conv_mode}; // @[Cat.scala 30:58:@110.4]
  assign _T_235 = {3'h0,io_field_skip_weight_rls,3'h0,io_field_skip_data_rls,3'h0,io_field_weight_reuse,3'h0,_T_228}; // @[Cat.scala 30:58:@117.4]
  assign _T_238 = {31'h0,io_op_en}; // @[Cat.scala 30:58:@118.4]
  assign _T_241 = {30'h0,io_field_y_extension}; // @[Cat.scala 30:58:@119.4]
  assign _T_244 = {30'h0,io_field_pra_truncate}; // @[Cat.scala 30:58:@120.4]
  assign _T_247 = {20'h0,io_field_rls_slices}; // @[Cat.scala 30:58:@121.4]
  assign _T_251 = {31'h0,io_field_weight_format}; // @[Cat.scala 30:58:@122.4]
  assign _T_257 = {11'h0,io_field_weight_height_ext,11'h0,io_field_weight_width_ext}; // @[Cat.scala 30:58:@125.4]
  assign _T_263 = {3'h0,io_field_weight_kernel,3'h0,io_field_weight_channel_ext}; // @[Cat.scala 30:58:@128.4]
  assign _T_266 = {4'h0,io_field_wmb_bytes}; // @[Cat.scala 30:58:@129.4]
  assign _T_272 = {11'h0,io_field_pad_top,11'h0,io_field_pad_left}; // @[Cat.scala 30:58:@132.4]
  assign _T_275 = {16'h0,io_field_pad_value}; // @[Cat.scala 30:58:@133.4]
  assign _T_276 = 32'h58 == _GEN_37; // @[Mux.scala 46:19:@134.4]
  assign _T_277 = _T_276 ? _T_275 : 32'h0; // @[Mux.scala 46:16:@135.4]
  assign _T_278 = 32'h54 == _GEN_37; // @[Mux.scala 46:19:@136.4]
  assign _T_279 = _T_278 ? _T_272 : _T_277; // @[Mux.scala 46:16:@137.4]
  assign _T_280 = 32'h38 == _GEN_37; // @[Mux.scala 46:19:@138.4]
  assign _T_281 = _T_280 ? _T_266 : _T_279; // @[Mux.scala 46:16:@139.4]
  assign _T_282 = 32'h30 == _GEN_37; // @[Mux.scala 46:19:@140.4]
  assign _T_283 = _T_282 ? _T_263 : _T_281; // @[Mux.scala 46:16:@141.4]
  assign _T_284 = 32'h2c == _GEN_37; // @[Mux.scala 46:19:@142.4]
  assign _T_285 = _T_284 ? _T_257 : _T_283; // @[Mux.scala 46:16:@143.4]
  assign _T_286 = 32'h28 == _GEN_37; // @[Mux.scala 46:19:@144.4]
  assign _T_287 = _T_286 ? _T_251 : _T_285; // @[Mux.scala 46:16:@145.4]
  assign _T_288 = 32'h34 == _GEN_37; // @[Mux.scala 46:19:@146.4]
  assign _T_289 = _T_288 ? io_field_weight_bytes : _T_287; // @[Mux.scala 46:16:@147.4]
  assign _T_290 = 32'h48 == _GEN_37; // @[Mux.scala 46:19:@148.4]
  assign _T_291 = _T_290 ? _T_247 : _T_289; // @[Mux.scala 46:16:@149.4]
  assign _T_292 = 32'h60 == _GEN_37; // @[Mux.scala 46:19:@150.4]
  assign _T_293 = _T_292 ? _T_244 : _T_291; // @[Mux.scala 46:16:@151.4]
  assign _T_294 = 32'h20 == _GEN_37; // @[Mux.scala 46:19:@152.4]
  assign _T_295 = _T_294 ? _T_241 : _T_293; // @[Mux.scala 46:16:@153.4]
  assign _T_296 = 32'h8 == _GEN_37; // @[Mux.scala 46:19:@154.4]
  assign _T_297 = _T_296 ? _T_238 : _T_295; // @[Mux.scala 46:16:@155.4]
  assign _T_298 = 32'hc == _GEN_37; // @[Mux.scala 46:19:@156.4]
  assign _T_299 = _T_298 ? _T_235 : _T_297; // @[Mux.scala 46:16:@157.4]
  assign _T_300 = 32'h24 == _GEN_37; // @[Mux.scala 46:19:@158.4]
  assign _T_301 = _T_300 ? _T_214 : _T_299; // @[Mux.scala 46:16:@159.4]
  assign _T_302 = 32'h50 == _GEN_37; // @[Mux.scala 46:19:@160.4]
  assign _T_303 = _T_302 ? _T_211 : _T_301; // @[Mux.scala 46:16:@161.4]
  assign _T_304 = 32'h40 == _GEN_37; // @[Mux.scala 46:19:@162.4]
  assign _T_305 = _T_304 ? _T_205 : _T_303; // @[Mux.scala 46:16:@163.4]
  assign _T_306 = 32'h3c == _GEN_37; // @[Mux.scala 46:19:@164.4]
  assign _T_307 = _T_306 ? _T_202 : _T_305; // @[Mux.scala 46:16:@165.4]
  assign _T_308 = 32'h18 == _GEN_37; // @[Mux.scala 46:19:@166.4]
  assign _T_309 = _T_308 ? _T_196 : _T_307; // @[Mux.scala 46:16:@167.4]
  assign _T_310 = 32'h14 == _GEN_37; // @[Mux.scala 46:19:@168.4]
  assign _T_311 = _T_310 ? _T_193 : _T_309; // @[Mux.scala 46:16:@169.4]
  assign _T_312 = 32'h10 == _GEN_37; // @[Mux.scala 46:19:@170.4]
  assign _T_313 = _T_312 ? _T_187 : _T_311; // @[Mux.scala 46:16:@171.4]
  assign _T_314 = 32'h64 == _GEN_37; // @[Mux.scala 46:19:@172.4]
  assign _T_315 = _T_314 ? io_field_cya : _T_313; // @[Mux.scala 46:16:@173.4]
  assign _T_316 = 32'h4c == _GEN_37; // @[Mux.scala 46:19:@174.4]
  assign _T_317 = _T_316 ? _T_183 : _T_315; // @[Mux.scala 46:16:@175.4]
  assign _T_318 = 32'h1c == _GEN_37; // @[Mux.scala 46:19:@176.4]
  assign _T_319 = _T_318 ? _T_177 : _T_317; // @[Mux.scala 46:16:@177.4]
  assign _T_320 = 32'h5c == _GEN_37; // @[Mux.scala 46:19:@178.4]
  assign _T_321 = _T_320 ? _T_174 : _T_319; // @[Mux.scala 46:16:@179.4]
  assign _T_322 = 32'h44 == _GEN_37; // @[Mux.scala 46:19:@180.4]
  assign _T_324 = io_reg_wr_data[20:0]; // @[NV_NVDLA_CSC_dual_reg.scala 132:49:@183.4]
  assign _GEN_0 = _T_95 ? _T_324 : _T_327; // @[Reg.scala 20:19:@185.4]
  assign _T_328 = io_reg_wr_data[4:0]; // @[NV_NVDLA_CSC_dual_reg.scala 134:51:@189.4]
  assign _GEN_1 = _T_98 ? _T_328 : _T_331; // @[Reg.scala 20:19:@191.4]
  assign _T_332 = io_reg_wr_data[20:16]; // @[NV_NVDLA_CSC_dual_reg.scala 136:53:@195.4]
  assign _GEN_2 = _T_98 ? _T_332 : _T_335; // @[Reg.scala 20:19:@197.4]
  assign _GEN_3 = _T_101 ? _T_328 : _T_339; // @[Reg.scala 20:19:@203.4]
  assign _T_340 = io_reg_wr_data[2:0]; // @[NV_NVDLA_CSC_dual_reg.scala 140:59:@207.4]
  assign _GEN_4 = _T_104 ? _T_340 : _T_343; // @[Reg.scala 20:19:@209.4]
  assign _T_344 = io_reg_wr_data[18:16]; // @[NV_NVDLA_CSC_dual_reg.scala 142:59:@213.4]
  assign _GEN_5 = _T_104 ? _T_344 : _T_347; // @[Reg.scala 20:19:@215.4]
  assign _GEN_6 = _T_107 ? io_reg_wr_data : _T_350; // @[Reg.scala 20:19:@220.4]
  assign _T_351 = io_reg_wr_data[0]; // @[NV_NVDLA_CSC_dual_reg.scala 146:55:@224.4]
  assign _GEN_7 = _T_110 ? _T_351 : _T_354; // @[Reg.scala 20:19:@226.4]
  assign _T_355 = io_reg_wr_data[28:16]; // @[NV_NVDLA_CSC_dual_reg.scala 148:59:@230.4]
  assign _GEN_8 = _T_113 ? _T_355 : _T_358; // @[Reg.scala 20:19:@232.4]
  assign _T_359 = io_reg_wr_data[12:0]; // @[NV_NVDLA_CSC_dual_reg.scala 150:58:@236.4]
  assign _GEN_9 = _T_113 ? _T_359 : _T_362; // @[Reg.scala 20:19:@238.4]
  assign _GEN_10 = _T_116 ? _T_359 : _T_366; // @[Reg.scala 20:19:@244.4]
  assign _GEN_11 = _T_119 ? _T_355 : _T_370; // @[Reg.scala 20:19:@250.4]
  assign _GEN_12 = _T_119 ? _T_359 : _T_374; // @[Reg.scala 20:19:@256.4]
  assign _GEN_13 = _T_122 ? _T_359 : _T_378; // @[Reg.scala 20:19:@262.4]
  assign _GEN_14 = _T_125 ? _T_328 : _T_382; // @[Reg.scala 20:19:@268.4]
  assign _GEN_15 = _T_125 ? _T_332 : _T_386; // @[Reg.scala 20:19:@274.4]
  assign _T_387 = io_reg_wr_data[13:0]; // @[NV_NVDLA_CSC_dual_reg.scala 164:49:@278.4]
  assign _GEN_16 = _T_128 ? _T_387 : _T_390; // @[Reg.scala 20:19:@280.4]
  assign _GEN_17 = _T_131 ? _T_351 : _T_394; // @[Reg.scala 20:19:@286.4]
  assign _T_395 = io_reg_wr_data[16]; // @[NV_NVDLA_CSC_dual_reg.scala 168:52:@290.4]
  assign _GEN_18 = _T_131 ? _T_395 : _T_398; // @[Reg.scala 20:19:@292.4]
  assign _T_399 = io_reg_wr_data[9:8]; // @[NV_NVDLA_CSC_dual_reg.scala 170:54:@296.4]
  assign _GEN_19 = _T_131 ? _T_399 : _T_402; // @[Reg.scala 20:19:@298.4]
  assign _T_403 = io_reg_wr_data[13:12]; // @[NV_NVDLA_CSC_dual_reg.scala 172:56:@302.4]
  assign _GEN_20 = _T_131 ? _T_403 : _T_406; // @[Reg.scala 20:19:@304.4]
  assign _T_407 = io_reg_wr_data[24]; // @[NV_NVDLA_CSC_dual_reg.scala 174:55:@308.4]
  assign _GEN_21 = _T_131 ? _T_407 : _T_410; // @[Reg.scala 20:19:@310.4]
  assign _T_411 = io_reg_wr_data[28]; // @[NV_NVDLA_CSC_dual_reg.scala 176:57:@314.4]
  assign _GEN_22 = _T_131 ? _T_411 : _T_414; // @[Reg.scala 20:19:@316.4]
  assign _T_415 = io_reg_wr_data[20]; // @[NV_NVDLA_CSC_dual_reg.scala 178:54:@320.4]
  assign _GEN_23 = _T_131 ? _T_415 : _T_418; // @[Reg.scala 20:19:@322.4]
  assign _T_419 = io_reg_wr_data[1:0]; // @[NV_NVDLA_CSC_dual_reg.scala 180:53:@326.4]
  assign _GEN_24 = _T_137 ? _T_419 : _T_422; // @[Reg.scala 20:19:@328.4]
  assign _GEN_25 = _T_140 ? _T_419 : _T_426; // @[Reg.scala 20:19:@334.4]
  assign _T_427 = io_reg_wr_data[11:0]; // @[NV_NVDLA_CSC_dual_reg.scala 184:52:@338.4]
  assign _GEN_26 = _T_143 ? _T_427 : _T_430; // @[Reg.scala 20:19:@340.4]
  assign _GEN_27 = _T_146 ? io_reg_wr_data : _T_434; // @[Reg.scala 20:19:@346.4]
  assign _GEN_28 = _T_149 ? _T_351 : _T_438; // @[Reg.scala 20:19:@352.4]
  assign _GEN_29 = _T_152 ? _T_332 : _T_442; // @[Reg.scala 20:19:@358.4]
  assign _GEN_30 = _T_152 ? _T_328 : _T_446; // @[Reg.scala 20:19:@364.4]
  assign _GEN_31 = _T_155 ? _T_359 : _T_450; // @[Reg.scala 20:19:@370.4]
  assign _GEN_32 = _T_155 ? _T_355 : _T_454; // @[Reg.scala 20:19:@376.4]
  assign _T_455 = io_reg_wr_data[27:0]; // @[NV_NVDLA_CSC_dual_reg.scala 198:51:@380.4]
  assign _GEN_33 = _T_158 ? _T_455 : _T_458; // @[Reg.scala 20:19:@382.4]
  assign _GEN_34 = _T_161 ? _T_328 : _T_462; // @[Reg.scala 20:19:@388.4]
  assign _GEN_35 = _T_161 ? _T_332 : _T_466; // @[Reg.scala 20:19:@394.4]
  assign _T_467 = io_reg_wr_data[15:0]; // @[NV_NVDLA_CSC_dual_reg.scala 204:51:@398.4]
  assign _GEN_36 = _T_164 ? _T_467 : _T_470; // @[Reg.scala 20:19:@400.4]
  assign io_reg_rd_data = _T_322 ? _T_168 : _T_321; // @[NV_NVDLA_CSC_dual_reg.scala 75:20:@182.4]
  assign io_field_atomics = _T_327; // @[NV_NVDLA_CSC_dual_reg.scala 132:22:@188.4]
  assign io_field_data_bank = _T_331; // @[NV_NVDLA_CSC_dual_reg.scala 134:24:@194.4]
  assign io_field_weight_bank = _T_335; // @[NV_NVDLA_CSC_dual_reg.scala 136:26:@200.4]
  assign io_field_batches = _T_339; // @[NV_NVDLA_CSC_dual_reg.scala 138:22:@206.4]
  assign io_field_conv_x_stride_ext = _T_343; // @[NV_NVDLA_CSC_dual_reg.scala 140:32:@212.4]
  assign io_field_conv_y_stride_ext = _T_347; // @[NV_NVDLA_CSC_dual_reg.scala 142:32:@218.4]
  assign io_field_cya = _T_350; // @[NV_NVDLA_CSC_dual_reg.scala 144:18:@223.4]
  assign io_field_datain_format = _T_354; // @[NV_NVDLA_CSC_dual_reg.scala 146:28:@229.4]
  assign io_field_datain_height_ext = _T_358; // @[NV_NVDLA_CSC_dual_reg.scala 148:32:@235.4]
  assign io_field_datain_width_ext = _T_362; // @[NV_NVDLA_CSC_dual_reg.scala 150:31:@241.4]
  assign io_field_datain_channel_ext = _T_366; // @[NV_NVDLA_CSC_dual_reg.scala 152:33:@247.4]
  assign io_field_dataout_height = _T_370; // @[NV_NVDLA_CSC_dual_reg.scala 154:29:@253.4]
  assign io_field_dataout_width = _T_374; // @[NV_NVDLA_CSC_dual_reg.scala 156:28:@259.4]
  assign io_field_dataout_channel = _T_378; // @[NV_NVDLA_CSC_dual_reg.scala 158:30:@265.4]
  assign io_field_x_dilation_ext = _T_382; // @[NV_NVDLA_CSC_dual_reg.scala 160:29:@271.4]
  assign io_field_y_dilation_ext = _T_386; // @[NV_NVDLA_CSC_dual_reg.scala 162:29:@277.4]
  assign io_field_entries = _T_390; // @[NV_NVDLA_CSC_dual_reg.scala 164:22:@283.4]
  assign io_field_conv_mode = _T_394; // @[NV_NVDLA_CSC_dual_reg.scala 166:24:@289.4]
  assign io_field_data_reuse = _T_398; // @[NV_NVDLA_CSC_dual_reg.scala 168:25:@295.4]
  assign io_field_in_precision = _T_402; // @[NV_NVDLA_CSC_dual_reg.scala 170:27:@301.4]
  assign io_field_proc_precision = _T_406; // @[NV_NVDLA_CSC_dual_reg.scala 172:29:@307.4]
  assign io_field_skip_data_rls = _T_410; // @[NV_NVDLA_CSC_dual_reg.scala 174:28:@313.4]
  assign io_field_skip_weight_rls = _T_414; // @[NV_NVDLA_CSC_dual_reg.scala 176:30:@319.4]
  assign io_field_weight_reuse = _T_418; // @[NV_NVDLA_CSC_dual_reg.scala 178:27:@325.4]
  assign io_field_y_extension = _T_422; // @[NV_NVDLA_CSC_dual_reg.scala 180:26:@331.4]
  assign io_field_pra_truncate = _T_426; // @[NV_NVDLA_CSC_dual_reg.scala 182:27:@337.4]
  assign io_field_rls_slices = _T_430; // @[NV_NVDLA_CSC_dual_reg.scala 184:25:@343.4]
  assign io_field_weight_bytes = _T_434; // @[NV_NVDLA_CSC_dual_reg.scala 186:27:@349.4]
  assign io_field_weight_format = _T_438; // @[NV_NVDLA_CSC_dual_reg.scala 188:28:@355.4]
  assign io_field_weight_height_ext = _T_442; // @[NV_NVDLA_CSC_dual_reg.scala 190:32:@361.4]
  assign io_field_weight_width_ext = _T_446; // @[NV_NVDLA_CSC_dual_reg.scala 192:31:@367.4]
  assign io_field_weight_channel_ext = _T_450; // @[NV_NVDLA_CSC_dual_reg.scala 194:33:@373.4]
  assign io_field_weight_kernel = _T_454; // @[NV_NVDLA_CSC_dual_reg.scala 196:28:@379.4]
  assign io_field_wmb_bytes = _T_458; // @[NV_NVDLA_CSC_dual_reg.scala 198:24:@385.4]
  assign io_field_pad_left = _T_462; // @[NV_NVDLA_CSC_dual_reg.scala 200:23:@391.4]
  assign io_field_pad_top = _T_466; // @[NV_NVDLA_CSC_dual_reg.scala 202:22:@397.4]
  assign io_field_pad_value = _T_470; // @[NV_NVDLA_CSC_dual_reg.scala 204:24:@403.4]
  assign io_op_en_trigger = _T_133 & io_reg_wr_en; // @[NV_NVDLA_CSC_dual_reg.scala 71:22:@83.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_327 = _RAND_0[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_331 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_335 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_339 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_343 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_347 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_350 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_354 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_358 = _RAND_8[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_362 = _RAND_9[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_366 = _RAND_10[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_370 = _RAND_11[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_374 = _RAND_12[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_378 = _RAND_13[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_382 = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_386 = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_390 = _RAND_16[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_394 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_398 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_402 = _RAND_19[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_406 = _RAND_20[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_410 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_414 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_418 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_422 = _RAND_24[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_426 = _RAND_25[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_430 = _RAND_26[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_434 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_438 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_442 = _RAND_29[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_446 = _RAND_30[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_450 = _RAND_31[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_454 = _RAND_32[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_458 = _RAND_33[27:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_462 = _RAND_34[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_466 = _RAND_35[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_470 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_327 <= 21'h1;
    end else begin
      if (_T_95) begin
        _T_327 <= _T_324;
      end
    end
    if (reset) begin
      _T_331 <= 5'h0;
    end else begin
      if (_T_98) begin
        _T_331 <= _T_328;
      end
    end
    if (reset) begin
      _T_335 <= 5'h0;
    end else begin
      if (_T_98) begin
        _T_335 <= _T_332;
      end
    end
    if (reset) begin
      _T_339 <= 5'h0;
    end else begin
      if (_T_101) begin
        _T_339 <= _T_328;
      end
    end
    if (reset) begin
      _T_343 <= 3'h0;
    end else begin
      if (_T_104) begin
        _T_343 <= _T_340;
      end
    end
    if (reset) begin
      _T_347 <= 3'h0;
    end else begin
      if (_T_104) begin
        _T_347 <= _T_344;
      end
    end
    if (reset) begin
      _T_350 <= 32'h0;
    end else begin
      if (_T_107) begin
        _T_350 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_354 <= 1'h0;
    end else begin
      if (_T_110) begin
        _T_354 <= _T_351;
      end
    end
    if (reset) begin
      _T_358 <= 13'h0;
    end else begin
      if (_T_113) begin
        _T_358 <= _T_355;
      end
    end
    if (reset) begin
      _T_362 <= 13'h0;
    end else begin
      if (_T_113) begin
        _T_362 <= _T_359;
      end
    end
    if (reset) begin
      _T_366 <= 13'h0;
    end else begin
      if (_T_116) begin
        _T_366 <= _T_359;
      end
    end
    if (reset) begin
      _T_370 <= 13'h0;
    end else begin
      if (_T_119) begin
        _T_370 <= _T_355;
      end
    end
    if (reset) begin
      _T_374 <= 13'h0;
    end else begin
      if (_T_119) begin
        _T_374 <= _T_359;
      end
    end
    if (reset) begin
      _T_378 <= 13'h0;
    end else begin
      if (_T_122) begin
        _T_378 <= _T_359;
      end
    end
    if (reset) begin
      _T_382 <= 5'h0;
    end else begin
      if (_T_125) begin
        _T_382 <= _T_328;
      end
    end
    if (reset) begin
      _T_386 <= 5'h0;
    end else begin
      if (_T_125) begin
        _T_386 <= _T_332;
      end
    end
    if (reset) begin
      _T_390 <= 14'h0;
    end else begin
      if (_T_128) begin
        _T_390 <= _T_387;
      end
    end
    if (reset) begin
      _T_394 <= 1'h0;
    end else begin
      if (_T_131) begin
        _T_394 <= _T_351;
      end
    end
    if (reset) begin
      _T_398 <= 1'h0;
    end else begin
      if (_T_131) begin
        _T_398 <= _T_395;
      end
    end
    if (reset) begin
      _T_402 <= 2'h1;
    end else begin
      if (_T_131) begin
        _T_402 <= _T_399;
      end
    end
    if (reset) begin
      _T_406 <= 2'h1;
    end else begin
      if (_T_131) begin
        _T_406 <= _T_403;
      end
    end
    if (reset) begin
      _T_410 <= 1'h0;
    end else begin
      if (_T_131) begin
        _T_410 <= _T_407;
      end
    end
    if (reset) begin
      _T_414 <= 1'h0;
    end else begin
      if (_T_131) begin
        _T_414 <= _T_411;
      end
    end
    if (reset) begin
      _T_418 <= 1'h0;
    end else begin
      if (_T_131) begin
        _T_418 <= _T_415;
      end
    end
    if (reset) begin
      _T_422 <= 2'h0;
    end else begin
      if (_T_137) begin
        _T_422 <= _T_419;
      end
    end
    if (reset) begin
      _T_426 <= 2'h0;
    end else begin
      if (_T_140) begin
        _T_426 <= _T_419;
      end
    end
    if (reset) begin
      _T_430 <= 12'h1;
    end else begin
      if (_T_143) begin
        _T_430 <= _T_427;
      end
    end
    if (reset) begin
      _T_434 <= 32'h0;
    end else begin
      if (_T_146) begin
        _T_434 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_438 <= 1'h0;
    end else begin
      if (_T_149) begin
        _T_438 <= _T_351;
      end
    end
    if (reset) begin
      _T_442 <= 5'h0;
    end else begin
      if (_T_152) begin
        _T_442 <= _T_332;
      end
    end
    if (reset) begin
      _T_446 <= 5'h0;
    end else begin
      if (_T_152) begin
        _T_446 <= _T_328;
      end
    end
    if (reset) begin
      _T_450 <= 13'h0;
    end else begin
      if (_T_155) begin
        _T_450 <= _T_359;
      end
    end
    if (reset) begin
      _T_454 <= 13'h0;
    end else begin
      if (_T_155) begin
        _T_454 <= _T_355;
      end
    end
    if (reset) begin
      _T_458 <= 28'h0;
    end else begin
      if (_T_158) begin
        _T_458 <= _T_455;
      end
    end
    if (reset) begin
      _T_462 <= 5'h0;
    end else begin
      if (_T_161) begin
        _T_462 <= _T_328;
      end
    end
    if (reset) begin
      _T_466 <= 5'h0;
    end else begin
      if (_T_161) begin
        _T_466 <= _T_332;
      end
    end
    if (reset) begin
      _T_470 <= 16'h0;
    end else begin
      if (_T_164) begin
        _T_470 <= _T_467;
      end
    end
  end
endmodule
module NV_NVDLA_CSB_LOGIC( // @[:@780.2]
  input         reset, // @[:@782.4]
  input         io_clk, // @[:@783.4]
  input         io_csb2dp_req_valid, // @[:@783.4]
  input  [62:0] io_csb2dp_req_bits, // @[:@783.4]
  output        io_csb2dp_resp_valid, // @[:@783.4]
  output [33:0] io_csb2dp_resp_bits, // @[:@783.4]
  input  [31:0] io_reg_rd_data, // @[:@783.4]
  output [11:0] io_reg_offset, // @[:@783.4]
  output [31:0] io_reg_wr_data, // @[:@783.4]
  output        io_reg_wr_en // @[:@783.4]
);
  reg  _T_43; // @[NV_NVDLA_CSB_LOGIC.scala 45:27:@785.4]
  reg [31:0] _RAND_0;
  reg [62:0] _T_46; // @[NV_NVDLA_CSB_LOGIC.scala 46:25:@786.4]
  reg [63:0] _RAND_1;
  wire [62:0] _GEN_0; // @[NV_NVDLA_CSB_LOGIC.scala 49:30:@788.4]
  wire [21:0] _T_47; // @[NV_NVDLA_CSB_LOGIC.scala 54:26:@791.4]
  wire  _T_49; // @[NV_NVDLA_CSB_LOGIC.scala 56:27:@793.4]
  wire  _T_50; // @[NV_NVDLA_CSB_LOGIC.scala 57:29:@794.4]
  wire [23:0] _T_56; // @[Cat.scala 30:58:@799.4]
  wire  _T_58; // @[NV_NVDLA_CSB_LOGIC.scala 68:32:@804.4]
  wire  _T_59; // @[NV_NVDLA_CSB_LOGIC.scala 68:30:@805.4]
  wire [33:0] _T_63; // @[Cat.scala 30:58:@807.4]
  reg [33:0] _T_71; // @[NV_NVDLA_CSB_LOGIC.scala 83:37:@810.4]
  reg [63:0] _RAND_2;
  reg  _T_74; // @[NV_NVDLA_CSB_LOGIC.scala 84:40:@811.4]
  reg [31:0] _RAND_3;
  wire  _T_75; // @[NV_NVDLA_CSB_LOGIC.scala 89:28:@816.6]
  wire [33:0] _GEN_1; // @[NV_NVDLA_CSB_LOGIC.scala 89:42:@817.6]
  wire [33:0] _GEN_2; // @[NV_NVDLA_CSB_LOGIC.scala 86:20:@812.4]
  wire  _T_77; // @[NV_NVDLA_CSB_LOGIC.scala 92:59:@821.4]
  assign _GEN_0 = io_csb2dp_req_valid ? io_csb2dp_req_bits : _T_46; // @[NV_NVDLA_CSB_LOGIC.scala 49:30:@788.4]
  assign _T_47 = _T_46[21:0]; // @[NV_NVDLA_CSB_LOGIC.scala 54:26:@791.4]
  assign _T_49 = _T_46[54]; // @[NV_NVDLA_CSB_LOGIC.scala 56:27:@793.4]
  assign _T_50 = _T_46[55]; // @[NV_NVDLA_CSB_LOGIC.scala 57:29:@794.4]
  assign _T_56 = {_T_47,2'h0}; // @[Cat.scala 30:58:@799.4]
  assign _T_58 = ~ _T_49; // @[NV_NVDLA_CSB_LOGIC.scala 68:32:@804.4]
  assign _T_59 = _T_43 & _T_58; // @[NV_NVDLA_CSB_LOGIC.scala 68:30:@805.4]
  assign _T_63 = {2'h0,io_reg_rd_data}; // @[Cat.scala 30:58:@807.4]
  assign _T_75 = io_reg_wr_en & _T_50; // @[NV_NVDLA_CSB_LOGIC.scala 89:28:@816.6]
  assign _GEN_1 = _T_75 ? 34'h200000000 : _T_71; // @[NV_NVDLA_CSB_LOGIC.scala 89:42:@817.6]
  assign _GEN_2 = _T_59 ? _T_63 : _GEN_1; // @[NV_NVDLA_CSB_LOGIC.scala 86:20:@812.4]
  assign _T_77 = _T_75 | _T_59; // @[NV_NVDLA_CSB_LOGIC.scala 92:59:@821.4]
  assign io_csb2dp_resp_valid = _T_74; // @[NV_NVDLA_CSB_LOGIC.scala 95:26:@824.4]
  assign io_csb2dp_resp_bits = _T_71; // @[NV_NVDLA_CSB_LOGIC.scala 94:25:@823.4]
  assign io_reg_offset = _T_56[11:0]; // @[NV_NVDLA_CSB_LOGIC.scala 65:19:@800.4]
  assign io_reg_wr_data = _T_46[53:22]; // @[NV_NVDLA_CSB_LOGIC.scala 66:20:@801.4]
  assign io_reg_wr_en = _T_43 & _T_49; // @[NV_NVDLA_CSB_LOGIC.scala 67:18:@803.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_43 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  _T_46 = _RAND_1[62:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  _T_71 = _RAND_2[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_74 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_clk) begin
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      _T_43 <= io_csb2dp_req_valid;
    end
    if (reset) begin
      _T_46 <= 63'h0;
    end else begin
      if (io_csb2dp_req_valid) begin
        _T_46 <= io_csb2dp_req_bits;
      end
    end
    if (reset) begin
      _T_71 <= 34'h0;
    end else begin
      if (_T_59) begin
        _T_71 <= _T_63;
      end else begin
        if (_T_75) begin
          _T_71 <= 34'h200000000;
        end
      end
    end
    if (reset) begin
      _T_74 <= 1'h0;
    end else begin
      _T_74 <= _T_77;
    end
  end
endmodule
module NV_NVDLA_CSC_regfile( // @[:@826.2]
  input         reset, // @[:@828.4]
  input         io_nvdla_core_clk, // @[:@829.4]
  input         io_csb2csc_req_valid, // @[:@829.4]
  input  [62:0] io_csb2csc_req_bits, // @[:@829.4]
  output        io_csb2csc_resp_valid, // @[:@829.4]
  output [33:0] io_csb2csc_resp_bits, // @[:@829.4]
  output        io_reg2dp_op_en, // @[:@829.4]
  output [20:0] io_reg2dp_field_atomics, // @[:@829.4]
  output [4:0]  io_reg2dp_field_data_bank, // @[:@829.4]
  output [4:0]  io_reg2dp_field_weight_bank, // @[:@829.4]
  output [2:0]  io_reg2dp_field_conv_x_stride_ext, // @[:@829.4]
  output [2:0]  io_reg2dp_field_conv_y_stride_ext, // @[:@829.4]
  output        io_reg2dp_field_datain_format, // @[:@829.4]
  output [12:0] io_reg2dp_field_datain_height_ext, // @[:@829.4]
  output [12:0] io_reg2dp_field_datain_width_ext, // @[:@829.4]
  output [12:0] io_reg2dp_field_datain_channel_ext, // @[:@829.4]
  output [12:0] io_reg2dp_field_dataout_height, // @[:@829.4]
  output [12:0] io_reg2dp_field_dataout_width, // @[:@829.4]
  output [4:0]  io_reg2dp_field_x_dilation_ext, // @[:@829.4]
  output [4:0]  io_reg2dp_field_y_dilation_ext, // @[:@829.4]
  output [13:0] io_reg2dp_field_entries, // @[:@829.4]
  output        io_reg2dp_field_conv_mode, // @[:@829.4]
  output        io_reg2dp_field_data_reuse, // @[:@829.4]
  output        io_reg2dp_field_skip_data_rls, // @[:@829.4]
  output        io_reg2dp_field_skip_weight_rls, // @[:@829.4]
  output        io_reg2dp_field_weight_reuse, // @[:@829.4]
  output [1:0]  io_reg2dp_field_y_extension, // @[:@829.4]
  output [11:0] io_reg2dp_field_rls_slices, // @[:@829.4]
  output [31:0] io_reg2dp_field_weight_bytes, // @[:@829.4]
  output        io_reg2dp_field_weight_format, // @[:@829.4]
  output [4:0]  io_reg2dp_field_weight_height_ext, // @[:@829.4]
  output [4:0]  io_reg2dp_field_weight_width_ext, // @[:@829.4]
  output [12:0] io_reg2dp_field_weight_channel_ext, // @[:@829.4]
  output [12:0] io_reg2dp_field_weight_kernel, // @[:@829.4]
  output [27:0] io_reg2dp_field_wmb_bytes, // @[:@829.4]
  output [4:0]  io_reg2dp_field_pad_left, // @[:@829.4]
  output [4:0]  io_reg2dp_field_pad_top, // @[:@829.4]
  output [15:0] io_reg2dp_field_pad_value, // @[:@829.4]
  input         io_dp2reg_done // @[:@829.4]
);
  wire  NV_NVDLA_BASIC_REG_single_reset; // @[NV_NVDLA_CSC_regfile.scala 58:30:@837.4]
  wire  NV_NVDLA_BASIC_REG_single_io_nvdla_core_clk; // @[NV_NVDLA_CSC_regfile.scala 58:30:@837.4]
  wire [31:0] NV_NVDLA_BASIC_REG_single_io_reg_rd_data; // @[NV_NVDLA_CSC_regfile.scala 58:30:@837.4]
  wire [11:0] NV_NVDLA_BASIC_REG_single_io_reg_offset; // @[NV_NVDLA_CSC_regfile.scala 58:30:@837.4]
  wire [31:0] NV_NVDLA_BASIC_REG_single_io_reg_wr_data; // @[NV_NVDLA_CSC_regfile.scala 58:30:@837.4]
  wire  NV_NVDLA_BASIC_REG_single_io_reg_wr_en; // @[NV_NVDLA_CSC_regfile.scala 58:30:@837.4]
  wire  NV_NVDLA_BASIC_REG_single_io_producer; // @[NV_NVDLA_CSC_regfile.scala 58:30:@837.4]
  wire  NV_NVDLA_BASIC_REG_single_io_consumer; // @[NV_NVDLA_CSC_regfile.scala 58:30:@837.4]
  wire [1:0] NV_NVDLA_BASIC_REG_single_io_status_0; // @[NV_NVDLA_CSC_regfile.scala 58:30:@837.4]
  wire [1:0] NV_NVDLA_BASIC_REG_single_io_status_1; // @[NV_NVDLA_CSC_regfile.scala 58:30:@837.4]
  wire  NV_NVDLA_CSC_dual_reg_reset; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire  NV_NVDLA_CSC_dual_reg_io_nvdla_core_clk; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [31:0] NV_NVDLA_CSC_dual_reg_io_reg_rd_data; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [11:0] NV_NVDLA_CSC_dual_reg_io_reg_offset; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [31:0] NV_NVDLA_CSC_dual_reg_io_reg_wr_data; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire  NV_NVDLA_CSC_dual_reg_io_reg_wr_en; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [20:0] NV_NVDLA_CSC_dual_reg_io_field_atomics; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_io_field_data_bank; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_io_field_weight_bank; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_io_field_batches; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [2:0] NV_NVDLA_CSC_dual_reg_io_field_conv_x_stride_ext; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [2:0] NV_NVDLA_CSC_dual_reg_io_field_conv_y_stride_ext; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [31:0] NV_NVDLA_CSC_dual_reg_io_field_cya; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire  NV_NVDLA_CSC_dual_reg_io_field_datain_format; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [12:0] NV_NVDLA_CSC_dual_reg_io_field_datain_height_ext; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [12:0] NV_NVDLA_CSC_dual_reg_io_field_datain_width_ext; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [12:0] NV_NVDLA_CSC_dual_reg_io_field_datain_channel_ext; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [12:0] NV_NVDLA_CSC_dual_reg_io_field_dataout_height; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [12:0] NV_NVDLA_CSC_dual_reg_io_field_dataout_width; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [12:0] NV_NVDLA_CSC_dual_reg_io_field_dataout_channel; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_io_field_x_dilation_ext; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_io_field_y_dilation_ext; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [13:0] NV_NVDLA_CSC_dual_reg_io_field_entries; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire  NV_NVDLA_CSC_dual_reg_io_field_conv_mode; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire  NV_NVDLA_CSC_dual_reg_io_field_data_reuse; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [1:0] NV_NVDLA_CSC_dual_reg_io_field_in_precision; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [1:0] NV_NVDLA_CSC_dual_reg_io_field_proc_precision; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire  NV_NVDLA_CSC_dual_reg_io_field_skip_data_rls; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire  NV_NVDLA_CSC_dual_reg_io_field_skip_weight_rls; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire  NV_NVDLA_CSC_dual_reg_io_field_weight_reuse; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [1:0] NV_NVDLA_CSC_dual_reg_io_field_y_extension; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [1:0] NV_NVDLA_CSC_dual_reg_io_field_pra_truncate; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [11:0] NV_NVDLA_CSC_dual_reg_io_field_rls_slices; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [31:0] NV_NVDLA_CSC_dual_reg_io_field_weight_bytes; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire  NV_NVDLA_CSC_dual_reg_io_field_weight_format; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_io_field_weight_height_ext; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_io_field_weight_width_ext; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [12:0] NV_NVDLA_CSC_dual_reg_io_field_weight_channel_ext; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [12:0] NV_NVDLA_CSC_dual_reg_io_field_weight_kernel; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [27:0] NV_NVDLA_CSC_dual_reg_io_field_wmb_bytes; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_io_field_pad_left; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_io_field_pad_top; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire [15:0] NV_NVDLA_CSC_dual_reg_io_field_pad_value; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire  NV_NVDLA_CSC_dual_reg_io_op_en_trigger; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire  NV_NVDLA_CSC_dual_reg_io_op_en; // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
  wire  NV_NVDLA_CSC_dual_reg_1_reset; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire  NV_NVDLA_CSC_dual_reg_1_io_nvdla_core_clk; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [31:0] NV_NVDLA_CSC_dual_reg_1_io_reg_rd_data; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [11:0] NV_NVDLA_CSC_dual_reg_1_io_reg_offset; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [31:0] NV_NVDLA_CSC_dual_reg_1_io_reg_wr_data; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire  NV_NVDLA_CSC_dual_reg_1_io_reg_wr_en; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [20:0] NV_NVDLA_CSC_dual_reg_1_io_field_atomics; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_1_io_field_data_bank; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_1_io_field_weight_bank; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_1_io_field_batches; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [2:0] NV_NVDLA_CSC_dual_reg_1_io_field_conv_x_stride_ext; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [2:0] NV_NVDLA_CSC_dual_reg_1_io_field_conv_y_stride_ext; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [31:0] NV_NVDLA_CSC_dual_reg_1_io_field_cya; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire  NV_NVDLA_CSC_dual_reg_1_io_field_datain_format; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [12:0] NV_NVDLA_CSC_dual_reg_1_io_field_datain_height_ext; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [12:0] NV_NVDLA_CSC_dual_reg_1_io_field_datain_width_ext; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [12:0] NV_NVDLA_CSC_dual_reg_1_io_field_datain_channel_ext; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [12:0] NV_NVDLA_CSC_dual_reg_1_io_field_dataout_height; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [12:0] NV_NVDLA_CSC_dual_reg_1_io_field_dataout_width; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [12:0] NV_NVDLA_CSC_dual_reg_1_io_field_dataout_channel; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_1_io_field_x_dilation_ext; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_1_io_field_y_dilation_ext; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [13:0] NV_NVDLA_CSC_dual_reg_1_io_field_entries; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire  NV_NVDLA_CSC_dual_reg_1_io_field_conv_mode; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire  NV_NVDLA_CSC_dual_reg_1_io_field_data_reuse; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [1:0] NV_NVDLA_CSC_dual_reg_1_io_field_in_precision; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [1:0] NV_NVDLA_CSC_dual_reg_1_io_field_proc_precision; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire  NV_NVDLA_CSC_dual_reg_1_io_field_skip_data_rls; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire  NV_NVDLA_CSC_dual_reg_1_io_field_skip_weight_rls; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire  NV_NVDLA_CSC_dual_reg_1_io_field_weight_reuse; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [1:0] NV_NVDLA_CSC_dual_reg_1_io_field_y_extension; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [1:0] NV_NVDLA_CSC_dual_reg_1_io_field_pra_truncate; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [11:0] NV_NVDLA_CSC_dual_reg_1_io_field_rls_slices; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [31:0] NV_NVDLA_CSC_dual_reg_1_io_field_weight_bytes; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire  NV_NVDLA_CSC_dual_reg_1_io_field_weight_format; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_1_io_field_weight_height_ext; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_1_io_field_weight_width_ext; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [12:0] NV_NVDLA_CSC_dual_reg_1_io_field_weight_channel_ext; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [12:0] NV_NVDLA_CSC_dual_reg_1_io_field_weight_kernel; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [27:0] NV_NVDLA_CSC_dual_reg_1_io_field_wmb_bytes; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_1_io_field_pad_left; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [4:0] NV_NVDLA_CSC_dual_reg_1_io_field_pad_top; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire [15:0] NV_NVDLA_CSC_dual_reg_1_io_field_pad_value; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire  NV_NVDLA_CSC_dual_reg_1_io_op_en_trigger; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire  NV_NVDLA_CSC_dual_reg_1_io_op_en; // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
  wire  NV_NVDLA_CSB_LOGIC_reset; // @[NV_NVDLA_CSC_regfile.scala 162:27:@953.4]
  wire  NV_NVDLA_CSB_LOGIC_io_clk; // @[NV_NVDLA_CSC_regfile.scala 162:27:@953.4]
  wire  NV_NVDLA_CSB_LOGIC_io_csb2dp_req_valid; // @[NV_NVDLA_CSC_regfile.scala 162:27:@953.4]
  wire [62:0] NV_NVDLA_CSB_LOGIC_io_csb2dp_req_bits; // @[NV_NVDLA_CSC_regfile.scala 162:27:@953.4]
  wire  NV_NVDLA_CSB_LOGIC_io_csb2dp_resp_valid; // @[NV_NVDLA_CSC_regfile.scala 162:27:@953.4]
  wire [33:0] NV_NVDLA_CSB_LOGIC_io_csb2dp_resp_bits; // @[NV_NVDLA_CSC_regfile.scala 162:27:@953.4]
  wire [31:0] NV_NVDLA_CSB_LOGIC_io_reg_rd_data; // @[NV_NVDLA_CSC_regfile.scala 162:27:@953.4]
  wire [11:0] NV_NVDLA_CSB_LOGIC_io_reg_offset; // @[NV_NVDLA_CSC_regfile.scala 162:27:@953.4]
  wire [31:0] NV_NVDLA_CSB_LOGIC_io_reg_wr_data; // @[NV_NVDLA_CSC_regfile.scala 162:27:@953.4]
  wire  NV_NVDLA_CSB_LOGIC_io_reg_wr_en; // @[NV_NVDLA_CSC_regfile.scala 162:27:@953.4]
  reg  _T_105; // @[NV_NVDLA_CSC_regfile.scala 50:34:@831.4]
  reg [31:0] _RAND_0;
  reg  _T_120; // @[NV_NVDLA_CSC_regfile.scala 72:34:@848.4]
  reg [31:0] _RAND_1;
  reg  _T_125; // @[NV_NVDLA_CSC_regfile.scala 85:34:@858.4]
  reg [31:0] _RAND_2;
  wire  _T_126; // @[NV_NVDLA_CSC_regfile.scala 103:28:@868.6]
  wire  _GEN_0; // @[NV_NVDLA_CSC_regfile.scala 102:25:@867.4]
  wire  _T_128; // @[NV_NVDLA_CSC_regfile.scala 111:44:@871.4]
  wire [1:0] _T_134; // @[NV_NVDLA_CSC_regfile.scala 112:27:@873.4]
  wire  _T_137; // @[NV_NVDLA_CSC_regfile.scala 115:44:@876.4]
  wire  _T_140; // @[NV_NVDLA_CSC_regfile.scala 116:44:@877.4]
  wire [1:0] _T_143; // @[NV_NVDLA_CSC_regfile.scala 116:27:@878.4]
  reg [2:0] _T_147; // @[NV_NVDLA_CSC_regfile.scala 124:35:@881.4]
  reg [31:0] _RAND_3;
  wire  _T_148; // @[NV_NVDLA_CSC_regfile.scala 126:28:@882.4]
  wire  _T_149; // @[NV_NVDLA_CSC_regfile.scala 126:45:@883.4]
  wire [31:0] _T_113; // @[NV_NVDLA_CSC_regfile.scala 55:27:@835.4 NV_NVDLA_CSC_regfile.scala 167:17:@964.4]
  wire  _T_150; // @[NV_NVDLA_CSC_regfile.scala 126:83:@884.4]
  wire  _T_153; // @[NV_NVDLA_CSC_regfile.scala 127:43:@886.4]
  wire  _T_155; // @[NV_NVDLA_CSC_regfile.scala 127:27:@887.4]
  wire  _T_156; // @[NV_NVDLA_CSC_regfile.scala 126:27:@888.4]
  wire  _T_157; // @[NV_NVDLA_CSC_regfile.scala 129:28:@890.4]
  wire  _T_158; // @[NV_NVDLA_CSC_regfile.scala 129:45:@891.4]
  wire  _T_162; // @[NV_NVDLA_CSC_regfile.scala 130:43:@894.4]
  wire  _T_164; // @[NV_NVDLA_CSC_regfile.scala 130:27:@895.4]
  wire  _T_165; // @[NV_NVDLA_CSC_regfile.scala 129:27:@896.4]
  wire  _T_166; // @[NV_NVDLA_CSC_regfile.scala 132:31:@898.4]
  wire [1:0] _T_168; // @[NV_NVDLA_CSC_regfile.scala 134:83:@899.4]
  wire [2:0] _T_169; // @[Cat.scala 30:58:@900.4]
  wire [2:0] _T_170; // @[NV_NVDLA_CSC_regfile.scala 134:28:@901.4]
  wire [11:0] _T_111; // @[NV_NVDLA_CSC_regfile.scala 54:26:@834.4 NV_NVDLA_CSC_regfile.scala 165:16:@962.4]
  wire [31:0] _GEN_4; // @[NV_NVDLA_CSC_regfile.scala 145:41:@922.4]
  wire  _T_187; // @[NV_NVDLA_CSC_regfile.scala 145:41:@922.4]
  wire  _T_193; // @[NV_NVDLA_CSC_regfile.scala 146:39:@925.4]
  wire  _T_195; // @[NV_NVDLA_CSC_regfile.scala 146:83:@926.4]
  wire  _T_196; // @[NV_NVDLA_CSC_regfile.scala 146:64:@927.4]
  wire  _T_201; // @[NV_NVDLA_CSC_regfile.scala 147:83:@930.4]
  wire  _T_202; // @[NV_NVDLA_CSC_regfile.scala 147:64:@931.4]
  wire  _T_184; // @[NV_NVDLA_CSC_regfile.scala 144:25:@920.4 NV_NVDLA_CSC_regfile.scala 166:15:@963.4]
  wire  _T_204; // @[NV_NVDLA_CSC_regfile.scala 150:31:@934.4]
  wire  _T_208; // @[NV_NVDLA_CSC_regfile.scala 151:31:@938.4]
  wire [31:0] _T_215; // @[Bitwise.scala 72:12:@943.4]
  wire [31:0] _T_216; // @[NV_NVDLA_CSC_regfile.scala 153:43:@944.4]
  wire [31:0] _T_220; // @[Bitwise.scala 72:12:@946.4]
  wire [31:0] _T_221; // @[NV_NVDLA_CSC_regfile.scala 154:44:@947.4]
  wire [31:0] _T_222; // @[NV_NVDLA_CSC_regfile.scala 153:59:@948.4]
  wire [31:0] _T_226; // @[Bitwise.scala 72:12:@950.4]
  wire [31:0] _T_227; // @[NV_NVDLA_CSC_regfile.scala 155:43:@951.4]
  NV_NVDLA_BASIC_REG_single NV_NVDLA_BASIC_REG_single ( // @[NV_NVDLA_CSC_regfile.scala 58:30:@837.4]
    .reset(NV_NVDLA_BASIC_REG_single_reset),
    .io_nvdla_core_clk(NV_NVDLA_BASIC_REG_single_io_nvdla_core_clk),
    .io_reg_rd_data(NV_NVDLA_BASIC_REG_single_io_reg_rd_data),
    .io_reg_offset(NV_NVDLA_BASIC_REG_single_io_reg_offset),
    .io_reg_wr_data(NV_NVDLA_BASIC_REG_single_io_reg_wr_data),
    .io_reg_wr_en(NV_NVDLA_BASIC_REG_single_io_reg_wr_en),
    .io_producer(NV_NVDLA_BASIC_REG_single_io_producer),
    .io_consumer(NV_NVDLA_BASIC_REG_single_io_consumer),
    .io_status_0(NV_NVDLA_BASIC_REG_single_io_status_0),
    .io_status_1(NV_NVDLA_BASIC_REG_single_io_status_1)
  );
  NV_NVDLA_CSC_dual_reg NV_NVDLA_CSC_dual_reg ( // @[NV_NVDLA_CSC_regfile.scala 74:31:@849.4]
    .reset(NV_NVDLA_CSC_dual_reg_reset),
    .io_nvdla_core_clk(NV_NVDLA_CSC_dual_reg_io_nvdla_core_clk),
    .io_reg_rd_data(NV_NVDLA_CSC_dual_reg_io_reg_rd_data),
    .io_reg_offset(NV_NVDLA_CSC_dual_reg_io_reg_offset),
    .io_reg_wr_data(NV_NVDLA_CSC_dual_reg_io_reg_wr_data),
    .io_reg_wr_en(NV_NVDLA_CSC_dual_reg_io_reg_wr_en),
    .io_field_atomics(NV_NVDLA_CSC_dual_reg_io_field_atomics),
    .io_field_data_bank(NV_NVDLA_CSC_dual_reg_io_field_data_bank),
    .io_field_weight_bank(NV_NVDLA_CSC_dual_reg_io_field_weight_bank),
    .io_field_batches(NV_NVDLA_CSC_dual_reg_io_field_batches),
    .io_field_conv_x_stride_ext(NV_NVDLA_CSC_dual_reg_io_field_conv_x_stride_ext),
    .io_field_conv_y_stride_ext(NV_NVDLA_CSC_dual_reg_io_field_conv_y_stride_ext),
    .io_field_cya(NV_NVDLA_CSC_dual_reg_io_field_cya),
    .io_field_datain_format(NV_NVDLA_CSC_dual_reg_io_field_datain_format),
    .io_field_datain_height_ext(NV_NVDLA_CSC_dual_reg_io_field_datain_height_ext),
    .io_field_datain_width_ext(NV_NVDLA_CSC_dual_reg_io_field_datain_width_ext),
    .io_field_datain_channel_ext(NV_NVDLA_CSC_dual_reg_io_field_datain_channel_ext),
    .io_field_dataout_height(NV_NVDLA_CSC_dual_reg_io_field_dataout_height),
    .io_field_dataout_width(NV_NVDLA_CSC_dual_reg_io_field_dataout_width),
    .io_field_dataout_channel(NV_NVDLA_CSC_dual_reg_io_field_dataout_channel),
    .io_field_x_dilation_ext(NV_NVDLA_CSC_dual_reg_io_field_x_dilation_ext),
    .io_field_y_dilation_ext(NV_NVDLA_CSC_dual_reg_io_field_y_dilation_ext),
    .io_field_entries(NV_NVDLA_CSC_dual_reg_io_field_entries),
    .io_field_conv_mode(NV_NVDLA_CSC_dual_reg_io_field_conv_mode),
    .io_field_data_reuse(NV_NVDLA_CSC_dual_reg_io_field_data_reuse),
    .io_field_in_precision(NV_NVDLA_CSC_dual_reg_io_field_in_precision),
    .io_field_proc_precision(NV_NVDLA_CSC_dual_reg_io_field_proc_precision),
    .io_field_skip_data_rls(NV_NVDLA_CSC_dual_reg_io_field_skip_data_rls),
    .io_field_skip_weight_rls(NV_NVDLA_CSC_dual_reg_io_field_skip_weight_rls),
    .io_field_weight_reuse(NV_NVDLA_CSC_dual_reg_io_field_weight_reuse),
    .io_field_y_extension(NV_NVDLA_CSC_dual_reg_io_field_y_extension),
    .io_field_pra_truncate(NV_NVDLA_CSC_dual_reg_io_field_pra_truncate),
    .io_field_rls_slices(NV_NVDLA_CSC_dual_reg_io_field_rls_slices),
    .io_field_weight_bytes(NV_NVDLA_CSC_dual_reg_io_field_weight_bytes),
    .io_field_weight_format(NV_NVDLA_CSC_dual_reg_io_field_weight_format),
    .io_field_weight_height_ext(NV_NVDLA_CSC_dual_reg_io_field_weight_height_ext),
    .io_field_weight_width_ext(NV_NVDLA_CSC_dual_reg_io_field_weight_width_ext),
    .io_field_weight_channel_ext(NV_NVDLA_CSC_dual_reg_io_field_weight_channel_ext),
    .io_field_weight_kernel(NV_NVDLA_CSC_dual_reg_io_field_weight_kernel),
    .io_field_wmb_bytes(NV_NVDLA_CSC_dual_reg_io_field_wmb_bytes),
    .io_field_pad_left(NV_NVDLA_CSC_dual_reg_io_field_pad_left),
    .io_field_pad_top(NV_NVDLA_CSC_dual_reg_io_field_pad_top),
    .io_field_pad_value(NV_NVDLA_CSC_dual_reg_io_field_pad_value),
    .io_op_en_trigger(NV_NVDLA_CSC_dual_reg_io_op_en_trigger),
    .io_op_en(NV_NVDLA_CSC_dual_reg_io_op_en)
  );
  NV_NVDLA_CSC_dual_reg NV_NVDLA_CSC_dual_reg_1 ( // @[NV_NVDLA_CSC_regfile.scala 87:31:@859.4]
    .reset(NV_NVDLA_CSC_dual_reg_1_reset),
    .io_nvdla_core_clk(NV_NVDLA_CSC_dual_reg_1_io_nvdla_core_clk),
    .io_reg_rd_data(NV_NVDLA_CSC_dual_reg_1_io_reg_rd_data),
    .io_reg_offset(NV_NVDLA_CSC_dual_reg_1_io_reg_offset),
    .io_reg_wr_data(NV_NVDLA_CSC_dual_reg_1_io_reg_wr_data),
    .io_reg_wr_en(NV_NVDLA_CSC_dual_reg_1_io_reg_wr_en),
    .io_field_atomics(NV_NVDLA_CSC_dual_reg_1_io_field_atomics),
    .io_field_data_bank(NV_NVDLA_CSC_dual_reg_1_io_field_data_bank),
    .io_field_weight_bank(NV_NVDLA_CSC_dual_reg_1_io_field_weight_bank),
    .io_field_batches(NV_NVDLA_CSC_dual_reg_1_io_field_batches),
    .io_field_conv_x_stride_ext(NV_NVDLA_CSC_dual_reg_1_io_field_conv_x_stride_ext),
    .io_field_conv_y_stride_ext(NV_NVDLA_CSC_dual_reg_1_io_field_conv_y_stride_ext),
    .io_field_cya(NV_NVDLA_CSC_dual_reg_1_io_field_cya),
    .io_field_datain_format(NV_NVDLA_CSC_dual_reg_1_io_field_datain_format),
    .io_field_datain_height_ext(NV_NVDLA_CSC_dual_reg_1_io_field_datain_height_ext),
    .io_field_datain_width_ext(NV_NVDLA_CSC_dual_reg_1_io_field_datain_width_ext),
    .io_field_datain_channel_ext(NV_NVDLA_CSC_dual_reg_1_io_field_datain_channel_ext),
    .io_field_dataout_height(NV_NVDLA_CSC_dual_reg_1_io_field_dataout_height),
    .io_field_dataout_width(NV_NVDLA_CSC_dual_reg_1_io_field_dataout_width),
    .io_field_dataout_channel(NV_NVDLA_CSC_dual_reg_1_io_field_dataout_channel),
    .io_field_x_dilation_ext(NV_NVDLA_CSC_dual_reg_1_io_field_x_dilation_ext),
    .io_field_y_dilation_ext(NV_NVDLA_CSC_dual_reg_1_io_field_y_dilation_ext),
    .io_field_entries(NV_NVDLA_CSC_dual_reg_1_io_field_entries),
    .io_field_conv_mode(NV_NVDLA_CSC_dual_reg_1_io_field_conv_mode),
    .io_field_data_reuse(NV_NVDLA_CSC_dual_reg_1_io_field_data_reuse),
    .io_field_in_precision(NV_NVDLA_CSC_dual_reg_1_io_field_in_precision),
    .io_field_proc_precision(NV_NVDLA_CSC_dual_reg_1_io_field_proc_precision),
    .io_field_skip_data_rls(NV_NVDLA_CSC_dual_reg_1_io_field_skip_data_rls),
    .io_field_skip_weight_rls(NV_NVDLA_CSC_dual_reg_1_io_field_skip_weight_rls),
    .io_field_weight_reuse(NV_NVDLA_CSC_dual_reg_1_io_field_weight_reuse),
    .io_field_y_extension(NV_NVDLA_CSC_dual_reg_1_io_field_y_extension),
    .io_field_pra_truncate(NV_NVDLA_CSC_dual_reg_1_io_field_pra_truncate),
    .io_field_rls_slices(NV_NVDLA_CSC_dual_reg_1_io_field_rls_slices),
    .io_field_weight_bytes(NV_NVDLA_CSC_dual_reg_1_io_field_weight_bytes),
    .io_field_weight_format(NV_NVDLA_CSC_dual_reg_1_io_field_weight_format),
    .io_field_weight_height_ext(NV_NVDLA_CSC_dual_reg_1_io_field_weight_height_ext),
    .io_field_weight_width_ext(NV_NVDLA_CSC_dual_reg_1_io_field_weight_width_ext),
    .io_field_weight_channel_ext(NV_NVDLA_CSC_dual_reg_1_io_field_weight_channel_ext),
    .io_field_weight_kernel(NV_NVDLA_CSC_dual_reg_1_io_field_weight_kernel),
    .io_field_wmb_bytes(NV_NVDLA_CSC_dual_reg_1_io_field_wmb_bytes),
    .io_field_pad_left(NV_NVDLA_CSC_dual_reg_1_io_field_pad_left),
    .io_field_pad_top(NV_NVDLA_CSC_dual_reg_1_io_field_pad_top),
    .io_field_pad_value(NV_NVDLA_CSC_dual_reg_1_io_field_pad_value),
    .io_op_en_trigger(NV_NVDLA_CSC_dual_reg_1_io_op_en_trigger),
    .io_op_en(NV_NVDLA_CSC_dual_reg_1_io_op_en)
  );
  NV_NVDLA_CSB_LOGIC NV_NVDLA_CSB_LOGIC ( // @[NV_NVDLA_CSC_regfile.scala 162:27:@953.4]
    .reset(NV_NVDLA_CSB_LOGIC_reset),
    .io_clk(NV_NVDLA_CSB_LOGIC_io_clk),
    .io_csb2dp_req_valid(NV_NVDLA_CSB_LOGIC_io_csb2dp_req_valid),
    .io_csb2dp_req_bits(NV_NVDLA_CSB_LOGIC_io_csb2dp_req_bits),
    .io_csb2dp_resp_valid(NV_NVDLA_CSB_LOGIC_io_csb2dp_resp_valid),
    .io_csb2dp_resp_bits(NV_NVDLA_CSB_LOGIC_io_csb2dp_resp_bits),
    .io_reg_rd_data(NV_NVDLA_CSB_LOGIC_io_reg_rd_data),
    .io_reg_offset(NV_NVDLA_CSB_LOGIC_io_reg_offset),
    .io_reg_wr_data(NV_NVDLA_CSB_LOGIC_io_reg_wr_data),
    .io_reg_wr_en(NV_NVDLA_CSB_LOGIC_io_reg_wr_en)
  );
  assign _T_126 = ~ _T_105; // @[NV_NVDLA_CSC_regfile.scala 103:28:@868.6]
  assign _GEN_0 = io_dp2reg_done ? _T_126 : _T_105; // @[NV_NVDLA_CSC_regfile.scala 102:25:@867.4]
  assign _T_128 = _T_120 == 1'h0; // @[NV_NVDLA_CSC_regfile.scala 111:44:@871.4]
  assign _T_134 = _T_105 ? 2'h2 : 2'h1; // @[NV_NVDLA_CSC_regfile.scala 112:27:@873.4]
  assign _T_137 = _T_125 == 1'h0; // @[NV_NVDLA_CSC_regfile.scala 115:44:@876.4]
  assign _T_140 = _T_105 == 1'h0; // @[NV_NVDLA_CSC_regfile.scala 116:44:@877.4]
  assign _T_143 = _T_140 ? 2'h2 : 2'h1; // @[NV_NVDLA_CSC_regfile.scala 116:27:@878.4]
  assign _T_148 = ~ _T_120; // @[NV_NVDLA_CSC_regfile.scala 126:28:@882.4]
  assign _T_149 = _T_148 & NV_NVDLA_CSC_dual_reg_io_op_en_trigger; // @[NV_NVDLA_CSC_regfile.scala 126:45:@883.4]
  assign _T_113 = NV_NVDLA_CSB_LOGIC_io_reg_wr_data; // @[NV_NVDLA_CSC_regfile.scala 55:27:@835.4 NV_NVDLA_CSC_regfile.scala 167:17:@964.4]
  assign _T_150 = _T_113[0]; // @[NV_NVDLA_CSC_regfile.scala 126:83:@884.4]
  assign _T_153 = io_dp2reg_done & _T_140; // @[NV_NVDLA_CSC_regfile.scala 127:43:@886.4]
  assign _T_155 = _T_153 ? 1'h0 : _T_120; // @[NV_NVDLA_CSC_regfile.scala 127:27:@887.4]
  assign _T_156 = _T_149 ? _T_150 : _T_155; // @[NV_NVDLA_CSC_regfile.scala 126:27:@888.4]
  assign _T_157 = ~ _T_125; // @[NV_NVDLA_CSC_regfile.scala 129:28:@890.4]
  assign _T_158 = _T_157 & NV_NVDLA_CSC_dual_reg_1_io_op_en_trigger; // @[NV_NVDLA_CSC_regfile.scala 129:45:@891.4]
  assign _T_162 = io_dp2reg_done & _T_105; // @[NV_NVDLA_CSC_regfile.scala 130:43:@894.4]
  assign _T_164 = _T_162 ? 1'h0 : _T_125; // @[NV_NVDLA_CSC_regfile.scala 130:27:@895.4]
  assign _T_165 = _T_158 ? _T_150 : _T_164; // @[NV_NVDLA_CSC_regfile.scala 129:27:@896.4]
  assign _T_166 = _T_105 ? _T_125 : _T_120; // @[NV_NVDLA_CSC_regfile.scala 132:31:@898.4]
  assign _T_168 = _T_147[1:0]; // @[NV_NVDLA_CSC_regfile.scala 134:83:@899.4]
  assign _T_169 = {_T_168,_T_166}; // @[Cat.scala 30:58:@900.4]
  assign _T_170 = io_dp2reg_done ? 3'h0 : _T_169; // @[NV_NVDLA_CSC_regfile.scala 134:28:@901.4]
  assign _T_111 = NV_NVDLA_CSB_LOGIC_io_reg_offset; // @[NV_NVDLA_CSC_regfile.scala 54:26:@834.4 NV_NVDLA_CSC_regfile.scala 165:16:@962.4]
  assign _GEN_4 = {{20'd0}, _T_111}; // @[NV_NVDLA_CSC_regfile.scala 145:41:@922.4]
  assign _T_187 = _GEN_4 < 32'h8; // @[NV_NVDLA_CSC_regfile.scala 145:41:@922.4]
  assign _T_193 = _GEN_4 >= 32'h8; // @[NV_NVDLA_CSC_regfile.scala 146:39:@925.4]
  assign _T_195 = NV_NVDLA_BASIC_REG_single_io_producer == 1'h0; // @[NV_NVDLA_CSC_regfile.scala 146:83:@926.4]
  assign _T_196 = _T_193 & _T_195; // @[NV_NVDLA_CSC_regfile.scala 146:64:@927.4]
  assign _T_201 = NV_NVDLA_BASIC_REG_single_io_producer; // @[NV_NVDLA_CSC_regfile.scala 147:83:@930.4]
  assign _T_202 = _T_193 & _T_201; // @[NV_NVDLA_CSC_regfile.scala 147:64:@931.4]
  assign _T_184 = NV_NVDLA_CSB_LOGIC_io_reg_wr_en; // @[NV_NVDLA_CSC_regfile.scala 144:25:@920.4 NV_NVDLA_CSC_regfile.scala 166:15:@963.4]
  assign _T_204 = _T_184 & _T_196; // @[NV_NVDLA_CSC_regfile.scala 150:31:@934.4]
  assign _T_208 = _T_184 & _T_202; // @[NV_NVDLA_CSC_regfile.scala 151:31:@938.4]
  assign _T_215 = _T_187 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@943.4]
  assign _T_216 = _T_215 & NV_NVDLA_BASIC_REG_single_io_reg_rd_data; // @[NV_NVDLA_CSC_regfile.scala 153:43:@944.4]
  assign _T_220 = _T_196 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@946.4]
  assign _T_221 = _T_220 & NV_NVDLA_CSC_dual_reg_io_reg_rd_data; // @[NV_NVDLA_CSC_regfile.scala 154:44:@947.4]
  assign _T_222 = _T_216 | _T_221; // @[NV_NVDLA_CSC_regfile.scala 153:59:@948.4]
  assign _T_226 = _T_202 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@950.4]
  assign _T_227 = _T_226 & NV_NVDLA_CSC_dual_reg_1_io_reg_rd_data; // @[NV_NVDLA_CSC_regfile.scala 155:43:@951.4]
  assign io_csb2csc_resp_valid = NV_NVDLA_CSB_LOGIC_io_csb2dp_resp_valid; // @[NV_NVDLA_CSC_regfile.scala 164:25:@958.4]
  assign io_csb2csc_resp_bits = NV_NVDLA_CSB_LOGIC_io_csb2dp_resp_bits; // @[NV_NVDLA_CSC_regfile.scala 164:25:@957.4]
  assign io_reg2dp_op_en = _T_147[2]; // @[NV_NVDLA_CSC_regfile.scala 135:21:@904.4]
  assign io_reg2dp_field_atomics = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_atomics : NV_NVDLA_CSC_dual_reg_io_field_atomics; // @[NV_NVDLA_CSC_regfile.scala 175:21:@1003.4]
  assign io_reg2dp_field_data_bank = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_data_bank : NV_NVDLA_CSC_dual_reg_io_field_data_bank; // @[NV_NVDLA_CSC_regfile.scala 175:21:@1002.4]
  assign io_reg2dp_field_weight_bank = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_weight_bank : NV_NVDLA_CSC_dual_reg_io_field_weight_bank; // @[NV_NVDLA_CSC_regfile.scala 175:21:@1001.4]
  assign io_reg2dp_field_conv_x_stride_ext = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_conv_x_stride_ext : NV_NVDLA_CSC_dual_reg_io_field_conv_x_stride_ext; // @[NV_NVDLA_CSC_regfile.scala 175:21:@999.4]
  assign io_reg2dp_field_conv_y_stride_ext = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_conv_y_stride_ext : NV_NVDLA_CSC_dual_reg_io_field_conv_y_stride_ext; // @[NV_NVDLA_CSC_regfile.scala 175:21:@998.4]
  assign io_reg2dp_field_datain_format = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_datain_format : NV_NVDLA_CSC_dual_reg_io_field_datain_format; // @[NV_NVDLA_CSC_regfile.scala 175:21:@996.4]
  assign io_reg2dp_field_datain_height_ext = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_datain_height_ext : NV_NVDLA_CSC_dual_reg_io_field_datain_height_ext; // @[NV_NVDLA_CSC_regfile.scala 175:21:@995.4]
  assign io_reg2dp_field_datain_width_ext = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_datain_width_ext : NV_NVDLA_CSC_dual_reg_io_field_datain_width_ext; // @[NV_NVDLA_CSC_regfile.scala 175:21:@994.4]
  assign io_reg2dp_field_datain_channel_ext = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_datain_channel_ext : NV_NVDLA_CSC_dual_reg_io_field_datain_channel_ext; // @[NV_NVDLA_CSC_regfile.scala 175:21:@993.4]
  assign io_reg2dp_field_dataout_height = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_dataout_height : NV_NVDLA_CSC_dual_reg_io_field_dataout_height; // @[NV_NVDLA_CSC_regfile.scala 175:21:@992.4]
  assign io_reg2dp_field_dataout_width = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_dataout_width : NV_NVDLA_CSC_dual_reg_io_field_dataout_width; // @[NV_NVDLA_CSC_regfile.scala 175:21:@991.4]
  assign io_reg2dp_field_x_dilation_ext = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_x_dilation_ext : NV_NVDLA_CSC_dual_reg_io_field_x_dilation_ext; // @[NV_NVDLA_CSC_regfile.scala 175:21:@989.4]
  assign io_reg2dp_field_y_dilation_ext = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_y_dilation_ext : NV_NVDLA_CSC_dual_reg_io_field_y_dilation_ext; // @[NV_NVDLA_CSC_regfile.scala 175:21:@988.4]
  assign io_reg2dp_field_entries = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_entries : NV_NVDLA_CSC_dual_reg_io_field_entries; // @[NV_NVDLA_CSC_regfile.scala 175:21:@987.4]
  assign io_reg2dp_field_conv_mode = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_conv_mode : NV_NVDLA_CSC_dual_reg_io_field_conv_mode; // @[NV_NVDLA_CSC_regfile.scala 175:21:@986.4]
  assign io_reg2dp_field_data_reuse = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_data_reuse : NV_NVDLA_CSC_dual_reg_io_field_data_reuse; // @[NV_NVDLA_CSC_regfile.scala 175:21:@985.4]
  assign io_reg2dp_field_skip_data_rls = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_skip_data_rls : NV_NVDLA_CSC_dual_reg_io_field_skip_data_rls; // @[NV_NVDLA_CSC_regfile.scala 175:21:@982.4]
  assign io_reg2dp_field_skip_weight_rls = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_skip_weight_rls : NV_NVDLA_CSC_dual_reg_io_field_skip_weight_rls; // @[NV_NVDLA_CSC_regfile.scala 175:21:@981.4]
  assign io_reg2dp_field_weight_reuse = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_weight_reuse : NV_NVDLA_CSC_dual_reg_io_field_weight_reuse; // @[NV_NVDLA_CSC_regfile.scala 175:21:@980.4]
  assign io_reg2dp_field_y_extension = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_y_extension : NV_NVDLA_CSC_dual_reg_io_field_y_extension; // @[NV_NVDLA_CSC_regfile.scala 175:21:@979.4]
  assign io_reg2dp_field_rls_slices = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_rls_slices : NV_NVDLA_CSC_dual_reg_io_field_rls_slices; // @[NV_NVDLA_CSC_regfile.scala 175:21:@977.4]
  assign io_reg2dp_field_weight_bytes = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_weight_bytes : NV_NVDLA_CSC_dual_reg_io_field_weight_bytes; // @[NV_NVDLA_CSC_regfile.scala 175:21:@976.4]
  assign io_reg2dp_field_weight_format = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_weight_format : NV_NVDLA_CSC_dual_reg_io_field_weight_format; // @[NV_NVDLA_CSC_regfile.scala 175:21:@975.4]
  assign io_reg2dp_field_weight_height_ext = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_weight_height_ext : NV_NVDLA_CSC_dual_reg_io_field_weight_height_ext; // @[NV_NVDLA_CSC_regfile.scala 175:21:@974.4]
  assign io_reg2dp_field_weight_width_ext = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_weight_width_ext : NV_NVDLA_CSC_dual_reg_io_field_weight_width_ext; // @[NV_NVDLA_CSC_regfile.scala 175:21:@973.4]
  assign io_reg2dp_field_weight_channel_ext = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_weight_channel_ext : NV_NVDLA_CSC_dual_reg_io_field_weight_channel_ext; // @[NV_NVDLA_CSC_regfile.scala 175:21:@972.4]
  assign io_reg2dp_field_weight_kernel = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_weight_kernel : NV_NVDLA_CSC_dual_reg_io_field_weight_kernel; // @[NV_NVDLA_CSC_regfile.scala 175:21:@971.4]
  assign io_reg2dp_field_wmb_bytes = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_wmb_bytes : NV_NVDLA_CSC_dual_reg_io_field_wmb_bytes; // @[NV_NVDLA_CSC_regfile.scala 175:21:@970.4]
  assign io_reg2dp_field_pad_left = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_pad_left : NV_NVDLA_CSC_dual_reg_io_field_pad_left; // @[NV_NVDLA_CSC_regfile.scala 175:21:@969.4]
  assign io_reg2dp_field_pad_top = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_pad_top : NV_NVDLA_CSC_dual_reg_io_field_pad_top; // @[NV_NVDLA_CSC_regfile.scala 175:21:@968.4]
  assign io_reg2dp_field_pad_value = _T_105 ? NV_NVDLA_CSC_dual_reg_1_io_field_pad_value : NV_NVDLA_CSC_dual_reg_io_field_pad_value; // @[NV_NVDLA_CSC_regfile.scala 175:21:@967.4]
  assign NV_NVDLA_BASIC_REG_single_reset = reset; // @[:@839.4]
  assign NV_NVDLA_BASIC_REG_single_io_nvdla_core_clk = io_nvdla_core_clk; // @[NV_NVDLA_CSC_regfile.scala 60:36:@840.4]
  assign NV_NVDLA_BASIC_REG_single_io_reg_offset = NV_NVDLA_CSB_LOGIC_io_reg_offset; // @[NV_NVDLA_CSC_regfile.scala 61:32:@841.4]
  assign NV_NVDLA_BASIC_REG_single_io_reg_wr_data = NV_NVDLA_CSB_LOGIC_io_reg_wr_data; // @[NV_NVDLA_CSC_regfile.scala 62:33:@842.4]
  assign NV_NVDLA_BASIC_REG_single_io_reg_wr_en = _T_184 & _T_187; // @[NV_NVDLA_CSC_regfile.scala 63:31:@843.4]
  assign NV_NVDLA_BASIC_REG_single_io_consumer = _T_105; // @[NV_NVDLA_CSC_regfile.scala 65:30:@844.4]
  assign NV_NVDLA_BASIC_REG_single_io_status_0 = _T_128 ? 2'h0 : _T_134; // @[NV_NVDLA_CSC_regfile.scala 66:30:@845.4]
  assign NV_NVDLA_BASIC_REG_single_io_status_1 = _T_137 ? 2'h0 : _T_143; // @[NV_NVDLA_CSC_regfile.scala 67:30:@846.4]
  assign NV_NVDLA_CSC_dual_reg_reset = reset; // @[:@851.4]
  assign NV_NVDLA_CSC_dual_reg_io_nvdla_core_clk = io_nvdla_core_clk; // @[NV_NVDLA_CSC_regfile.scala 75:37:@852.4]
  assign NV_NVDLA_CSC_dual_reg_io_reg_offset = NV_NVDLA_CSB_LOGIC_io_reg_offset; // @[NV_NVDLA_CSC_regfile.scala 76:33:@853.4]
  assign NV_NVDLA_CSC_dual_reg_io_reg_wr_data = NV_NVDLA_CSB_LOGIC_io_reg_wr_data; // @[NV_NVDLA_CSC_regfile.scala 77:34:@854.4]
  assign NV_NVDLA_CSC_dual_reg_io_reg_wr_en = _T_204 & _T_128; // @[NV_NVDLA_CSC_regfile.scala 78:32:@855.4]
  assign NV_NVDLA_CSC_dual_reg_io_op_en = _T_120; // @[NV_NVDLA_CSC_regfile.scala 80:28:@856.4]
  assign NV_NVDLA_CSC_dual_reg_1_reset = reset; // @[:@861.4]
  assign NV_NVDLA_CSC_dual_reg_1_io_nvdla_core_clk = io_nvdla_core_clk; // @[NV_NVDLA_CSC_regfile.scala 88:37:@862.4]
  assign NV_NVDLA_CSC_dual_reg_1_io_reg_offset = NV_NVDLA_CSB_LOGIC_io_reg_offset; // @[NV_NVDLA_CSC_regfile.scala 89:33:@863.4]
  assign NV_NVDLA_CSC_dual_reg_1_io_reg_wr_data = NV_NVDLA_CSB_LOGIC_io_reg_wr_data; // @[NV_NVDLA_CSC_regfile.scala 90:34:@864.4]
  assign NV_NVDLA_CSC_dual_reg_1_io_reg_wr_en = _T_208 & _T_137; // @[NV_NVDLA_CSC_regfile.scala 91:32:@865.4]
  assign NV_NVDLA_CSC_dual_reg_1_io_op_en = _T_125; // @[NV_NVDLA_CSC_regfile.scala 93:28:@866.4]
  assign NV_NVDLA_CSB_LOGIC_reset = reset; // @[:@955.4]
  assign NV_NVDLA_CSB_LOGIC_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CSC_regfile.scala 163:22:@956.4]
  assign NV_NVDLA_CSB_LOGIC_io_csb2dp_req_valid = io_csb2csc_req_valid; // @[NV_NVDLA_CSC_regfile.scala 164:25:@960.4]
  assign NV_NVDLA_CSB_LOGIC_io_csb2dp_req_bits = io_csb2csc_req_bits; // @[NV_NVDLA_CSC_regfile.scala 164:25:@959.4]
  assign NV_NVDLA_CSB_LOGIC_io_reg_rd_data = _T_222 | _T_227; // @[NV_NVDLA_CSC_regfile.scala 168:30:@965.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_105 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_120 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_125 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_147 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_105 <= 1'h0;
    end else begin
      if (io_dp2reg_done) begin
        _T_105 <= _T_126;
      end
    end
    if (reset) begin
      _T_120 <= 1'h0;
    end else begin
      if (_T_149) begin
        _T_120 <= _T_150;
      end else begin
        if (_T_153) begin
          _T_120 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      if (_T_158) begin
        _T_125 <= _T_150;
      end else begin
        if (_T_162) begin
          _T_125 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_147 <= 3'h0;
    end else begin
      if (io_dp2reg_done) begin
        _T_147 <= 3'h0;
      end else begin
        _T_147 <= _T_169;
      end
    end
  end
endmodule
module nv_ram_rwsp( // @[:@1036.2]
  input         io_clk, // @[:@1039.4]
  input         io_re, // @[:@1039.4]
  input         io_we, // @[:@1039.4]
  input         io_ore, // @[:@1039.4]
  input  [1:0]  io_ra, // @[:@1039.4]
  input  [1:0]  io_wa, // @[:@1039.4]
  input  [32:0] io_di, // @[:@1039.4]
  output [32:0] io_dout // @[:@1039.4]
);
  reg [32:0] _T_26_0; // @[nv_ram_rwsp.scala 31:18:@1041.4]
  reg [63:0] _RAND_0;
  reg [32:0] _T_26_1; // @[nv_ram_rwsp.scala 31:18:@1041.4]
  reg [63:0] _RAND_1;
  reg [32:0] _T_26_2; // @[nv_ram_rwsp.scala 31:18:@1041.4]
  reg [63:0] _RAND_2;
  reg [32:0] _T_26_3; // @[nv_ram_rwsp.scala 31:18:@1041.4]
  reg [63:0] _RAND_3;
  reg [1:0] _T_34; // @[nv_ram_rwsp.scala 32:19:@1042.4]
  reg [31:0] _RAND_4;
  reg [32:0] _T_36; // @[nv_ram_rwsp.scala 33:21:@1043.4]
  reg [63:0] _RAND_5;
  wire [32:0] _GEN_0; // @[nv_ram_rwsp.scala 36:20:@1045.6]
  wire [32:0] _GEN_1; // @[nv_ram_rwsp.scala 36:20:@1045.6]
  wire [32:0] _GEN_2; // @[nv_ram_rwsp.scala 36:20:@1045.6]
  wire [32:0] _GEN_3; // @[nv_ram_rwsp.scala 36:20:@1045.6]
  wire [32:0] _GEN_10; // @[nv_ram_rwsp.scala 43:16:@1051.6]
  wire [32:0] _GEN_11; // @[nv_ram_rwsp.scala 43:16:@1051.6]
  wire [32:0] _GEN_12; // @[nv_ram_rwsp.scala 43:16:@1051.6]
  assign _GEN_0 = 2'h0 == io_wa ? io_di : _T_26_0; // @[nv_ram_rwsp.scala 36:20:@1045.6]
  assign _GEN_1 = 2'h1 == io_wa ? io_di : _T_26_1; // @[nv_ram_rwsp.scala 36:20:@1045.6]
  assign _GEN_2 = 2'h2 == io_wa ? io_di : _T_26_2; // @[nv_ram_rwsp.scala 36:20:@1045.6]
  assign _GEN_3 = 2'h3 == io_wa ? io_di : _T_26_3; // @[nv_ram_rwsp.scala 36:20:@1045.6]
  assign _GEN_10 = 2'h1 == _T_34 ? _T_26_1 : _T_26_0; // @[nv_ram_rwsp.scala 43:16:@1051.6]
  assign _GEN_11 = 2'h2 == _T_34 ? _T_26_2 : _GEN_10; // @[nv_ram_rwsp.scala 43:16:@1051.6]
  assign _GEN_12 = 2'h3 == _T_34 ? _T_26_3 : _GEN_11; // @[nv_ram_rwsp.scala 43:16:@1051.6]
  assign io_dout = _T_36; // @[nv_ram_rwsp.scala 45:13:@1053.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_26_0 = _RAND_0[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  _T_26_1 = _RAND_1[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  _T_26_2 = _RAND_2[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  _T_26_3 = _RAND_3[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_34 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  _T_36 = _RAND_5[32:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_clk) begin
    if (io_we) begin
      if (2'h0 == io_wa) begin
        _T_26_0 <= io_di;
      end
    end
    if (io_we) begin
      if (2'h1 == io_wa) begin
        _T_26_1 <= io_di;
      end
    end
    if (io_we) begin
      if (2'h2 == io_wa) begin
        _T_26_2 <= io_di;
      end
    end
    if (io_we) begin
      if (2'h3 == io_wa) begin
        _T_26_3 <= io_di;
      end
    end
    if (io_re) begin
      _T_34 <= io_ra;
    end
    if (io_ore) begin
      if (2'h3 == _T_34) begin
        _T_36 <= _T_26_3;
      end else begin
        if (2'h2 == _T_34) begin
          _T_36 <= _T_26_2;
        end else begin
          if (2'h1 == _T_34) begin
            _T_36 <= _T_26_1;
          end else begin
            _T_36 <= _T_26_0;
          end
        end
      end
    end
  end
endmodule
module NV_NVDLA_fifo( // @[:@1055.2]
  input         clock, // @[:@1056.4]
  input         reset, // @[:@1057.4]
  input         io_clk, // @[:@1058.4]
  input         io_wr_pvld, // @[:@1058.4]
  output        io_wr_prdy, // @[:@1058.4]
  input  [32:0] io_wr_pd, // @[:@1058.4]
  output        io_wr_empty, // @[:@1058.4]
  output        io_rd_pvld, // @[:@1058.4]
  input         io_rd_prdy, // @[:@1058.4]
  output [32:0] io_rd_pd // @[:@1058.4]
);
  wire  nv_ram_rwsp_io_clk; // @[FIFO.scala 270:29:@1138.4]
  wire  nv_ram_rwsp_io_re; // @[FIFO.scala 270:29:@1138.4]
  wire  nv_ram_rwsp_io_we; // @[FIFO.scala 270:29:@1138.4]
  wire  nv_ram_rwsp_io_ore; // @[FIFO.scala 270:29:@1138.4]
  wire [1:0] nv_ram_rwsp_io_ra; // @[FIFO.scala 270:29:@1138.4]
  wire [1:0] nv_ram_rwsp_io_wa; // @[FIFO.scala 270:29:@1138.4]
  wire [32:0] nv_ram_rwsp_io_di; // @[FIFO.scala 270:29:@1138.4]
  wire [32:0] nv_ram_rwsp_io_dout; // @[FIFO.scala 270:29:@1138.4]
  reg  _T_28; // @[FIFO.scala 156:56:@1067.4]
  reg [31:0] _RAND_0;
  reg  _T_31; // @[FIFO.scala 158:52:@1068.4]
  reg [31:0] _RAND_1;
  reg [32:0] _T_33; // @[FIFO.scala 159:64:@1069.4]
  reg [63:0] _RAND_2;
  reg  _T_36; // @[FIFO.scala 160:52:@1070.4]
  reg [31:0] _RAND_3;
  wire  _T_135; // @[FIFO.scala 331:38:@1169.4]
  wire  _T_56; // @[FIFO.scala 183:39:@1091.4]
  wire  _T_57; // @[FIFO.scala 183:36:@1092.4]
  reg [2:0] _T_62; // @[FIFO.scala 186:53:@1095.4]
  reg [31:0] _RAND_4;
  wire [3:0] _T_69; // @[FIFO.scala 191:69:@1100.4]
  wire [2:0] _T_70; // @[FIFO.scala 191:69:@1101.4]
  wire [2:0] _T_71; // @[FIFO.scala 191:46:@1102.4]
  wire  _T_74; // @[FIFO.scala 194:80:@1104.4]
  wire  _T_76; // @[FIFO.scala 195:40:@1105.4]
  wire [3:0] _T_64; // @[FIFO.scala 190:76:@1096.4]
  wire [3:0] _T_65; // @[FIFO.scala 190:76:@1097.4]
  wire [2:0] _T_66; // @[FIFO.scala 190:76:@1098.4]
  wire [2:0] _T_67; // @[FIFO.scala 190:43:@1099.4]
  wire [2:0] _T_72; // @[FIFO.scala 192:32:@1103.4]
  wire  _T_39; // @[FIFO.scala 166:60:@1072.4]
  wire  _T_41; // @[FIFO.scala 166:80:@1073.4]
  wire  _T_42; // @[FIFO.scala 166:77:@1074.4]
  wire  _T_43; // @[FIFO.scala 167:38:@1075.4]
  wire  _T_44; // @[FIFO.scala 168:45:@1076.4]
  wire  _T_46; // @[FIFO.scala 171:18:@1078.4]
  wire  _T_48; // @[FIFO.scala 172:45:@1080.6]
  wire  _T_49; // @[FIFO.scala 172:42:@1081.6]
  wire  _GEN_0; // @[FIFO.scala 171:34:@1079.4]
  wire  _T_52; // @[FIFO.scala 176:34:@1085.4]
  wire  _T_84; // @[FIFO.scala 202:27:@1113.4]
  wire [2:0] _GEN_2; // @[FIFO.scala 202:40:@1114.4]
  wire  _T_86; // @[FIFO.scala 207:54:@1117.4]
  wire  _T_88; // @[FIFO.scala 207:65:@1118.4]
  wire  _T_89; // @[FIFO.scala 207:62:@1119.4]
  reg  _T_92; // @[FIFO.scala 207:39:@1120.4]
  reg [31:0] _RAND_5;
  reg [1:0] _T_95; // @[FIFO.scala 215:68:@1123.4]
  reg [31:0] _RAND_6;
  wire [2:0] _T_97; // @[FIFO.scala 217:42:@1124.4]
  wire [1:0] _T_98; // @[FIFO.scala 217:42:@1125.4]
  wire [1:0] _GEN_3; // @[FIFO.scala 218:29:@1126.4]
  reg [1:0] _T_103; // @[FIFO.scala 224:63:@1130.4]
  reg [31:0] _RAND_7;
  wire [2:0] _T_105; // @[FIFO.scala 225:42:@1131.4]
  wire [1:0] _T_106; // @[FIFO.scala 225:42:@1132.4]
  wire [1:0] _GEN_4; // @[FIFO.scala 227:29:@1133.4]
  reg  _T_114; // @[FIFO.scala 289:73:@1152.4]
  reg [31:0] _RAND_8;
  reg  _T_117; // @[FIFO.scala 295:72:@1154.4]
  reg [31:0] _RAND_9;
  reg  _T_120; // @[FIFO.scala 297:97:@1155.4]
  reg [31:0] _RAND_10;
  reg [2:0] _T_123; // @[FIFO.scala 299:53:@1156.4]
  reg [31:0] _RAND_11;
  wire [3:0] _T_125; // @[FIFO.scala 300:74:@1157.4]
  wire [3:0] _T_126; // @[FIFO.scala 300:74:@1158.4]
  wire [2:0] _T_127; // @[FIFO.scala 300:74:@1159.4]
  wire [2:0] _T_128; // @[FIFO.scala 300:43:@1160.4]
  wire [3:0] _T_130; // @[FIFO.scala 301:68:@1161.4]
  wire [2:0] _T_131; // @[FIFO.scala 301:68:@1162.4]
  wire [2:0] _T_132; // @[FIFO.scala 301:46:@1163.4]
  wire [2:0] _T_133; // @[FIFO.scala 302:32:@1164.4]
  wire  _T_134; // @[FIFO.scala 303:25:@1165.4]
  wire [2:0] _GEN_5; // @[FIFO.scala 303:39:@1166.4]
  wire  _T_137; // @[FIFO.scala 333:77:@1171.4]
  wire  _T_139; // @[FIFO.scala 334:83:@1172.4]
  wire  _T_140; // @[FIFO.scala 335:44:@1173.4]
  wire  _T_141; // @[FIFO.scala 336:60:@1174.4]
  wire  _T_143; // @[FIFO.scala 336:81:@1176.4]
  wire  _GEN_6; // @[FIFO.scala 338:43:@1180.4]
  wire  _T_147; // @[FIFO.scala 341:66:@1183.4]
  wire  _T_148; // @[FIFO.scala 341:63:@1184.4]
  wire  _T_149; // @[FIFO.scala 341:43:@1185.4]
  nv_ram_rwsp nv_ram_rwsp ( // @[FIFO.scala 270:29:@1138.4]
    .io_clk(nv_ram_rwsp_io_clk),
    .io_re(nv_ram_rwsp_io_re),
    .io_we(nv_ram_rwsp_io_we),
    .io_ore(nv_ram_rwsp_io_ore),
    .io_ra(nv_ram_rwsp_io_ra),
    .io_wa(nv_ram_rwsp_io_wa),
    .io_di(nv_ram_rwsp_io_di),
    .io_dout(nv_ram_rwsp_io_dout)
  );
  assign _T_135 = io_rd_pvld & io_rd_prdy; // @[FIFO.scala 331:38:@1169.4]
  assign _T_56 = _T_28 == 1'h0; // @[FIFO.scala 183:39:@1091.4]
  assign _T_57 = _T_31 & _T_56; // @[FIFO.scala 183:36:@1092.4]
  assign _T_69 = _T_62 + 3'h1; // @[FIFO.scala 191:69:@1100.4]
  assign _T_70 = _T_62 + 3'h1; // @[FIFO.scala 191:69:@1101.4]
  assign _T_71 = _T_57 ? _T_70 : _T_62; // @[FIFO.scala 191:46:@1102.4]
  assign _T_74 = _T_71 == 3'h4; // @[FIFO.scala 194:80:@1104.4]
  assign _T_76 = _T_135 ? 1'h0 : _T_74; // @[FIFO.scala 195:40:@1105.4]
  assign _T_64 = _T_62 - 3'h1; // @[FIFO.scala 190:76:@1096.4]
  assign _T_65 = $unsigned(_T_64); // @[FIFO.scala 190:76:@1097.4]
  assign _T_66 = _T_65[2:0]; // @[FIFO.scala 190:76:@1098.4]
  assign _T_67 = _T_57 ? _T_62 : _T_66; // @[FIFO.scala 190:43:@1099.4]
  assign _T_72 = _T_135 ? _T_67 : _T_71; // @[FIFO.scala 192:32:@1103.4]
  assign _T_39 = _T_31 & _T_76; // @[FIFO.scala 166:60:@1072.4]
  assign _T_41 = _T_57 == 1'h0; // @[FIFO.scala 166:80:@1073.4]
  assign _T_42 = _T_39 & _T_41; // @[FIFO.scala 166:77:@1074.4]
  assign _T_43 = io_wr_pvld ? _T_76 : _T_42; // @[FIFO.scala 167:38:@1075.4]
  assign _T_44 = _T_31 & _T_28; // @[FIFO.scala 168:45:@1076.4]
  assign _T_46 = _T_44 == 1'h0; // @[FIFO.scala 171:18:@1078.4]
  assign _T_48 = _T_36 == 1'h0; // @[FIFO.scala 172:45:@1080.6]
  assign _T_49 = io_wr_pvld & _T_48; // @[FIFO.scala 172:42:@1081.6]
  assign _GEN_0 = _T_46 ? _T_49 : _T_31; // @[FIFO.scala 171:34:@1079.4]
  assign _T_52 = _T_48 & io_wr_pvld; // @[FIFO.scala 176:34:@1085.4]
  assign _T_84 = _T_57 ^ _T_135; // @[FIFO.scala 202:27:@1113.4]
  assign _GEN_2 = _T_84 ? _T_72 : _T_62; // @[FIFO.scala 202:40:@1114.4]
  assign _T_86 = _T_72 == 3'h0; // @[FIFO.scala 207:54:@1117.4]
  assign _T_88 = io_wr_pvld == 1'h0; // @[FIFO.scala 207:65:@1118.4]
  assign _T_89 = _T_86 & _T_88; // @[FIFO.scala 207:62:@1119.4]
  assign _T_97 = _T_95 + 2'h1; // @[FIFO.scala 217:42:@1124.4]
  assign _T_98 = _T_95 + 2'h1; // @[FIFO.scala 217:42:@1125.4]
  assign _GEN_3 = _T_57 ? _T_98 : _T_95; // @[FIFO.scala 218:29:@1126.4]
  assign _T_105 = _T_103 + 2'h1; // @[FIFO.scala 225:42:@1131.4]
  assign _T_106 = _T_103 + 2'h1; // @[FIFO.scala 225:42:@1132.4]
  assign _GEN_4 = _T_135 ? _T_106 : _T_103; // @[FIFO.scala 227:29:@1133.4]
  assign _T_125 = _T_123 - 3'h1; // @[FIFO.scala 300:74:@1157.4]
  assign _T_126 = $unsigned(_T_125); // @[FIFO.scala 300:74:@1158.4]
  assign _T_127 = _T_126[2:0]; // @[FIFO.scala 300:74:@1159.4]
  assign _T_128 = _T_114 ? _T_123 : _T_127; // @[FIFO.scala 300:43:@1160.4]
  assign _T_130 = _T_123 + 3'h1; // @[FIFO.scala 301:68:@1161.4]
  assign _T_131 = _T_123 + 3'h1; // @[FIFO.scala 301:68:@1162.4]
  assign _T_132 = _T_114 ? _T_131 : _T_123; // @[FIFO.scala 301:46:@1163.4]
  assign _T_133 = _T_135 ? _T_128 : _T_132; // @[FIFO.scala 302:32:@1164.4]
  assign _T_134 = _T_114 | _T_135; // @[FIFO.scala 303:25:@1165.4]
  assign _GEN_5 = _T_134 ? _T_133 : _T_123; // @[FIFO.scala 303:39:@1166.4]
  assign _T_137 = _T_128 != 3'h0; // @[FIFO.scala 333:77:@1171.4]
  assign _T_139 = _T_132 != 3'h0; // @[FIFO.scala 334:83:@1172.4]
  assign _T_140 = _T_135 ? _T_137 : _T_139; // @[FIFO.scala 335:44:@1173.4]
  assign _T_141 = ~ _T_117; // @[FIFO.scala 336:60:@1174.4]
  assign _T_143 = _T_141 | _T_135; // @[FIFO.scala 336:81:@1176.4]
  assign _GEN_6 = _T_134 ? _T_140 : _T_117; // @[FIFO.scala 338:43:@1180.4]
  assign _T_147 = io_rd_prdy == 1'h0; // @[FIFO.scala 341:66:@1183.4]
  assign _T_148 = _T_120 & _T_147; // @[FIFO.scala 341:63:@1184.4]
  assign _T_149 = _T_117 | _T_148; // @[FIFO.scala 341:43:@1185.4]
  assign io_wr_prdy = _T_36 == 1'h0; // @[FIFO.scala 182:20:@1090.4]
  assign io_wr_empty = _T_92; // @[FIFO.scala 207:29:@1122.4]
  assign io_rd_pvld = _T_120; // @[FIFO.scala 344:24:@1187.4]
  assign io_rd_pd = nv_ram_rwsp_io_dout; // @[FIFO.scala 345:22:@1188.4]
  assign nv_ram_rwsp_io_clk = io_clk; // @[FIFO.scala 271:24:@1141.4]
  assign nv_ram_rwsp_io_re = _T_140 & _T_143; // @[FIFO.scala 279:23:@1148.4]
  assign nv_ram_rwsp_io_we = _T_31 & _T_56; // @[FIFO.scala 276:23:@1144.4]
  assign nv_ram_rwsp_io_ore = io_rd_pvld & io_rd_prdy; // @[FIFO.scala 280:24:@1149.4]
  assign nv_ram_rwsp_io_ra = _T_135 ? _T_106 : _T_103; // @[FIFO.scala 278:23:@1147.4]
  assign nv_ram_rwsp_io_wa = _T_95; // @[FIFO.scala 274:27:@1143.4]
  assign nv_ram_rwsp_io_di = _T_33; // @[FIFO.scala 277:23:@1145.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_28 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_31 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  _T_33 = _RAND_2[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_36 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_62 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_92 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_95 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_103 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_114 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_117 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_120 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_123 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_135) begin
        _T_28 <= 1'h0;
      end else begin
        _T_28 <= _T_74;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_46) begin
        _T_31 <= _T_49;
      end
    end
    if (_T_52) begin
      _T_33 <= io_wr_pd;
    end
    if (reset) begin
      _T_36 <= 1'h0;
    end else begin
      if (io_wr_pvld) begin
        if (_T_135) begin
          _T_36 <= 1'h0;
        end else begin
          _T_36 <= _T_74;
        end
      end else begin
        _T_36 <= _T_42;
      end
    end
    if (reset) begin
      _T_62 <= 3'h0;
    end else begin
      if (_T_84) begin
        if (_T_135) begin
          if (!(_T_57)) begin
            _T_62 <= _T_66;
          end
        end else begin
          if (_T_57) begin
            _T_62 <= _T_70;
          end
        end
      end
    end
    if (reset) begin
      _T_92 <= 1'h1;
    end else begin
      _T_92 <= _T_89;
    end
    if (reset) begin
      _T_95 <= 2'h0;
    end else begin
      if (_T_57) begin
        _T_95 <= _T_98;
      end
    end
    if (reset) begin
      _T_103 <= 2'h0;
    end else begin
      if (_T_135) begin
        _T_103 <= _T_106;
      end
    end
    if (reset) begin
      _T_114 <= 1'h0;
    end else begin
      _T_114 <= _T_57;
    end
    if (reset) begin
      _T_117 <= 1'h0;
    end else begin
      if (_T_134) begin
        if (_T_135) begin
          _T_117 <= _T_137;
        end else begin
          _T_117 <= _T_139;
        end
      end
    end
    if (reset) begin
      _T_120 <= 1'h0;
    end else begin
      _T_120 <= _T_149;
    end
    if (reset) begin
      _T_123 <= 3'h0;
    end else begin
      if (_T_134) begin
        if (_T_135) begin
          if (!(_T_114)) begin
            _T_123 <= _T_127;
          end
        end else begin
          if (_T_114) begin
            _T_123 <= _T_131;
          end
        end
      end
    end
  end
endmodule
module nv_ram_rwsp_1( // @[:@1235.2]
  input         io_clk, // @[:@1238.4]
  input         io_re, // @[:@1238.4]
  input         io_we, // @[:@1238.4]
  input         io_ore, // @[:@1238.4]
  input  [1:0]  io_ra, // @[:@1238.4]
  input  [1:0]  io_wa, // @[:@1238.4]
  input  [19:0] io_di, // @[:@1238.4]
  output [19:0] io_dout // @[:@1238.4]
);
  reg [19:0] _T_26_0; // @[nv_ram_rwsp.scala 31:18:@1240.4]
  reg [31:0] _RAND_0;
  reg [19:0] _T_26_1; // @[nv_ram_rwsp.scala 31:18:@1240.4]
  reg [31:0] _RAND_1;
  reg [19:0] _T_26_2; // @[nv_ram_rwsp.scala 31:18:@1240.4]
  reg [31:0] _RAND_2;
  reg [19:0] _T_26_3; // @[nv_ram_rwsp.scala 31:18:@1240.4]
  reg [31:0] _RAND_3;
  reg [1:0] _T_34; // @[nv_ram_rwsp.scala 32:19:@1241.4]
  reg [31:0] _RAND_4;
  reg [19:0] _T_36; // @[nv_ram_rwsp.scala 33:21:@1242.4]
  reg [31:0] _RAND_5;
  wire [19:0] _GEN_0; // @[nv_ram_rwsp.scala 36:20:@1244.6]
  wire [19:0] _GEN_1; // @[nv_ram_rwsp.scala 36:20:@1244.6]
  wire [19:0] _GEN_2; // @[nv_ram_rwsp.scala 36:20:@1244.6]
  wire [19:0] _GEN_3; // @[nv_ram_rwsp.scala 36:20:@1244.6]
  wire [19:0] _GEN_10; // @[nv_ram_rwsp.scala 43:16:@1250.6]
  wire [19:0] _GEN_11; // @[nv_ram_rwsp.scala 43:16:@1250.6]
  wire [19:0] _GEN_12; // @[nv_ram_rwsp.scala 43:16:@1250.6]
  assign _GEN_0 = 2'h0 == io_wa ? io_di : _T_26_0; // @[nv_ram_rwsp.scala 36:20:@1244.6]
  assign _GEN_1 = 2'h1 == io_wa ? io_di : _T_26_1; // @[nv_ram_rwsp.scala 36:20:@1244.6]
  assign _GEN_2 = 2'h2 == io_wa ? io_di : _T_26_2; // @[nv_ram_rwsp.scala 36:20:@1244.6]
  assign _GEN_3 = 2'h3 == io_wa ? io_di : _T_26_3; // @[nv_ram_rwsp.scala 36:20:@1244.6]
  assign _GEN_10 = 2'h1 == _T_34 ? _T_26_1 : _T_26_0; // @[nv_ram_rwsp.scala 43:16:@1250.6]
  assign _GEN_11 = 2'h2 == _T_34 ? _T_26_2 : _GEN_10; // @[nv_ram_rwsp.scala 43:16:@1250.6]
  assign _GEN_12 = 2'h3 == _T_34 ? _T_26_3 : _GEN_11; // @[nv_ram_rwsp.scala 43:16:@1250.6]
  assign io_dout = _T_36; // @[nv_ram_rwsp.scala 45:13:@1252.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_26_0 = _RAND_0[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26_1 = _RAND_1[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_26_2 = _RAND_2[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_26_3 = _RAND_3[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_34 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_36 = _RAND_5[19:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_clk) begin
    if (io_we) begin
      if (2'h0 == io_wa) begin
        _T_26_0 <= io_di;
      end
    end
    if (io_we) begin
      if (2'h1 == io_wa) begin
        _T_26_1 <= io_di;
      end
    end
    if (io_we) begin
      if (2'h2 == io_wa) begin
        _T_26_2 <= io_di;
      end
    end
    if (io_we) begin
      if (2'h3 == io_wa) begin
        _T_26_3 <= io_di;
      end
    end
    if (io_re) begin
      _T_34 <= io_ra;
    end
    if (io_ore) begin
      if (2'h3 == _T_34) begin
        _T_36 <= _T_26_3;
      end else begin
        if (2'h2 == _T_34) begin
          _T_36 <= _T_26_2;
        end else begin
          if (2'h1 == _T_34) begin
            _T_36 <= _T_26_1;
          end else begin
            _T_36 <= _T_26_0;
          end
        end
      end
    end
  end
endmodule
module NV_NVDLA_fifo_1( // @[:@1254.2]
  input         clock, // @[:@1255.4]
  input         reset, // @[:@1256.4]
  input         io_clk, // @[:@1257.4]
  input         io_wr_pvld, // @[:@1257.4]
  output        io_wr_prdy, // @[:@1257.4]
  input  [19:0] io_wr_pd, // @[:@1257.4]
  output        io_wr_empty, // @[:@1257.4]
  output        io_rd_pvld, // @[:@1257.4]
  input         io_rd_prdy, // @[:@1257.4]
  output [19:0] io_rd_pd // @[:@1257.4]
);
  wire  nv_ram_rwsp_io_clk; // @[FIFO.scala 270:29:@1337.4]
  wire  nv_ram_rwsp_io_re; // @[FIFO.scala 270:29:@1337.4]
  wire  nv_ram_rwsp_io_we; // @[FIFO.scala 270:29:@1337.4]
  wire  nv_ram_rwsp_io_ore; // @[FIFO.scala 270:29:@1337.4]
  wire [1:0] nv_ram_rwsp_io_ra; // @[FIFO.scala 270:29:@1337.4]
  wire [1:0] nv_ram_rwsp_io_wa; // @[FIFO.scala 270:29:@1337.4]
  wire [19:0] nv_ram_rwsp_io_di; // @[FIFO.scala 270:29:@1337.4]
  wire [19:0] nv_ram_rwsp_io_dout; // @[FIFO.scala 270:29:@1337.4]
  reg  _T_28; // @[FIFO.scala 156:56:@1266.4]
  reg [31:0] _RAND_0;
  reg  _T_31; // @[FIFO.scala 158:52:@1267.4]
  reg [31:0] _RAND_1;
  reg [19:0] _T_33; // @[FIFO.scala 159:64:@1268.4]
  reg [31:0] _RAND_2;
  reg  _T_36; // @[FIFO.scala 160:52:@1269.4]
  reg [31:0] _RAND_3;
  wire  _T_135; // @[FIFO.scala 331:38:@1368.4]
  wire  _T_56; // @[FIFO.scala 183:39:@1290.4]
  wire  _T_57; // @[FIFO.scala 183:36:@1291.4]
  reg [2:0] _T_62; // @[FIFO.scala 186:53:@1294.4]
  reg [31:0] _RAND_4;
  wire [3:0] _T_69; // @[FIFO.scala 191:69:@1299.4]
  wire [2:0] _T_70; // @[FIFO.scala 191:69:@1300.4]
  wire [2:0] _T_71; // @[FIFO.scala 191:46:@1301.4]
  wire  _T_74; // @[FIFO.scala 194:80:@1303.4]
  wire  _T_76; // @[FIFO.scala 195:40:@1304.4]
  wire [3:0] _T_64; // @[FIFO.scala 190:76:@1295.4]
  wire [3:0] _T_65; // @[FIFO.scala 190:76:@1296.4]
  wire [2:0] _T_66; // @[FIFO.scala 190:76:@1297.4]
  wire [2:0] _T_67; // @[FIFO.scala 190:43:@1298.4]
  wire [2:0] _T_72; // @[FIFO.scala 192:32:@1302.4]
  wire  _T_39; // @[FIFO.scala 166:60:@1271.4]
  wire  _T_41; // @[FIFO.scala 166:80:@1272.4]
  wire  _T_42; // @[FIFO.scala 166:77:@1273.4]
  wire  _T_43; // @[FIFO.scala 167:38:@1274.4]
  wire  _T_44; // @[FIFO.scala 168:45:@1275.4]
  wire  _T_46; // @[FIFO.scala 171:18:@1277.4]
  wire  _T_48; // @[FIFO.scala 172:45:@1279.6]
  wire  _T_49; // @[FIFO.scala 172:42:@1280.6]
  wire  _GEN_0; // @[FIFO.scala 171:34:@1278.4]
  wire  _T_52; // @[FIFO.scala 176:34:@1284.4]
  wire  _T_84; // @[FIFO.scala 202:27:@1312.4]
  wire [2:0] _GEN_2; // @[FIFO.scala 202:40:@1313.4]
  wire  _T_86; // @[FIFO.scala 207:54:@1316.4]
  wire  _T_88; // @[FIFO.scala 207:65:@1317.4]
  wire  _T_89; // @[FIFO.scala 207:62:@1318.4]
  reg  _T_92; // @[FIFO.scala 207:39:@1319.4]
  reg [31:0] _RAND_5;
  reg [1:0] _T_95; // @[FIFO.scala 215:68:@1322.4]
  reg [31:0] _RAND_6;
  wire [2:0] _T_97; // @[FIFO.scala 217:42:@1323.4]
  wire [1:0] _T_98; // @[FIFO.scala 217:42:@1324.4]
  wire [1:0] _GEN_3; // @[FIFO.scala 218:29:@1325.4]
  reg [1:0] _T_103; // @[FIFO.scala 224:63:@1329.4]
  reg [31:0] _RAND_7;
  wire [2:0] _T_105; // @[FIFO.scala 225:42:@1330.4]
  wire [1:0] _T_106; // @[FIFO.scala 225:42:@1331.4]
  wire [1:0] _GEN_4; // @[FIFO.scala 227:29:@1332.4]
  reg  _T_114; // @[FIFO.scala 289:73:@1351.4]
  reg [31:0] _RAND_8;
  reg  _T_117; // @[FIFO.scala 295:72:@1353.4]
  reg [31:0] _RAND_9;
  reg  _T_120; // @[FIFO.scala 297:97:@1354.4]
  reg [31:0] _RAND_10;
  reg [2:0] _T_123; // @[FIFO.scala 299:53:@1355.4]
  reg [31:0] _RAND_11;
  wire [3:0] _T_125; // @[FIFO.scala 300:74:@1356.4]
  wire [3:0] _T_126; // @[FIFO.scala 300:74:@1357.4]
  wire [2:0] _T_127; // @[FIFO.scala 300:74:@1358.4]
  wire [2:0] _T_128; // @[FIFO.scala 300:43:@1359.4]
  wire [3:0] _T_130; // @[FIFO.scala 301:68:@1360.4]
  wire [2:0] _T_131; // @[FIFO.scala 301:68:@1361.4]
  wire [2:0] _T_132; // @[FIFO.scala 301:46:@1362.4]
  wire [2:0] _T_133; // @[FIFO.scala 302:32:@1363.4]
  wire  _T_134; // @[FIFO.scala 303:25:@1364.4]
  wire [2:0] _GEN_5; // @[FIFO.scala 303:39:@1365.4]
  wire  _T_137; // @[FIFO.scala 333:77:@1370.4]
  wire  _T_139; // @[FIFO.scala 334:83:@1371.4]
  wire  _T_140; // @[FIFO.scala 335:44:@1372.4]
  wire  _T_141; // @[FIFO.scala 336:60:@1373.4]
  wire  _T_143; // @[FIFO.scala 336:81:@1375.4]
  wire  _GEN_6; // @[FIFO.scala 338:43:@1379.4]
  wire  _T_147; // @[FIFO.scala 341:66:@1382.4]
  wire  _T_148; // @[FIFO.scala 341:63:@1383.4]
  wire  _T_149; // @[FIFO.scala 341:43:@1384.4]
  nv_ram_rwsp_1 nv_ram_rwsp ( // @[FIFO.scala 270:29:@1337.4]
    .io_clk(nv_ram_rwsp_io_clk),
    .io_re(nv_ram_rwsp_io_re),
    .io_we(nv_ram_rwsp_io_we),
    .io_ore(nv_ram_rwsp_io_ore),
    .io_ra(nv_ram_rwsp_io_ra),
    .io_wa(nv_ram_rwsp_io_wa),
    .io_di(nv_ram_rwsp_io_di),
    .io_dout(nv_ram_rwsp_io_dout)
  );
  assign _T_135 = io_rd_pvld & io_rd_prdy; // @[FIFO.scala 331:38:@1368.4]
  assign _T_56 = _T_28 == 1'h0; // @[FIFO.scala 183:39:@1290.4]
  assign _T_57 = _T_31 & _T_56; // @[FIFO.scala 183:36:@1291.4]
  assign _T_69 = _T_62 + 3'h1; // @[FIFO.scala 191:69:@1299.4]
  assign _T_70 = _T_62 + 3'h1; // @[FIFO.scala 191:69:@1300.4]
  assign _T_71 = _T_57 ? _T_70 : _T_62; // @[FIFO.scala 191:46:@1301.4]
  assign _T_74 = _T_71 == 3'h4; // @[FIFO.scala 194:80:@1303.4]
  assign _T_76 = _T_135 ? 1'h0 : _T_74; // @[FIFO.scala 195:40:@1304.4]
  assign _T_64 = _T_62 - 3'h1; // @[FIFO.scala 190:76:@1295.4]
  assign _T_65 = $unsigned(_T_64); // @[FIFO.scala 190:76:@1296.4]
  assign _T_66 = _T_65[2:0]; // @[FIFO.scala 190:76:@1297.4]
  assign _T_67 = _T_57 ? _T_62 : _T_66; // @[FIFO.scala 190:43:@1298.4]
  assign _T_72 = _T_135 ? _T_67 : _T_71; // @[FIFO.scala 192:32:@1302.4]
  assign _T_39 = _T_31 & _T_76; // @[FIFO.scala 166:60:@1271.4]
  assign _T_41 = _T_57 == 1'h0; // @[FIFO.scala 166:80:@1272.4]
  assign _T_42 = _T_39 & _T_41; // @[FIFO.scala 166:77:@1273.4]
  assign _T_43 = io_wr_pvld ? _T_76 : _T_42; // @[FIFO.scala 167:38:@1274.4]
  assign _T_44 = _T_31 & _T_28; // @[FIFO.scala 168:45:@1275.4]
  assign _T_46 = _T_44 == 1'h0; // @[FIFO.scala 171:18:@1277.4]
  assign _T_48 = _T_36 == 1'h0; // @[FIFO.scala 172:45:@1279.6]
  assign _T_49 = io_wr_pvld & _T_48; // @[FIFO.scala 172:42:@1280.6]
  assign _GEN_0 = _T_46 ? _T_49 : _T_31; // @[FIFO.scala 171:34:@1278.4]
  assign _T_52 = _T_48 & io_wr_pvld; // @[FIFO.scala 176:34:@1284.4]
  assign _T_84 = _T_57 ^ _T_135; // @[FIFO.scala 202:27:@1312.4]
  assign _GEN_2 = _T_84 ? _T_72 : _T_62; // @[FIFO.scala 202:40:@1313.4]
  assign _T_86 = _T_72 == 3'h0; // @[FIFO.scala 207:54:@1316.4]
  assign _T_88 = io_wr_pvld == 1'h0; // @[FIFO.scala 207:65:@1317.4]
  assign _T_89 = _T_86 & _T_88; // @[FIFO.scala 207:62:@1318.4]
  assign _T_97 = _T_95 + 2'h1; // @[FIFO.scala 217:42:@1323.4]
  assign _T_98 = _T_95 + 2'h1; // @[FIFO.scala 217:42:@1324.4]
  assign _GEN_3 = _T_57 ? _T_98 : _T_95; // @[FIFO.scala 218:29:@1325.4]
  assign _T_105 = _T_103 + 2'h1; // @[FIFO.scala 225:42:@1330.4]
  assign _T_106 = _T_103 + 2'h1; // @[FIFO.scala 225:42:@1331.4]
  assign _GEN_4 = _T_135 ? _T_106 : _T_103; // @[FIFO.scala 227:29:@1332.4]
  assign _T_125 = _T_123 - 3'h1; // @[FIFO.scala 300:74:@1356.4]
  assign _T_126 = $unsigned(_T_125); // @[FIFO.scala 300:74:@1357.4]
  assign _T_127 = _T_126[2:0]; // @[FIFO.scala 300:74:@1358.4]
  assign _T_128 = _T_114 ? _T_123 : _T_127; // @[FIFO.scala 300:43:@1359.4]
  assign _T_130 = _T_123 + 3'h1; // @[FIFO.scala 301:68:@1360.4]
  assign _T_131 = _T_123 + 3'h1; // @[FIFO.scala 301:68:@1361.4]
  assign _T_132 = _T_114 ? _T_131 : _T_123; // @[FIFO.scala 301:46:@1362.4]
  assign _T_133 = _T_135 ? _T_128 : _T_132; // @[FIFO.scala 302:32:@1363.4]
  assign _T_134 = _T_114 | _T_135; // @[FIFO.scala 303:25:@1364.4]
  assign _GEN_5 = _T_134 ? _T_133 : _T_123; // @[FIFO.scala 303:39:@1365.4]
  assign _T_137 = _T_128 != 3'h0; // @[FIFO.scala 333:77:@1370.4]
  assign _T_139 = _T_132 != 3'h0; // @[FIFO.scala 334:83:@1371.4]
  assign _T_140 = _T_135 ? _T_137 : _T_139; // @[FIFO.scala 335:44:@1372.4]
  assign _T_141 = ~ _T_117; // @[FIFO.scala 336:60:@1373.4]
  assign _T_143 = _T_141 | _T_135; // @[FIFO.scala 336:81:@1375.4]
  assign _GEN_6 = _T_134 ? _T_140 : _T_117; // @[FIFO.scala 338:43:@1379.4]
  assign _T_147 = io_rd_prdy == 1'h0; // @[FIFO.scala 341:66:@1382.4]
  assign _T_148 = _T_120 & _T_147; // @[FIFO.scala 341:63:@1383.4]
  assign _T_149 = _T_117 | _T_148; // @[FIFO.scala 341:43:@1384.4]
  assign io_wr_prdy = _T_36 == 1'h0; // @[FIFO.scala 182:20:@1289.4]
  assign io_wr_empty = _T_92; // @[FIFO.scala 207:29:@1321.4]
  assign io_rd_pvld = _T_120; // @[FIFO.scala 344:24:@1386.4]
  assign io_rd_pd = nv_ram_rwsp_io_dout; // @[FIFO.scala 345:22:@1387.4]
  assign nv_ram_rwsp_io_clk = io_clk; // @[FIFO.scala 271:24:@1340.4]
  assign nv_ram_rwsp_io_re = _T_140 & _T_143; // @[FIFO.scala 279:23:@1347.4]
  assign nv_ram_rwsp_io_we = _T_31 & _T_56; // @[FIFO.scala 276:23:@1343.4]
  assign nv_ram_rwsp_io_ore = io_rd_pvld & io_rd_prdy; // @[FIFO.scala 280:24:@1348.4]
  assign nv_ram_rwsp_io_ra = _T_135 ? _T_106 : _T_103; // @[FIFO.scala 278:23:@1346.4]
  assign nv_ram_rwsp_io_wa = _T_95; // @[FIFO.scala 274:27:@1342.4]
  assign nv_ram_rwsp_io_di = _T_33; // @[FIFO.scala 277:23:@1344.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_28 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_31 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_33 = _RAND_2[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_36 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_62 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_92 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_95 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_103 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_114 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_117 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_120 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_123 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_135) begin
        _T_28 <= 1'h0;
      end else begin
        _T_28 <= _T_74;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_46) begin
        _T_31 <= _T_49;
      end
    end
    if (_T_52) begin
      _T_33 <= io_wr_pd;
    end
    if (reset) begin
      _T_36 <= 1'h0;
    end else begin
      if (io_wr_pvld) begin
        if (_T_135) begin
          _T_36 <= 1'h0;
        end else begin
          _T_36 <= _T_74;
        end
      end else begin
        _T_36 <= _T_42;
      end
    end
    if (reset) begin
      _T_62 <= 3'h0;
    end else begin
      if (_T_84) begin
        if (_T_135) begin
          if (!(_T_57)) begin
            _T_62 <= _T_66;
          end
        end else begin
          if (_T_57) begin
            _T_62 <= _T_70;
          end
        end
      end
    end
    if (reset) begin
      _T_92 <= 1'h1;
    end else begin
      _T_92 <= _T_89;
    end
    if (reset) begin
      _T_95 <= 2'h0;
    end else begin
      if (_T_57) begin
        _T_95 <= _T_98;
      end
    end
    if (reset) begin
      _T_103 <= 2'h0;
    end else begin
      if (_T_135) begin
        _T_103 <= _T_106;
      end
    end
    if (reset) begin
      _T_114 <= 1'h0;
    end else begin
      _T_114 <= _T_57;
    end
    if (reset) begin
      _T_117 <= 1'h0;
    end else begin
      if (_T_134) begin
        if (_T_135) begin
          _T_117 <= _T_137;
        end else begin
          _T_117 <= _T_139;
        end
      end
    end
    if (reset) begin
      _T_120 <= 1'h0;
    end else begin
      _T_120 <= _T_149;
    end
    if (reset) begin
      _T_123 <= 3'h0;
    end else begin
      if (_T_134) begin
        if (_T_135) begin
          if (!(_T_114)) begin
            _T_123 <= _T_127;
          end
        end else begin
          if (_T_114) begin
            _T_123 <= _T_131;
          end
        end
      end
    end
  end
endmodule
module NV_NVDLA_CSC_sg( // @[:@1403.2]
  input         reset, // @[:@1405.4]
  input         io_nvdla_core_clk, // @[:@1406.4]
  input         io_nvdla_core_ng_clk, // @[:@1406.4]
  input         io_cdma2sc_dat_updt_valid, // @[:@1406.4]
  input  [13:0] io_cdma2sc_dat_updt_bits_slices, // @[:@1406.4]
  output        io_sc2cdma_dat_pending_req, // @[:@1406.4]
  input         io_cdma2sc_dat_pending_ack, // @[:@1406.4]
  input         io_cdma2sc_wt_updt_valid, // @[:@1406.4]
  input  [13:0] io_cdma2sc_wt_updt_bits_kernels, // @[:@1406.4]
  output        io_sc2cdma_wt_pending_req, // @[:@1406.4]
  input         io_cdma2sc_wt_pending_ack, // @[:@1406.4]
  output [1:0]  io_sc_state, // @[:@1406.4]
  output        io_sg2dl_pd_valid, // @[:@1406.4]
  output        io_sg2dl_reuse_rls, // @[:@1406.4]
  output        io_sg2wl_pd_valid, // @[:@1406.4]
  output [17:0] io_sg2wl_pd_bits, // @[:@1406.4]
  output        io_sg2wl_reuse_rls, // @[:@1406.4]
  input         io_accu2sc_credit_size_valid, // @[:@1406.4]
  input  [2:0]  io_accu2sc_credit_size_bits, // @[:@1406.4]
  input         io_reg2dp_op_en, // @[:@1406.4]
  input         io_reg2dp_conv_mode, // @[:@1406.4]
  input         io_reg2dp_data_reuse, // @[:@1406.4]
  input         io_reg2dp_skip_data_rls, // @[:@1406.4]
  input         io_reg2dp_weight_reuse, // @[:@1406.4]
  input         io_reg2dp_skip_weight_rls, // @[:@1406.4]
  input         io_reg2dp_datain_format, // @[:@1406.4]
  input  [12:0] io_reg2dp_datain_height_ext, // @[:@1406.4]
  input  [1:0]  io_reg2dp_y_extension, // @[:@1406.4]
  input  [4:0]  io_reg2dp_weight_width_ext, // @[:@1406.4]
  input  [4:0]  io_reg2dp_weight_height_ext, // @[:@1406.4]
  input  [12:0] io_reg2dp_weight_channel_ext, // @[:@1406.4]
  input  [12:0] io_reg2dp_weight_kernel, // @[:@1406.4]
  input  [12:0] io_reg2dp_dataout_width, // @[:@1406.4]
  input  [12:0] io_reg2dp_dataout_height, // @[:@1406.4]
  input  [4:0]  io_reg2dp_data_bank, // @[:@1406.4]
  input  [4:0]  io_reg2dp_weight_bank, // @[:@1406.4]
  input  [20:0] io_reg2dp_atomics, // @[:@1406.4]
  input  [11:0] io_reg2dp_rls_slices, // @[:@1406.4]
  output        io_dp2reg_done // @[:@1406.4]
);
  wire  NV_NVDLA_fifo_clock; // @[NV_NVDLA_CSC_sg.scala 433:28:@1885.4]
  wire  NV_NVDLA_fifo_reset; // @[NV_NVDLA_CSC_sg.scala 433:28:@1885.4]
  wire  NV_NVDLA_fifo_io_clk; // @[NV_NVDLA_CSC_sg.scala 433:28:@1885.4]
  wire  NV_NVDLA_fifo_io_wr_pvld; // @[NV_NVDLA_CSC_sg.scala 433:28:@1885.4]
  wire  NV_NVDLA_fifo_io_wr_prdy; // @[NV_NVDLA_CSC_sg.scala 433:28:@1885.4]
  wire [32:0] NV_NVDLA_fifo_io_wr_pd; // @[NV_NVDLA_CSC_sg.scala 433:28:@1885.4]
  wire  NV_NVDLA_fifo_io_wr_empty; // @[NV_NVDLA_CSC_sg.scala 433:28:@1885.4]
  wire  NV_NVDLA_fifo_io_rd_pvld; // @[NV_NVDLA_CSC_sg.scala 433:28:@1885.4]
  wire  NV_NVDLA_fifo_io_rd_prdy; // @[NV_NVDLA_CSC_sg.scala 433:28:@1885.4]
  wire [32:0] NV_NVDLA_fifo_io_rd_pd; // @[NV_NVDLA_CSC_sg.scala 433:28:@1885.4]
  wire  NV_NVDLA_fifo_1_clock; // @[NV_NVDLA_CSC_sg.scala 446:27:@1896.4]
  wire  NV_NVDLA_fifo_1_reset; // @[NV_NVDLA_CSC_sg.scala 446:27:@1896.4]
  wire  NV_NVDLA_fifo_1_io_clk; // @[NV_NVDLA_CSC_sg.scala 446:27:@1896.4]
  wire  NV_NVDLA_fifo_1_io_wr_pvld; // @[NV_NVDLA_CSC_sg.scala 446:27:@1896.4]
  wire  NV_NVDLA_fifo_1_io_wr_prdy; // @[NV_NVDLA_CSC_sg.scala 446:27:@1896.4]
  wire [19:0] NV_NVDLA_fifo_1_io_wr_pd; // @[NV_NVDLA_CSC_sg.scala 446:27:@1896.4]
  wire  NV_NVDLA_fifo_1_io_wr_empty; // @[NV_NVDLA_CSC_sg.scala 446:27:@1896.4]
  wire  NV_NVDLA_fifo_1_io_rd_pvld; // @[NV_NVDLA_CSC_sg.scala 446:27:@1896.4]
  wire  NV_NVDLA_fifo_1_io_rd_prdy; // @[NV_NVDLA_CSC_sg.scala 446:27:@1896.4]
  wire [19:0] NV_NVDLA_fifo_1_io_rd_pd; // @[NV_NVDLA_CSC_sg.scala 446:27:@1896.4]
  reg  _T_131; // @[NV_NVDLA_CSC_sg.scala 88:29:@1410.4]
  reg [31:0] _RAND_0;
  reg  _T_136; // @[NV_NVDLA_CSC_sg.scala 90:26:@1412.4]
  reg [31:0] _RAND_1;
  reg [1:0] _T_142; // @[NV_NVDLA_CSC_sg.scala 93:28:@1413.4]
  reg [31:0] _RAND_2;
  wire  _T_145; // @[Conditional.scala 37:30:@1416.4]
  reg [4:0] _T_165; // @[NV_NVDLA_CSC_sg.scala 121:33:@1457.4]
  reg [31:0] _RAND_3;
  wire  _T_209; // @[NV_NVDLA_CSC_sg.scala 138:43:@1478.4]
  reg [4:0] _T_168; // @[NV_NVDLA_CSC_sg.scala 122:35:@1458.4]
  reg [31:0] _RAND_4;
  wire  _T_210; // @[NV_NVDLA_CSC_sg.scala 139:44:@1479.4]
  wire  _T_211; // @[NV_NVDLA_CSC_sg.scala 140:38:@1480.4]
  wire  _T_146; // @[NV_NVDLA_CSC_sg.scala 98:31:@1418.6]
  wire [1:0] _GEN_0; // @[NV_NVDLA_CSC_sg.scala 99:37:@1423.8]
  wire [1:0] _GEN_1; // @[NV_NVDLA_CSC_sg.scala 98:47:@1419.6]
  wire  _T_147; // @[Conditional.scala 37:30:@1428.6]
  wire  _T_241; // @[NV_NVDLA_CSC_sg.scala 160:30:@1512.4]
  reg  _T_171; // @[NV_NVDLA_CSC_sg.scala 123:34:@1459.4]
  reg [31:0] _RAND_5;
  reg  _T_174; // @[NV_NVDLA_CSC_sg.scala 124:34:@1460.4]
  reg [31:0] _RAND_6;
  wire  _T_212; // @[NV_NVDLA_CSC_sg.scala 141:51:@1482.4]
  wire  _T_213; // @[NV_NVDLA_CSC_sg.scala 141:34:@1483.4]
  wire  _T_214; // @[NV_NVDLA_CSC_sg.scala 141:32:@1484.4]
  reg  _T_180; // @[NV_NVDLA_CSC_sg.scala 126:33:@1462.4]
  reg [31:0] _RAND_7;
  reg  _T_183; // @[NV_NVDLA_CSC_sg.scala 127:33:@1463.4]
  reg [31:0] _RAND_8;
  wire  _T_215; // @[NV_NVDLA_CSC_sg.scala 141:87:@1485.4]
  wire  _T_216; // @[NV_NVDLA_CSC_sg.scala 141:71:@1486.4]
  wire  _T_217; // @[NV_NVDLA_CSC_sg.scala 141:69:@1487.4]
  wire [1:0] _GEN_2; // @[NV_NVDLA_CSC_sg.scala 102:29:@1430.8]
  wire  _T_148; // @[Conditional.scala 37:30:@1435.8]
  wire  _T_154; // @[NV_NVDLA_CSC_sg.scala 116:27:@1452.4 NV_NVDLA_CSC_sg.scala 441:17:@1893.4]
  wire  _T_204; // @[NV_NVDLA_CSC_sg.scala 137:22:@1472.4]
  wire  _T_160; // @[NV_NVDLA_CSC_sg.scala 119:26:@1455.4 NV_NVDLA_CSC_sg.scala 454:16:@1904.4]
  wire  _T_205; // @[NV_NVDLA_CSC_sg.scala 137:37:@1473.4]
  wire  _T_206; // @[NV_NVDLA_CSC_sg.scala 137:35:@1474.4]
  wire  _T_156; // @[NV_NVDLA_CSC_sg.scala 117:30:@1453.4 NV_NVDLA_CSC_sg.scala 444:20:@1895.4]
  wire  _T_207; // @[NV_NVDLA_CSC_sg.scala 137:49:@1475.4]
  wire  _T_162; // @[NV_NVDLA_CSC_sg.scala 120:29:@1456.4 NV_NVDLA_CSC_sg.scala 457:19:@1906.4]
  wire  _T_208; // @[NV_NVDLA_CSC_sg.scala 137:66:@1476.4]
  wire  _T_149; // @[NV_NVDLA_CSC_sg.scala 105:26:@1437.10]
  wire  _T_150; // @[NV_NVDLA_CSC_sg.scala 105:44:@1438.10]
  wire  _T_151; // @[NV_NVDLA_CSC_sg.scala 105:42:@1439.10]
  wire [1:0] _GEN_3; // @[NV_NVDLA_CSC_sg.scala 105:54:@1440.10]
  wire [1:0] _GEN_6; // @[Conditional.scala 39:67:@1436.8]
  wire [1:0] _GEN_7; // @[Conditional.scala 39:67:@1429.6]
  wire [1:0] _GEN_8; // @[Conditional.scala 40:58:@1417.4]
  reg  _T_177; // @[NV_NVDLA_CSC_sg.scala 125:34:@1461.4]
  reg [31:0] _RAND_9;
  reg  _T_186; // @[NV_NVDLA_CSC_sg.scala 128:33:@1464.4]
  reg [31:0] _RAND_10;
  reg [6:0] _T_191; // @[NV_NVDLA_CSC_sg.scala 130:34:@1466.4]
  reg [31:0] _RAND_11;
  reg [7:0] _T_198; // @[NV_NVDLA_CSC_sg.scala 133:31:@1469.4]
  reg [31:0] _RAND_12;
  reg [7:0] _T_201; // @[NV_NVDLA_CSC_sg.scala 134:28:@1470.4]
  reg [31:0] _RAND_13;
  wire  _T_243; // @[NV_NVDLA_CSC_sg.scala 162:27:@1515.4]
  wire  _T_218; // @[NV_NVDLA_CSC_sg.scala 144:26:@1490.6]
  wire  _T_244; // @[NV_NVDLA_CSC_sg.scala 163:31:@1517.4]
  wire  _T_219; // @[NV_NVDLA_CSC_sg.scala 144:35:@1491.6]
  wire [8:0] _T_221; // @[NV_NVDLA_CSC_sg.scala 144:74:@1492.6]
  wire [8:0] _T_222; // @[NV_NVDLA_CSC_sg.scala 144:74:@1493.6]
  wire [7:0] _T_223; // @[NV_NVDLA_CSC_sg.scala 144:74:@1494.6]
  wire [7:0] _T_224; // @[NV_NVDLA_CSC_sg.scala 144:25:@1495.6]
  wire [7:0] _GEN_9; // @[NV_NVDLA_CSC_sg.scala 143:22:@1489.4]
  reg [5:0] _T_799; // @[NV_NVDLA_CSC_sg.scala 501:26:@1946.4]
  reg [31:0] _RAND_14;
  wire  _T_861; // @[NV_NVDLA_CSC_sg.scala 521:45:@1986.4]
  wire  _T_862; // @[NV_NVDLA_CSC_sg.scala 521:34:@1987.4]
  wire [30:0] _T_748; // @[NV_NVDLA_CSC_sg.scala 463:34:@1908.4]
  wire  _T_757; // @[NV_NVDLA_CSC_sg.scala 474:40:@1917.4]
  wire  _T_883; // @[NV_NVDLA_CSC_sg.scala 561:21:@2023.4]
  reg [8:0] _T_870; // @[NV_NVDLA_CSC_sg.scala 548:61:@2012.4]
  reg [31:0] _RAND_15;
  wire [8:0] _T_877; // @[Cat.scala 30:58:@2019.4]
  wire  _T_884; // @[NV_NVDLA_CSC_sg.scala 561:55:@2024.4]
  wire  _T_885; // @[NV_NVDLA_CSC_sg.scala 561:41:@2025.4]
  wire  _T_863; // @[NV_NVDLA_CSC_sg.scala 521:54:@1988.4]
  wire [1:0] _T_747; // @[NV_NVDLA_CSC_sg.scala 462:35:@1907.4]
  wire [1:0] _T_749; // @[NV_NVDLA_CSC_sg.scala 464:33:@1909.4]
  wire  _T_864; // @[NV_NVDLA_CSC_sg.scala 521:85:@1989.4]
  wire  _T_866; // @[NV_NVDLA_CSC_sg.scala 521:101:@1991.4]
  wire  _T_867; // @[NV_NVDLA_CSC_sg.scala 521:69:@1992.4]
  wire  _T_225; // @[NV_NVDLA_CSC_sg.scala 148:22:@1500.4]
  wire  _T_759; // @[NV_NVDLA_CSC_sg.scala 476:35:@1919.4]
  wire  _T_226; // @[NV_NVDLA_CSC_sg.scala 148:38:@1501.4]
  wire [7:0] _T_228; // @[NV_NVDLA_CSC_sg.scala 149:41:@1503.6]
  wire [7:0] _GEN_10; // @[NV_NVDLA_CSC_sg.scala 148:57:@1502.4]
  reg [2:0] _T_237; // @[NV_NVDLA_CSC_sg.scala 156:28:@1508.4]
  reg [31:0] _RAND_16;
  wire  _T_238; // @[NV_NVDLA_CSC_sg.scala 158:49:@1509.4]
  wire  _T_239; // @[NV_NVDLA_CSC_sg.scala 158:36:@1510.4]
  wire  _T_242; // @[NV_NVDLA_CSC_sg.scala 161:33:@1514.4]
  wire  _T_245; // @[NV_NVDLA_CSC_sg.scala 164:37:@1519.4]
  wire [1:0] _T_250; // @[NV_NVDLA_CSC_sg.scala 165:90:@1520.4]
  wire [1:0] _T_251; // @[NV_NVDLA_CSC_sg.scala 165:55:@1521.4]
  wire  _T_312; // @[NV_NVDLA_CSC_sg.scala 199:40:@1568.4]
  wire  _T_313; // @[NV_NVDLA_CSC_sg.scala 200:26:@1569.4]
  wire  _T_314; // @[NV_NVDLA_CSC_sg.scala 201:27:@1570.4]
  wire  _T_315; // @[NV_NVDLA_CSC_sg.scala 201:25:@1571.4]
  wire [2:0] _T_318; // @[Cat.scala 30:58:@1573.4]
  wire  _T_253; // @[NV_NVDLA_CSC_sg.scala 166:37:@1524.4]
  wire  _T_255; // @[NV_NVDLA_CSC_sg.scala 168:53:@1525.4]
  wire  _T_256; // @[NV_NVDLA_CSC_sg.scala 168:39:@1526.4]
  reg  _T_259; // @[NV_NVDLA_CSC_sg.scala 168:30:@1527.4]
  reg [31:0] _RAND_17;
  wire  _T_260; // @[NV_NVDLA_CSC_sg.scala 169:43:@1530.4]
  wire  _T_262; // @[NV_NVDLA_CSC_sg.scala 169:85:@1531.4]
  wire  _T_264; // @[NV_NVDLA_CSC_sg.scala 169:83:@1532.4]
  wire  _T_265; // @[NV_NVDLA_CSC_sg.scala 169:27:@1533.4]
  wire  _T_269; // @[NV_NVDLA_CSC_sg.scala 170:64:@1536.4]
  wire  _T_270; // @[NV_NVDLA_CSC_sg.scala 170:26:@1537.4]
  wire  _T_271; // @[NV_NVDLA_CSC_sg.scala 171:39:@1539.4]
  wire  _T_275; // @[NV_NVDLA_CSC_sg.scala 171:79:@1541.4]
  wire  _T_276; // @[NV_NVDLA_CSC_sg.scala 171:27:@1542.4]
  wire  _T_277; // @[NV_NVDLA_CSC_sg.scala 172:38:@1544.4]
  wire  _T_281; // @[NV_NVDLA_CSC_sg.scala 172:77:@1546.4]
  wire  _T_282; // @[NV_NVDLA_CSC_sg.scala 172:26:@1547.4]
  reg [13:0] _T_289; // @[NV_NVDLA_CSC_sg.scala 181:30:@1552.4]
  reg [31:0] _RAND_18;
  reg [13:0] _T_296; // @[NV_NVDLA_CSC_sg.scala 182:29:@1554.4]
  reg [31:0] _RAND_19;
  reg [13:0] _T_303; // @[NV_NVDLA_CSC_sg.scala 183:31:@1556.4]
  reg [31:0] _RAND_20;
  reg  _T_306; // @[NV_NVDLA_CSC_sg.scala 184:39:@1557.4]
  reg [31:0] _RAND_21;
  wire [13:0] _T_308; // @[NV_NVDLA_CSC_sg.scala 190:49:@1562.6]
  wire [4:0] _GEN_11; // @[NV_NVDLA_CSC_sg.scala 186:25:@1558.4]
  wire [4:0] _GEN_12; // @[NV_NVDLA_CSC_sg.scala 186:25:@1558.4]
  wire [13:0] _GEN_13; // @[NV_NVDLA_CSC_sg.scala 186:25:@1558.4]
  wire [13:0] _GEN_14; // @[NV_NVDLA_CSC_sg.scala 186:25:@1558.4]
  wire  _GEN_15; // @[NV_NVDLA_CSC_sg.scala 186:25:@1558.4]
  wire [2:0] _GEN_16; // @[NV_NVDLA_CSC_sg.scala 186:25:@1558.4]
  reg [13:0] _T_326; // @[NV_NVDLA_CSC_sg.scala 207:33:@1576.4]
  reg [31:0] _RAND_22;
  reg [21:0] _T_333; // @[NV_NVDLA_CSC_sg.scala 208:34:@1578.4]
  reg [31:0] _RAND_23;
  reg [4:0] _T_347; // @[NV_NVDLA_CSC_sg.scala 210:35:@1582.4]
  reg [31:0] _RAND_24;
  reg [4:0] _T_354; // @[NV_NVDLA_CSC_sg.scala 211:36:@1584.4]
  reg [31:0] _RAND_25;
  reg [13:0] _T_361; // @[NV_NVDLA_CSC_sg.scala 212:33:@1586.4]
  reg [31:0] _RAND_26;
  reg [9:0] _T_368; // @[NV_NVDLA_CSC_sg.scala 213:32:@1588.4]
  reg [31:0] _RAND_27;
  reg [2:0] _T_371; // @[NV_NVDLA_CSC_sg.scala 214:31:@1589.4]
  reg [31:0] _RAND_28;
  reg [2:0] _T_374; // @[NV_NVDLA_CSC_sg.scala 215:32:@1590.4]
  reg [31:0] _RAND_29;
  reg [13:0] _T_381; // @[NV_NVDLA_CSC_sg.scala 216:29:@1592.4]
  reg [31:0] _RAND_30;
  reg  _T_384; // @[NV_NVDLA_CSC_sg.scala 217:28:@1593.4]
  reg [31:0] _RAND_31;
  reg [5:0] _T_387; // @[NV_NVDLA_CSC_sg.scala 218:30:@1594.4]
  reg [31:0] _RAND_32;
  reg [6:0] _T_390; // @[NV_NVDLA_CSC_sg.scala 219:30:@1595.4]
  reg [31:0] _RAND_33;
  wire [8:0] _T_392; // @[NV_NVDLA_CSC_sg.scala 221:44:@1596.4]
  wire [2:0] _T_393; // @[NV_NVDLA_CSC_sg.scala 221:69:@1597.4]
  wire [13:0] _T_395; // @[NV_NVDLA_CSC_sg.scala 224:55:@1599.6]
  wire [13:0] _T_397; // @[NV_NVDLA_CSC_sg.scala 225:64:@1601.6]
  wire [21:0] _T_399; // @[NV_NVDLA_CSC_sg.scala 225:90:@1602.6]
  wire [21:0] _T_400; // @[NV_NVDLA_CSC_sg.scala 225:31:@1603.6]
  wire [4:0] _T_403; // @[NV_NVDLA_CSC_sg.scala 227:32:@1606.6]
  wire [13:0] _T_405; // @[NV_NVDLA_CSC_sg.scala 229:56:@1609.6]
  wire [7:0] _T_406; // @[NV_NVDLA_CSC_sg.scala 230:49:@1611.6]
  wire [8:0] _T_408; // @[NV_NVDLA_CSC_sg.scala 230:71:@1612.6]
  wire  _T_409; // @[NV_NVDLA_CSC_sg.scala 232:44:@1615.6]
  wire  _T_411; // @[NV_NVDLA_CSC_sg.scala 233:44:@1616.6]
  wire  _T_413; // @[NV_NVDLA_CSC_sg.scala 233:98:@1617.6]
  wire [1:0] _T_414; // @[Cat.scala 30:58:@1618.6]
  wire [1:0] _T_415; // @[NV_NVDLA_CSC_sg.scala 234:55:@1619.6]
  wire [1:0] _T_416; // @[NV_NVDLA_CSC_sg.scala 233:29:@1620.6]
  wire [1:0] _T_417; // @[NV_NVDLA_CSC_sg.scala 232:29:@1621.6]
  wire [12:0] _T_419; // @[NV_NVDLA_CSC_sg.scala 235:44:@1623.6]
  wire [11:0] _T_420; // @[NV_NVDLA_CSC_sg.scala 235:44:@1624.6]
  wire [12:0] _GEN_62; // @[NV_NVDLA_CSC_sg.scala 236:116:@1627.6]
  wire [13:0] _T_423; // @[NV_NVDLA_CSC_sg.scala 236:116:@1627.6]
  wire [13:0] _T_424; // @[NV_NVDLA_CSC_sg.scala 236:116:@1628.6]
  wire [13:0] _T_425; // @[NV_NVDLA_CSC_sg.scala 236:26:@1629.6]
  wire [6:0] _T_428; // @[NV_NVDLA_CSC_sg.scala 240:27:@1632.6]
  wire [13:0] _GEN_17; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  wire [21:0] _GEN_18; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  wire [4:0] _GEN_20; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  wire [4:0] _GEN_21; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  wire [13:0] _GEN_22; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  wire [9:0] _GEN_23; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  wire [2:0] _GEN_24; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  wire [2:0] _GEN_25; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  wire [13:0] _GEN_26; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  wire [13:0] _GEN_27; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  wire  _GEN_28; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  wire [6:0] _GEN_29; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  wire [6:0] _GEN_30; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  reg [13:0] _T_593; // @[NV_NVDLA_CSC_sg.scala 333:29:@1747.4]
  reg [31:0] _RAND_34;
  wire  _T_600; // @[NV_NVDLA_CSC_sg.scala 337:38:@1750.4]
  reg [13:0] _T_596; // @[NV_NVDLA_CSC_sg.scala 334:35:@1748.4]
  reg [31:0] _RAND_35;
  reg [9:0] _T_449; // @[NV_NVDLA_CSC_sg.scala 257:31:@1647.4]
  reg [31:0] _RAND_36;
  wire [10:0] _T_451; // @[NV_NVDLA_CSC_sg.scala 258:41:@1648.4]
  wire [9:0] _T_452; // @[NV_NVDLA_CSC_sg.scala 258:41:@1649.4]
  wire  _T_453; // @[NV_NVDLA_CSC_sg.scala 259:40:@1650.4]
  wire  _T_454; // @[NV_NVDLA_CSC_sg.scala 260:26:@1652.4]
  wire [4:0] _T_456; // @[NV_NVDLA_CSC_sg.scala 260:87:@1653.4]
  wire [5:0] _T_458; // @[NV_NVDLA_CSC_sg.scala 260:110:@1654.4]
  wire [5:0] _T_459; // @[NV_NVDLA_CSC_sg.scala 260:25:@1655.4]
  wire [13:0] _GEN_63; // @[NV_NVDLA_CSC_sg.scala 338:49:@1751.4]
  wire [14:0] _T_601; // @[NV_NVDLA_CSC_sg.scala 338:49:@1751.4]
  wire [13:0] _T_602; // @[NV_NVDLA_CSC_sg.scala 338:49:@1752.4]
  reg [14:0] _T_599; // @[NV_NVDLA_CSC_sg.scala 335:30:@1749.4]
  reg [31:0] _RAND_37;
  wire [14:0] _GEN_64; // @[NV_NVDLA_CSC_sg.scala 339:46:@1753.4]
  wire  _T_603; // @[NV_NVDLA_CSC_sg.scala 339:46:@1753.4]
  wire  _T_615; // @[NV_NVDLA_CSC_sg.scala 350:37:@1765.4]
  wire  _T_616; // @[NV_NVDLA_CSC_sg.scala 351:30:@1766.4]
  wire  _T_617; // @[NV_NVDLA_CSC_sg.scala 351:45:@1767.4]
  wire  _T_618; // @[NV_NVDLA_CSC_sg.scala 351:43:@1768.4]
  wire  _T_611; // @[NV_NVDLA_CSC_sg.scala 346:30:@1762.4 NV_NVDLA_CSC_sg.scala 439:20:@1891.4]
  wire  _T_613; // @[NV_NVDLA_CSC_sg.scala 347:29:@1763.4 NV_NVDLA_CSC_sg.scala 452:19:@1902.4]
  wire  _T_614; // @[NV_NVDLA_CSC_sg.scala 349:42:@1764.4]
  wire  _T_620; // @[NV_NVDLA_CSC_sg.scala 351:69:@1770.4]
  wire  _T_621; // @[NV_NVDLA_CSC_sg.scala 351:57:@1771.4]
  reg [4:0] _T_554; // @[NV_NVDLA_CSC_sg.scala 308:34:@1721.4]
  reg [31:0] _RAND_38;
  wire  _T_570; // @[NV_NVDLA_CSC_sg.scala 315:38:@1729.4]
  reg [4:0] _T_561; // @[NV_NVDLA_CSC_sg.scala 309:34:@1723.4]
  reg [31:0] _RAND_39;
  wire [4:0] _GEN_65; // @[NV_NVDLA_CSC_sg.scala 314:47:@1728.4]
  wire [5:0] _T_569; // @[NV_NVDLA_CSC_sg.scala 314:47:@1728.4]
  wire [5:0] _GEN_66; // @[NV_NVDLA_CSC_sg.scala 316:42:@1730.4]
  wire  _T_571; // @[NV_NVDLA_CSC_sg.scala 316:42:@1730.4]
  wire  _T_580; // @[NV_NVDLA_CSC_sg.scala 322:35:@1736.4]
  wire  _T_634; // @[NV_NVDLA_CSC_sg.scala 358:28:@1790.4]
  reg [13:0] _T_524; // @[NV_NVDLA_CSC_sg.scala 297:33:@1704.4]
  reg [31:0] _RAND_40;
  wire [14:0] _T_526; // @[NV_NVDLA_CSC_sg.scala 298:45:@1705.4]
  wire [13:0] _T_527; // @[NV_NVDLA_CSC_sg.scala 298:45:@1706.4]
  wire  _T_528; // @[NV_NVDLA_CSC_sg.scala 299:47:@1707.4]
  wire  _T_635; // @[NV_NVDLA_CSC_sg.scala 358:44:@1791.4]
  reg [21:0] _T_489; // @[NV_NVDLA_CSC_sg.scala 278:32:@1676.4]
  reg [31:0] _RAND_41;
  wire [21:0] _GEN_67; // @[NV_NVDLA_CSC_sg.scala 280:47:@1680.4]
  wire [22:0] _T_494; // @[NV_NVDLA_CSC_sg.scala 280:47:@1680.4]
  wire [21:0] _T_495; // @[NV_NVDLA_CSC_sg.scala 280:47:@1681.4]
  wire  _T_497; // @[NV_NVDLA_CSC_sg.scala 282:49:@1683.4]
  wire  _T_636; // @[NV_NVDLA_CSC_sg.scala 358:62:@1792.4]
  wire  _T_472; // @[NV_NVDLA_CSC_sg.scala 270:24:@1664.4]
  reg [12:0] _T_469; // @[NV_NVDLA_CSC_sg.scala 267:35:@1662.4]
  reg [31:0] _RAND_42;
  wire  _T_473; // @[NV_NVDLA_CSC_sg.scala 270:55:@1665.4]
  wire  _T_474; // @[NV_NVDLA_CSC_sg.scala 270:35:@1666.4]
  wire  _T_637; // @[NV_NVDLA_CSC_sg.scala 358:79:@1793.4]
  wire  _T_638; // @[NV_NVDLA_CSC_sg.scala 358:94:@1794.4]
  wire  _T_436; // @[NV_NVDLA_CSC_sg.scala 251:19:@1639.4]
  wire  _T_439; // @[NV_NVDLA_CSC_sg.scala 252:48:@1641.6]
  wire  _T_440; // @[NV_NVDLA_CSC_sg.scala 252:25:@1642.6]
  wire  _GEN_31; // @[NV_NVDLA_CSC_sg.scala 251:33:@1640.4]
  wire  _T_460; // @[NV_NVDLA_CSC_sg.scala 262:19:@1656.4]
  wire [9:0] _T_462; // @[NV_NVDLA_CSC_sg.scala 263:27:@1658.6]
  wire [9:0] _GEN_32; // @[NV_NVDLA_CSC_sg.scala 262:33:@1657.4]
  wire  _T_626; // @[NV_NVDLA_CSC_sg.scala 356:29:@1780.4]
  wire  _T_627; // @[NV_NVDLA_CSC_sg.scala 356:39:@1781.4]
  wire  _T_628; // @[NV_NVDLA_CSC_sg.scala 356:55:@1782.4]
  wire  _T_629; // @[NV_NVDLA_CSC_sg.scala 356:73:@1783.4]
  wire  _T_475; // @[NV_NVDLA_CSC_sg.scala 271:19:@1667.4]
  wire [13:0] _T_479; // @[NV_NVDLA_CSC_sg.scala 274:47:@1669.6]
  wire [12:0] _T_480; // @[NV_NVDLA_CSC_sg.scala 274:47:@1670.6]
  wire [12:0] _T_481; // @[NV_NVDLA_CSC_sg.scala 273:32:@1671.6]
  wire [12:0] _T_482; // @[NV_NVDLA_CSC_sg.scala 272:32:@1672.6]
  wire [12:0] _GEN_33; // @[NV_NVDLA_CSC_sg.scala 271:32:@1668.4]
  wire [7:0] _T_491; // @[Cat.scala 30:58:@1677.4]
  wire [21:0] _GEN_68; // @[NV_NVDLA_CSC_sg.scala 279:46:@1678.4]
  wire [22:0] _T_492; // @[NV_NVDLA_CSC_sg.scala 279:46:@1678.4]
  wire [21:0] _T_493; // @[NV_NVDLA_CSC_sg.scala 279:46:@1679.4]
  wire  _T_496; // @[NV_NVDLA_CSC_sg.scala 281:49:@1682.4]
  wire [22:0] _T_498; // @[NV_NVDLA_CSC_sg.scala 284:43:@1684.4]
  wire [22:0] _T_499; // @[NV_NVDLA_CSC_sg.scala 284:43:@1685.4]
  wire [21:0] _T_500; // @[NV_NVDLA_CSC_sg.scala 284:43:@1686.4]
  wire [6:0] _T_501; // @[NV_NVDLA_CSC_sg.scala 284:60:@1687.4]
  wire [6:0] _T_502; // @[NV_NVDLA_CSC_sg.scala 285:59:@1688.4]
  wire [6:0] _T_503; // @[NV_NVDLA_CSC_sg.scala 285:25:@1689.4]
  wire  _T_506; // @[NV_NVDLA_CSC_sg.scala 288:19:@1691.4]
  wire [21:0] _GEN_70; // @[NV_NVDLA_CSC_sg.scala 292:41:@1695.6]
  wire [22:0] _T_511; // @[NV_NVDLA_CSC_sg.scala 292:41:@1695.6]
  wire [21:0] _T_512; // @[NV_NVDLA_CSC_sg.scala 292:41:@1696.6]
  wire [21:0] _T_513; // @[NV_NVDLA_CSC_sg.scala 291:29:@1697.6]
  wire [21:0] _T_514; // @[NV_NVDLA_CSC_sg.scala 290:29:@1698.6]
  wire [21:0] _T_515; // @[NV_NVDLA_CSC_sg.scala 289:29:@1699.6]
  wire [21:0] _GEN_34; // @[NV_NVDLA_CSC_sg.scala 288:34:@1692.4]
  wire  _T_529; // @[NV_NVDLA_CSC_sg.scala 301:27:@1708.4]
  wire [5:0] _T_531; // @[NV_NVDLA_CSC_sg.scala 301:93:@1709.4]
  wire [6:0] _T_533; // @[NV_NVDLA_CSC_sg.scala 301:117:@1710.4]
  wire [6:0] _T_534; // @[NV_NVDLA_CSC_sg.scala 301:26:@1711.4]
  wire  _T_535; // @[NV_NVDLA_CSC_sg.scala 303:19:@1712.4]
  wire [13:0] _T_546; // @[NV_NVDLA_CSC_sg.scala 304:63:@1716.6]
  wire [13:0] _T_547; // @[NV_NVDLA_CSC_sg.scala 304:30:@1717.6]
  wire [13:0] _GEN_35; // @[NV_NVDLA_CSC_sg.scala 303:35:@1713.4]
  wire [5:0] _T_567; // @[NV_NVDLA_CSC_sg.scala 313:47:@1726.4]
  wire [4:0] _T_568; // @[NV_NVDLA_CSC_sg.scala 313:47:@1727.4]
  wire  _T_572; // @[NV_NVDLA_CSC_sg.scala 318:33:@1731.4]
  wire  _T_574; // @[NV_NVDLA_CSC_sg.scala 319:33:@1732.4]
  wire [1:0] _T_577; // @[NV_NVDLA_CSC_sg.scala 319:20:@1733.4]
  wire [1:0] _T_578; // @[NV_NVDLA_CSC_sg.scala 318:20:@1734.4]
  wire [2:0] _T_579; // @[NV_NVDLA_CSC_sg.scala 317:20:@1735.4]
  wire  _T_581; // @[NV_NVDLA_CSC_sg.scala 324:19:@1737.4]
  wire [4:0] _T_584; // @[NV_NVDLA_CSC_sg.scala 326:32:@1739.6]
  wire [4:0] _T_585; // @[NV_NVDLA_CSC_sg.scala 325:31:@1740.6]
  wire [4:0] _T_588; // @[NV_NVDLA_CSC_sg.scala 330:48:@1742.6]
  wire [4:0] _T_589; // @[NV_NVDLA_CSC_sg.scala 329:32:@1743.6]
  wire [4:0] _T_590; // @[NV_NVDLA_CSC_sg.scala 328:31:@1744.6]
  wire [4:0] _GEN_36; // @[NV_NVDLA_CSC_sg.scala 324:29:@1738.4]
  wire [4:0] _GEN_37; // @[NV_NVDLA_CSC_sg.scala 324:29:@1738.4]
  wire  _T_605; // @[NV_NVDLA_CSC_sg.scala 342:43:@1756.6]
  wire  _T_606; // @[NV_NVDLA_CSC_sg.scala 342:61:@1757.6]
  wire  _T_607; // @[NV_NVDLA_CSC_sg.scala 342:59:@1758.6]
  wire [13:0] _T_609; // @[NV_NVDLA_CSC_sg.scala 342:32:@1759.6]
  wire [13:0] _GEN_38; // @[NV_NVDLA_CSC_sg.scala 341:33:@1755.4]
  wire  _T_639; // @[NV_NVDLA_CSC_sg.scala 360:20:@1796.4]
  wire  _T_642; // @[NV_NVDLA_CSC_sg.scala 360:57:@1798.4]
  wire  _T_645; // @[NV_NVDLA_CSC_sg.scala 360:83:@1799.4]
  wire  _T_646; // @[NV_NVDLA_CSC_sg.scala 360:45:@1800.4]
  wire  _T_647; // @[NV_NVDLA_CSC_sg.scala 360:19:@1801.4]
  reg [1:0] _T_654; // @[NV_NVDLA_CSC_sg.scala 363:26:@1804.4]
  reg [31:0] _RAND_43;
  reg [4:0] _T_657; // @[NV_NVDLA_CSC_sg.scala 364:35:@1805.4]
  reg [31:0] _RAND_44;
  reg [4:0] _T_660; // @[NV_NVDLA_CSC_sg.scala 365:35:@1806.4]
  reg [31:0] _RAND_45;
  reg [6:0] _T_663; // @[NV_NVDLA_CSC_sg.scala 366:39:@1807.4]
  reg [31:0] _RAND_46;
  reg [6:0] _T_666; // @[NV_NVDLA_CSC_sg.scala 367:40:@1808.4]
  reg [31:0] _RAND_47;
  reg [2:0] _T_669; // @[NV_NVDLA_CSC_sg.scala 368:36:@1809.4]
  reg [31:0] _RAND_48;
  reg  _T_672; // @[NV_NVDLA_CSC_sg.scala 369:36:@1810.4]
  reg [31:0] _RAND_49;
  reg  _T_675; // @[NV_NVDLA_CSC_sg.scala 370:38:@1811.4]
  reg [31:0] _RAND_50;
  reg  _T_678; // @[NV_NVDLA_CSC_sg.scala 371:36:@1812.4]
  reg [31:0] _RAND_51;
  reg  _T_681; // @[NV_NVDLA_CSC_sg.scala 372:36:@1813.4]
  reg [31:0] _RAND_52;
  reg  _T_684; // @[NV_NVDLA_CSC_sg.scala 373:38:@1814.4]
  reg [31:0] _RAND_53;
  wire [2:0] _T_687; // @[NV_NVDLA_CSC_sg.scala 375:61:@1815.4]
  wire [1:0] _T_688; // @[NV_NVDLA_CSC_sg.scala 375:61:@1816.4]
  wire [1:0] _T_689; // @[NV_NVDLA_CSC_sg.scala 375:24:@1817.4]
  wire  _T_690; // @[NV_NVDLA_CSC_sg.scala 379:43:@1818.4]
  wire  _T_692; // @[NV_NVDLA_CSC_sg.scala 380:59:@1820.4]
  wire  _T_693; // @[NV_NVDLA_CSC_sg.scala 380:76:@1821.4]
  wire  _T_697; // @[NV_NVDLA_CSC_sg.scala 381:91:@1825.4]
  wire [1:0] _GEN_39; // @[NV_NVDLA_CSC_sg.scala 383:29:@1827.4]
  wire  _T_704; // @[NV_NVDLA_CSC_sg.scala 396:32:@1843.6]
  wire  _T_705; // @[NV_NVDLA_CSC_sg.scala 396:57:@1844.6]
  wire [4:0] _GEN_40; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  wire [4:0] _GEN_41; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  wire [6:0] _GEN_42; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  wire [6:0] _GEN_43; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  wire [2:0] _GEN_44; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  wire  _GEN_45; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  wire  _GEN_46; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  wire  _GEN_47; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  wire  _GEN_48; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  wire  _GEN_49; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  reg [6:0] _T_708; // @[NV_NVDLA_CSC_sg.scala 400:37:@1847.4]
  reg [31:0] _RAND_54;
  reg [6:0] _T_711; // @[NV_NVDLA_CSC_sg.scala 401:37:@1848.4]
  reg [31:0] _RAND_55;
  reg [2:0] _T_714; // @[NV_NVDLA_CSC_sg.scala 402:35:@1849.4]
  reg [31:0] _RAND_56;
  reg  _T_717; // @[NV_NVDLA_CSC_sg.scala 403:36:@1850.4]
  reg [31:0] _RAND_57;
  wire [1:0] _T_718; // @[NV_NVDLA_CSC_sg.scala 406:42:@1851.4]
  wire [30:0] _T_731; // @[Cat.scala 30:58:@1864.4]
  wire  _T_734; // @[NV_NVDLA_CSC_sg.scala 415:57:@1871.6]
  wire [6:0] _GEN_50; // @[NV_NVDLA_CSC_sg.scala 411:18:@1866.4]
  wire [6:0] _GEN_51; // @[NV_NVDLA_CSC_sg.scala 411:18:@1866.4]
  wire [2:0] _GEN_52; // @[NV_NVDLA_CSC_sg.scala 411:18:@1866.4]
  wire  _GEN_53; // @[NV_NVDLA_CSC_sg.scala 411:18:@1866.4]
  wire [1:0] _T_735; // @[NV_NVDLA_CSC_sg.scala 423:41:@1874.4]
  wire [5:0] _T_736; // @[NV_NVDLA_CSC_sg.scala 423:67:@1875.4]
  wire [17:0] _T_741; // @[Cat.scala 30:58:@1880.4]
  wire [17:0] _T_750; // @[NV_NVDLA_CSC_sg.scala 465:32:@1910.4]
  wire [6:0] _T_754; // @[NV_NVDLA_CSC_sg.scala 471:42:@1914.4]
  wire [5:0] _T_762; // @[NV_NVDLA_CSC_sg.scala 481:38:@1923.4]
  wire  _T_774; // @[NV_NVDLA_CSC_sg.scala 492:61:@1932.4]
  wire [7:0] _T_776; // @[NV_NVDLA_CSC_sg.scala 492:106:@1933.4]
  wire [7:0] _T_778; // @[NV_NVDLA_CSC_sg.scala 492:127:@1934.4]
  wire [6:0] _T_779; // @[NV_NVDLA_CSC_sg.scala 492:147:@1935.4]
  wire  _T_781; // @[NV_NVDLA_CSC_sg.scala 493:61:@1936.4]
  wire [7:0] _T_783; // @[NV_NVDLA_CSC_sg.scala 493:106:@1937.4]
  wire [7:0] _T_785; // @[NV_NVDLA_CSC_sg.scala 493:127:@1938.4]
  wire [6:0] _T_786; // @[NV_NVDLA_CSC_sg.scala 493:147:@1939.4]
  wire [6:0] _T_787; // @[NV_NVDLA_CSC_sg.scala 493:38:@1940.4]
  wire [6:0] _T_788; // @[NV_NVDLA_CSC_sg.scala 492:38:@1941.4]
  wire [6:0] _T_789; // @[NV_NVDLA_CSC_sg.scala 491:38:@1942.4]
  wire [6:0] _T_790; // @[NV_NVDLA_CSC_sg.scala 496:34:@1943.4]
  reg  _T_793; // @[NV_NVDLA_CSC_sg.scala 499:34:@1944.4]
  reg [31:0] _RAND_58;
  reg [6:0] _T_796; // @[NV_NVDLA_CSC_sg.scala 500:36:@1945.4]
  reg [31:0] _RAND_59;
  reg  _T_802; // @[NV_NVDLA_CSC_sg.scala 502:33:@1947.4]
  reg [31:0] _RAND_60;
  reg  _T_808; // @[NV_NVDLA_CSC_sg.scala 504:33:@1949.4]
  reg [31:0] _RAND_61;
  reg [17:0] _T_811; // @[NV_NVDLA_CSC_sg.scala 505:31:@1950.4]
  reg [31:0] _RAND_62;
  wire  _T_814; // @[NV_NVDLA_CSC_sg.scala 508:30:@1952.4]
  wire  _T_817; // @[NV_NVDLA_CSC_sg.scala 509:49:@1953.4]
  wire [6:0] _T_819; // @[NV_NVDLA_CSC_sg.scala 509:29:@1954.4]
  wire [6:0] _T_820; // @[NV_NVDLA_CSC_sg.scala 508:29:@1955.4]
  wire  _T_856; // @[NV_NVDLA_CSC_sg.scala 520:54:@1981.4]
  wire  _T_857; // @[NV_NVDLA_CSC_sg.scala 520:85:@1982.4]
  wire  _T_858; // @[NV_NVDLA_CSC_sg.scala 520:70:@1983.4]
  wire  _T_859; // @[NV_NVDLA_CSC_sg.scala 520:32:@1984.4]
  wire  _T_821; // @[NV_NVDLA_CSC_sg.scala 513:29:@1956.4]
  wire  _T_824; // @[NV_NVDLA_CSC_sg.scala 514:41:@1957.4]
  wire  _T_826; // @[NV_NVDLA_CSC_sg.scala 514:73:@1958.4]
  wire  _T_827; // @[NV_NVDLA_CSC_sg.scala 514:62:@1959.4]
  wire  _T_829; // @[NV_NVDLA_CSC_sg.scala 515:41:@1960.4]
  wire [5:0] _T_830; // @[NV_NVDLA_CSC_sg.scala 515:29:@1961.4]
  wire [5:0] _T_831; // @[NV_NVDLA_CSC_sg.scala 514:29:@1962.4]
  wire [5:0] _T_832; // @[NV_NVDLA_CSC_sg.scala 513:28:@1963.4]
  wire [6:0] _GEN_71; // @[NV_NVDLA_CSC_sg.scala 517:41:@1964.4]
  wire  _T_833; // @[NV_NVDLA_CSC_sg.scala 517:41:@1964.4]
  wire [7:0] _T_835; // @[NV_NVDLA_CSC_sg.scala 517:76:@1965.4]
  wire [7:0] _T_836; // @[NV_NVDLA_CSC_sg.scala 517:76:@1966.4]
  wire [6:0] _T_837; // @[NV_NVDLA_CSC_sg.scala 517:76:@1967.4]
  wire [6:0] _T_839; // @[NV_NVDLA_CSC_sg.scala 517:99:@1968.4]
  wire [6:0] _T_840; // @[NV_NVDLA_CSC_sg.scala 517:99:@1969.4]
  wire [5:0] _T_841; // @[NV_NVDLA_CSC_sg.scala 517:99:@1970.4]
  wire [6:0] _T_842; // @[NV_NVDLA_CSC_sg.scala 517:25:@1971.4]
  wire [5:0] _T_843; // @[NV_NVDLA_CSC_sg.scala 517:106:@1972.4]
  wire [6:0] _T_845; // @[NV_NVDLA_CSC_sg.scala 518:31:@1973.4]
  wire [6:0] _T_846; // @[NV_NVDLA_CSC_sg.scala 518:31:@1974.4]
  wire [5:0] _T_847; // @[NV_NVDLA_CSC_sg.scala 518:31:@1975.4]
  wire  _T_848; // @[NV_NVDLA_CSC_sg.scala 519:39:@1976.4]
  wire [5:0] _T_852; // @[NV_NVDLA_CSC_sg.scala 519:70:@1978.4]
  wire [5:0] _T_853; // @[NV_NVDLA_CSC_sg.scala 519:24:@1979.4]
  wire [6:0] _GEN_54; // @[NV_NVDLA_CSC_sg.scala 525:26:@1995.4]
  wire [6:0] _GEN_55; // @[NV_NVDLA_CSC_sg.scala 525:26:@1995.4]
  wire [17:0] _GEN_57; // @[NV_NVDLA_CSC_sg.scala 535:23:@2005.4]
  reg  _T_873; // @[NV_NVDLA_CSC_sg.scala 549:61:@2013.4]
  reg [31:0] _RAND_63;
  reg [2:0] _T_875; // @[NV_NVDLA_CSC_sg.scala 550:58:@2014.4]
  reg [31:0] _RAND_64;
  wire [3:0] _T_879; // @[NV_NVDLA_CSC_sg.scala 559:29:@2020.4]
  wire  _T_880; // @[NV_NVDLA_CSC_sg.scala 560:43:@2021.4]
  wire [8:0] _T_882; // @[NV_NVDLA_CSC_sg.scala 560:29:@2022.4]
  wire  _T_886; // @[NV_NVDLA_CSC_sg.scala 563:24:@2027.4]
  wire [8:0] _GEN_72; // @[NV_NVDLA_CSC_sg.scala 564:34:@2029.6]
  wire [9:0] _T_887; // @[NV_NVDLA_CSC_sg.scala 564:34:@2029.6]
  wire [8:0] _T_888; // @[NV_NVDLA_CSC_sg.scala 564:34:@2030.6]
  wire [9:0] _T_889; // @[NV_NVDLA_CSC_sg.scala 564:51:@2031.6]
  wire [9:0] _T_890; // @[NV_NVDLA_CSC_sg.scala 564:51:@2032.6]
  wire [8:0] _T_891; // @[NV_NVDLA_CSC_sg.scala 564:51:@2033.6]
  wire [8:0] _GEN_59; // @[NV_NVDLA_CSC_sg.scala 563:37:@2028.4]
  wire  _T_892; // @[NV_NVDLA_CSC_sg.scala 570:31:@2036.4]
  wire  _T_894; // @[NV_NVDLA_CSC_sg.scala 570:49:@2038.4]
  wire  _T_895; // @[NV_NVDLA_CSC_sg.scala 571:37:@2039.4]
  wire  _T_896; // @[NV_NVDLA_CSC_sg.scala 571:58:@2040.4]
  wire  _T_897; // @[NV_NVDLA_CSC_sg.scala 571:80:@2041.4]
  wire  _T_898; // @[NV_NVDLA_CSC_sg.scala 571:55:@2042.4]
  wire  _T_900; // @[NV_NVDLA_CSC_sg.scala 571:113:@2043.4]
  wire  _T_901; // @[NV_NVDLA_CSC_sg.scala 571:98:@2044.4]
  wire [13:0] _T_903; // @[NV_NVDLA_CSC_sg.scala 572:29:@2045.4]
  wire [13:0] _T_905; // @[NV_NVDLA_CSC_sg.scala 573:58:@2046.4]
  wire [13:0] _T_906; // @[NV_NVDLA_CSC_sg.scala 573:29:@2047.4]
  wire  _T_908; // @[NV_NVDLA_CSC_sg.scala 574:30:@2049.4]
  wire  _T_909; // @[NV_NVDLA_CSC_sg.scala 574:59:@2050.4]
  wire  _T_911; // @[NV_NVDLA_CSC_sg.scala 575:56:@2052.4]
  wire  _T_912; // @[NV_NVDLA_CSC_sg.scala 575:54:@2053.4]
  wire  _T_913; // @[NV_NVDLA_CSC_sg.scala 575:80:@2054.4]
  wire [13:0] _T_915; // @[NV_NVDLA_CSC_sg.scala 576:30:@2055.4]
  wire [12:0] _T_917; // @[Cat.scala 30:58:@2056.4]
  wire [13:0] _T_919; // @[NV_NVDLA_CSC_sg.scala 577:81:@2057.4]
  wire [13:0] _T_920; // @[NV_NVDLA_CSC_sg.scala 577:30:@2058.4]
  wire  _T_921; // @[NV_NVDLA_CSC_sg.scala 579:26:@2059.4]
  wire  _T_922; // @[NV_NVDLA_CSC_sg.scala 579:40:@2060.4]
  wire  _T_923; // @[NV_NVDLA_CSC_sg.scala 579:60:@2061.4]
  wire [14:0] _T_925; // @[NV_NVDLA_CSC_sg.scala 580:75:@2063.6]
  wire [13:0] _T_926; // @[NV_NVDLA_CSC_sg.scala 580:75:@2064.6]
  wire [14:0] _T_927; // @[NV_NVDLA_CSC_sg.scala 580:92:@2065.6]
  wire [14:0] _T_928; // @[NV_NVDLA_CSC_sg.scala 580:92:@2066.6]
  wire [13:0] _T_929; // @[NV_NVDLA_CSC_sg.scala 580:92:@2067.6]
  wire [13:0] _T_930; // @[NV_NVDLA_CSC_sg.scala 580:26:@2068.6]
  wire [13:0] _GEN_60; // @[NV_NVDLA_CSC_sg.scala 579:88:@2062.4]
  wire  _T_931; // @[NV_NVDLA_CSC_sg.scala 582:25:@2071.4]
  wire  _T_932; // @[NV_NVDLA_CSC_sg.scala 582:38:@2072.4]
  wire  _T_933; // @[NV_NVDLA_CSC_sg.scala 582:57:@2073.4]
  wire [14:0] _GEN_73; // @[NV_NVDLA_CSC_sg.scala 583:75:@2075.6]
  wire [15:0] _T_935; // @[NV_NVDLA_CSC_sg.scala 583:75:@2075.6]
  wire [14:0] _T_936; // @[NV_NVDLA_CSC_sg.scala 583:75:@2076.6]
  wire [14:0] _GEN_74; // @[NV_NVDLA_CSC_sg.scala 583:93:@2077.6]
  wire [15:0] _T_937; // @[NV_NVDLA_CSC_sg.scala 583:93:@2077.6]
  wire [15:0] _T_938; // @[NV_NVDLA_CSC_sg.scala 583:93:@2078.6]
  wire [14:0] _T_939; // @[NV_NVDLA_CSC_sg.scala 583:93:@2079.6]
  wire [14:0] _T_940; // @[NV_NVDLA_CSC_sg.scala 583:27:@2080.6]
  wire [14:0] _GEN_61; // @[NV_NVDLA_CSC_sg.scala 582:84:@2074.4]
  reg  _T_943; // @[NV_NVDLA_CSC_sg.scala 586:66:@2083.4]
  reg [31:0] _RAND_65;
  reg  _T_946; // @[NV_NVDLA_CSC_sg.scala 587:66:@2086.4]
  reg [31:0] _RAND_66;
  NV_NVDLA_fifo NV_NVDLA_fifo ( // @[NV_NVDLA_CSC_sg.scala 433:28:@1885.4]
    .clock(NV_NVDLA_fifo_clock),
    .reset(NV_NVDLA_fifo_reset),
    .io_clk(NV_NVDLA_fifo_io_clk),
    .io_wr_pvld(NV_NVDLA_fifo_io_wr_pvld),
    .io_wr_prdy(NV_NVDLA_fifo_io_wr_prdy),
    .io_wr_pd(NV_NVDLA_fifo_io_wr_pd),
    .io_wr_empty(NV_NVDLA_fifo_io_wr_empty),
    .io_rd_pvld(NV_NVDLA_fifo_io_rd_pvld),
    .io_rd_prdy(NV_NVDLA_fifo_io_rd_prdy),
    .io_rd_pd(NV_NVDLA_fifo_io_rd_pd)
  );
  NV_NVDLA_fifo_1 NV_NVDLA_fifo_1 ( // @[NV_NVDLA_CSC_sg.scala 446:27:@1896.4]
    .clock(NV_NVDLA_fifo_1_clock),
    .reset(NV_NVDLA_fifo_1_reset),
    .io_clk(NV_NVDLA_fifo_1_io_clk),
    .io_wr_pvld(NV_NVDLA_fifo_1_io_wr_pvld),
    .io_wr_prdy(NV_NVDLA_fifo_1_io_wr_prdy),
    .io_wr_pd(NV_NVDLA_fifo_1_io_wr_pd),
    .io_wr_empty(NV_NVDLA_fifo_1_io_wr_empty),
    .io_rd_pvld(NV_NVDLA_fifo_1_io_rd_pvld),
    .io_rd_prdy(NV_NVDLA_fifo_1_io_rd_prdy),
    .io_rd_pd(NV_NVDLA_fifo_1_io_rd_pd)
  );
  assign _T_145 = 2'h0 == _T_142; // @[Conditional.scala 37:30:@1416.4]
  assign _T_209 = _T_165 != io_reg2dp_data_bank; // @[NV_NVDLA_CSC_sg.scala 138:43:@1478.4]
  assign _T_210 = _T_168 != io_reg2dp_weight_bank; // @[NV_NVDLA_CSC_sg.scala 139:44:@1479.4]
  assign _T_211 = _T_209 | _T_210; // @[NV_NVDLA_CSC_sg.scala 140:38:@1480.4]
  assign _T_146 = io_reg2dp_op_en & _T_211; // @[NV_NVDLA_CSC_sg.scala 98:31:@1418.6]
  assign _GEN_0 = io_reg2dp_op_en ? 2'h2 : 2'h0; // @[NV_NVDLA_CSC_sg.scala 99:37:@1423.8]
  assign _GEN_1 = _T_146 ? 2'h1 : _GEN_0; // @[NV_NVDLA_CSC_sg.scala 98:47:@1419.6]
  assign _T_147 = 2'h1 == _T_142; // @[Conditional.scala 37:30:@1428.6]
  assign _T_241 = _T_142 == 2'h1; // @[NV_NVDLA_CSC_sg.scala 160:30:@1512.4]
  assign _T_212 = _T_171 ^ _T_174; // @[NV_NVDLA_CSC_sg.scala 141:51:@1482.4]
  assign _T_213 = ~ _T_212; // @[NV_NVDLA_CSC_sg.scala 141:34:@1483.4]
  assign _T_214 = _T_241 & _T_213; // @[NV_NVDLA_CSC_sg.scala 141:32:@1484.4]
  assign _T_215 = _T_180 ^ _T_183; // @[NV_NVDLA_CSC_sg.scala 141:87:@1485.4]
  assign _T_216 = ~ _T_215; // @[NV_NVDLA_CSC_sg.scala 141:71:@1486.4]
  assign _T_217 = _T_214 & _T_216; // @[NV_NVDLA_CSC_sg.scala 141:69:@1487.4]
  assign _GEN_2 = _T_217 ? 2'h2 : 2'h0; // @[NV_NVDLA_CSC_sg.scala 102:29:@1430.8]
  assign _T_148 = 2'h2 == _T_142; // @[Conditional.scala 37:30:@1435.8]
  assign _T_154 = NV_NVDLA_fifo_io_rd_pvld; // @[NV_NVDLA_CSC_sg.scala 116:27:@1452.4 NV_NVDLA_CSC_sg.scala 441:17:@1893.4]
  assign _T_204 = ~ _T_154; // @[NV_NVDLA_CSC_sg.scala 137:22:@1472.4]
  assign _T_160 = NV_NVDLA_fifo_1_io_rd_pvld; // @[NV_NVDLA_CSC_sg.scala 119:26:@1455.4 NV_NVDLA_CSC_sg.scala 454:16:@1904.4]
  assign _T_205 = ~ _T_160; // @[NV_NVDLA_CSC_sg.scala 137:37:@1473.4]
  assign _T_206 = _T_204 & _T_205; // @[NV_NVDLA_CSC_sg.scala 137:35:@1474.4]
  assign _T_156 = NV_NVDLA_fifo_io_wr_empty; // @[NV_NVDLA_CSC_sg.scala 117:30:@1453.4 NV_NVDLA_CSC_sg.scala 444:20:@1895.4]
  assign _T_207 = _T_206 & _T_156; // @[NV_NVDLA_CSC_sg.scala 137:49:@1475.4]
  assign _T_162 = NV_NVDLA_fifo_1_io_wr_empty; // @[NV_NVDLA_CSC_sg.scala 120:29:@1456.4 NV_NVDLA_CSC_sg.scala 457:19:@1906.4]
  assign _T_208 = _T_207 & _T_162; // @[NV_NVDLA_CSC_sg.scala 137:66:@1476.4]
  assign _T_149 = _T_131 & _T_208; // @[NV_NVDLA_CSC_sg.scala 105:26:@1437.10]
  assign _T_150 = ~ _T_136; // @[NV_NVDLA_CSC_sg.scala 105:44:@1438.10]
  assign _T_151 = _T_149 & _T_150; // @[NV_NVDLA_CSC_sg.scala 105:42:@1439.10]
  assign _GEN_3 = _T_151 ? 2'h3 : 2'h0; // @[NV_NVDLA_CSC_sg.scala 105:54:@1440.10]
  assign _GEN_6 = _T_148 ? _GEN_3 : 2'h0; // @[Conditional.scala 39:67:@1436.8]
  assign _GEN_7 = _T_147 ? _GEN_2 : _GEN_6; // @[Conditional.scala 39:67:@1429.6]
  assign _GEN_8 = _T_145 ? _GEN_1 : _GEN_7; // @[Conditional.scala 40:58:@1417.4]
  assign _T_243 = _T_142 == 2'h3; // @[NV_NVDLA_CSC_sg.scala 162:27:@1515.4]
  assign _T_218 = ~ _T_243; // @[NV_NVDLA_CSC_sg.scala 144:26:@1490.6]
  assign _T_244 = _GEN_8 == 2'h3; // @[NV_NVDLA_CSC_sg.scala 163:31:@1517.4]
  assign _T_219 = _T_218 & _T_244; // @[NV_NVDLA_CSC_sg.scala 144:35:@1491.6]
  assign _T_221 = _T_201 - 8'h1; // @[NV_NVDLA_CSC_sg.scala 144:74:@1492.6]
  assign _T_222 = $unsigned(_T_221); // @[NV_NVDLA_CSC_sg.scala 144:74:@1493.6]
  assign _T_223 = _T_222[7:0]; // @[NV_NVDLA_CSC_sg.scala 144:74:@1494.6]
  assign _T_224 = _T_219 ? _T_198 : _T_223; // @[NV_NVDLA_CSC_sg.scala 144:25:@1495.6]
  assign _GEN_9 = _T_244 ? _T_224 : _T_201; // @[NV_NVDLA_CSC_sg.scala 143:22:@1489.4]
  assign _T_861 = _T_799 == 6'h0; // @[NV_NVDLA_CSC_sg.scala 521:45:@1986.4]
  assign _T_862 = _T_154 & _T_861; // @[NV_NVDLA_CSC_sg.scala 521:34:@1987.4]
  assign _T_748 = NV_NVDLA_fifo_io_rd_pd[30:0]; // @[NV_NVDLA_CSC_sg.scala 463:34:@1908.4]
  assign _T_757 = _T_748[27]; // @[NV_NVDLA_CSC_sg.scala 474:40:@1917.4]
  assign _T_883 = ~ _T_757; // @[NV_NVDLA_CSC_sg.scala 561:21:@2023.4]
  assign _T_877 = {2'h0,_T_191}; // @[Cat.scala 30:58:@2019.4]
  assign _T_884 = _T_870 >= _T_877; // @[NV_NVDLA_CSC_sg.scala 561:55:@2024.4]
  assign _T_885 = _T_883 | _T_884; // @[NV_NVDLA_CSC_sg.scala 561:41:@2025.4]
  assign _T_863 = _T_862 & _T_885; // @[NV_NVDLA_CSC_sg.scala 521:54:@1988.4]
  assign _T_747 = NV_NVDLA_fifo_io_rd_pd[32:31]; // @[NV_NVDLA_CSC_sg.scala 462:35:@1907.4]
  assign _T_749 = NV_NVDLA_fifo_1_io_rd_pd[19:18]; // @[NV_NVDLA_CSC_sg.scala 464:33:@1909.4]
  assign _T_864 = _T_747 != _T_749; // @[NV_NVDLA_CSC_sg.scala 521:85:@1989.4]
  assign _T_866 = _T_864 | _T_205; // @[NV_NVDLA_CSC_sg.scala 521:101:@1991.4]
  assign _T_867 = _T_863 & _T_866; // @[NV_NVDLA_CSC_sg.scala 521:69:@1992.4]
  assign _T_225 = _T_154 & _T_867; // @[NV_NVDLA_CSC_sg.scala 148:22:@1500.4]
  assign _T_759 = _T_748[29]; // @[NV_NVDLA_CSC_sg.scala 476:35:@1919.4]
  assign _T_226 = _T_225 & _T_759; // @[NV_NVDLA_CSC_sg.scala 148:38:@1501.4]
  assign _T_228 = _T_191 + 7'h30; // @[NV_NVDLA_CSC_sg.scala 149:41:@1503.6]
  assign _GEN_10 = _T_226 ? _T_228 : _T_198; // @[NV_NVDLA_CSC_sg.scala 148:57:@1502.4]
  assign _T_238 = _T_142 == 2'h0; // @[NV_NVDLA_CSC_sg.scala 158:49:@1509.4]
  assign _T_239 = io_reg2dp_op_en & _T_238; // @[NV_NVDLA_CSC_sg.scala 158:36:@1510.4]
  assign _T_242 = _T_142 == 2'h2; // @[NV_NVDLA_CSC_sg.scala 161:33:@1514.4]
  assign _T_245 = _GEN_8 == 2'h1; // @[NV_NVDLA_CSC_sg.scala 164:37:@1519.4]
  assign _T_250 = _T_242 ? 2'h2 : 2'h3; // @[NV_NVDLA_CSC_sg.scala 165:90:@1520.4]
  assign _T_251 = _T_241 ? 2'h1 : _T_250; // @[NV_NVDLA_CSC_sg.scala 165:55:@1521.4]
  assign _T_312 = io_reg2dp_conv_mode == 1'h0; // @[NV_NVDLA_CSC_sg.scala 199:40:@1568.4]
  assign _T_313 = _T_312 & io_reg2dp_datain_format; // @[NV_NVDLA_CSC_sg.scala 200:26:@1569.4]
  assign _T_314 = ~ io_reg2dp_datain_format; // @[NV_NVDLA_CSC_sg.scala 201:27:@1570.4]
  assign _T_315 = _T_312 & _T_314; // @[NV_NVDLA_CSC_sg.scala 201:25:@1571.4]
  assign _T_318 = {_T_313,1'h0,_T_315}; // @[Cat.scala 30:58:@1573.4]
  assign _T_253 = _T_237 != _T_318; // @[NV_NVDLA_CSC_sg.scala 166:37:@1524.4]
  assign _T_255 = _T_201 == 8'h1; // @[NV_NVDLA_CSC_sg.scala 168:53:@1525.4]
  assign _T_256 = _T_243 & _T_255; // @[NV_NVDLA_CSC_sg.scala 168:39:@1526.4]
  assign _T_260 = _T_245 & _T_209; // @[NV_NVDLA_CSC_sg.scala 169:43:@1530.4]
  assign _T_262 = ~ _T_245; // @[NV_NVDLA_CSC_sg.scala 169:85:@1531.4]
  assign _T_264 = _T_262 ? 1'h0 : _T_174; // @[NV_NVDLA_CSC_sg.scala 169:83:@1532.4]
  assign _T_265 = _T_260 ? 1'h1 : _T_264; // @[NV_NVDLA_CSC_sg.scala 169:27:@1533.4]
  assign _T_269 = _T_262 ? 1'h0 : _T_183; // @[NV_NVDLA_CSC_sg.scala 170:64:@1536.4]
  assign _T_270 = _T_245 ? 1'h1 : _T_269; // @[NV_NVDLA_CSC_sg.scala 170:26:@1537.4]
  assign _T_271 = _T_241 & _T_177; // @[NV_NVDLA_CSC_sg.scala 171:39:@1539.4]
  assign _T_275 = _T_262 ? 1'h0 : _T_171; // @[NV_NVDLA_CSC_sg.scala 171:79:@1541.4]
  assign _T_276 = _T_271 ? 1'h1 : _T_275; // @[NV_NVDLA_CSC_sg.scala 171:27:@1542.4]
  assign _T_277 = _T_241 & _T_186; // @[NV_NVDLA_CSC_sg.scala 172:38:@1544.4]
  assign _T_281 = _T_262 ? 1'h0 : _T_180; // @[NV_NVDLA_CSC_sg.scala 172:77:@1546.4]
  assign _T_282 = _T_277 ? 1'h1 : _T_281; // @[NV_NVDLA_CSC_sg.scala 172:26:@1547.4]
  assign _T_308 = io_reg2dp_weight_kernel + 13'h1; // @[NV_NVDLA_CSC_sg.scala 190:49:@1562.6]
  assign _GEN_11 = io_dp2reg_done ? io_reg2dp_data_bank : _T_165; // @[NV_NVDLA_CSC_sg.scala 186:25:@1558.4]
  assign _GEN_12 = io_dp2reg_done ? io_reg2dp_weight_bank : _T_168; // @[NV_NVDLA_CSC_sg.scala 186:25:@1558.4]
  assign _GEN_13 = io_dp2reg_done ? _T_296 : _T_289; // @[NV_NVDLA_CSC_sg.scala 186:25:@1558.4]
  assign _GEN_14 = io_dp2reg_done ? _T_308 : _T_303; // @[NV_NVDLA_CSC_sg.scala 186:25:@1558.4]
  assign _GEN_15 = io_dp2reg_done ? io_reg2dp_skip_weight_rls : _T_306; // @[NV_NVDLA_CSC_sg.scala 186:25:@1558.4]
  assign _GEN_16 = io_dp2reg_done ? _T_318 : _T_237; // @[NV_NVDLA_CSC_sg.scala 186:25:@1558.4]
  assign _T_392 = 9'h9 << io_reg2dp_y_extension; // @[NV_NVDLA_CSC_sg.scala 221:44:@1596.4]
  assign _T_393 = _T_392[5:3]; // @[NV_NVDLA_CSC_sg.scala 221:69:@1597.4]
  assign _T_395 = io_reg2dp_datain_height_ext + 13'h1; // @[NV_NVDLA_CSC_sg.scala 224:55:@1599.6]
  assign _T_397 = io_reg2dp_dataout_width + 13'h1; // @[NV_NVDLA_CSC_sg.scala 225:64:@1601.6]
  assign _T_399 = io_reg2dp_atomics + 21'h1; // @[NV_NVDLA_CSC_sg.scala 225:90:@1602.6]
  assign _T_400 = _T_313 ? {{8'd0}, _T_397} : _T_399; // @[NV_NVDLA_CSC_sg.scala 225:31:@1603.6]
  assign _T_403 = _T_313 ? 5'h0 : io_reg2dp_weight_width_ext; // @[NV_NVDLA_CSC_sg.scala 227:32:@1606.6]
  assign _T_405 = io_reg2dp_weight_channel_ext + 13'h1; // @[NV_NVDLA_CSC_sg.scala 229:56:@1609.6]
  assign _T_406 = io_reg2dp_weight_kernel[12:5]; // @[NV_NVDLA_CSC_sg.scala 230:49:@1611.6]
  assign _T_408 = _T_406 + 8'h1; // @[NV_NVDLA_CSC_sg.scala 230:71:@1612.6]
  assign _T_409 = _T_393[0]; // @[NV_NVDLA_CSC_sg.scala 232:44:@1615.6]
  assign _T_411 = _T_393[1]; // @[NV_NVDLA_CSC_sg.scala 233:44:@1616.6]
  assign _T_413 = io_reg2dp_weight_height_ext[0]; // @[NV_NVDLA_CSC_sg.scala 233:98:@1617.6]
  assign _T_414 = {1'h0,_T_413}; // @[Cat.scala 30:58:@1618.6]
  assign _T_415 = io_reg2dp_weight_height_ext[1:0]; // @[NV_NVDLA_CSC_sg.scala 234:55:@1619.6]
  assign _T_416 = _T_411 ? _T_414 : _T_415; // @[NV_NVDLA_CSC_sg.scala 233:29:@1620.6]
  assign _T_417 = _T_409 ? 2'h0 : _T_416; // @[NV_NVDLA_CSC_sg.scala 232:29:@1621.6]
  assign _T_419 = io_reg2dp_rls_slices + 12'h1; // @[NV_NVDLA_CSC_sg.scala 235:44:@1623.6]
  assign _T_420 = io_reg2dp_rls_slices + 12'h1; // @[NV_NVDLA_CSC_sg.scala 235:44:@1624.6]
  assign _GEN_62 = {{1'd0}, io_reg2dp_rls_slices}; // @[NV_NVDLA_CSC_sg.scala 236:116:@1627.6]
  assign _T_423 = io_reg2dp_datain_height_ext - _GEN_62; // @[NV_NVDLA_CSC_sg.scala 236:116:@1627.6]
  assign _T_424 = $unsigned(_T_423); // @[NV_NVDLA_CSC_sg.scala 236:116:@1628.6]
  assign _T_425 = io_reg2dp_skip_data_rls ? _T_395 : _T_424; // @[NV_NVDLA_CSC_sg.scala 236:26:@1629.6]
  assign _T_428 = _T_313 ? 7'h40 : 7'h20; // @[NV_NVDLA_CSC_sg.scala 240:27:@1632.6]
  assign _GEN_17 = _T_239 ? _T_395 : _T_326; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  assign _GEN_18 = _T_239 ? _T_400 : _T_333; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  assign _GEN_20 = _T_239 ? _T_403 : _T_347; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  assign _GEN_21 = _T_239 ? io_reg2dp_weight_height_ext : _T_354; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  assign _GEN_22 = _T_239 ? _T_405 : _T_361; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  assign _GEN_23 = _T_239 ? {{1'd0}, _T_408} : _T_368; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  assign _GEN_24 = _T_239 ? _T_393 : _T_371; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  assign _GEN_25 = _T_239 ? {{1'd0}, _T_417} : _T_374; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  assign _GEN_26 = _T_239 ? {{2'd0}, _T_420} : _T_381; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  assign _GEN_27 = _T_239 ? _T_425 : _T_296; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  assign _GEN_28 = _T_239 ? _T_313 : _T_384; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  assign _GEN_29 = _T_239 ? _T_428 : {{1'd0}, _T_387}; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  assign _GEN_30 = _T_239 ? 7'h40 : _T_390; // @[NV_NVDLA_CSC_sg.scala 223:19:@1598.4]
  assign _T_600 = _T_593 >= _T_326; // @[NV_NVDLA_CSC_sg.scala 337:38:@1750.4]
  assign _T_451 = _T_449 + 10'h1; // @[NV_NVDLA_CSC_sg.scala 258:41:@1648.4]
  assign _T_452 = _T_449 + 10'h1; // @[NV_NVDLA_CSC_sg.scala 258:41:@1649.4]
  assign _T_453 = _T_452 == _T_368; // @[NV_NVDLA_CSC_sg.scala 259:40:@1650.4]
  assign _T_454 = ~ _T_453; // @[NV_NVDLA_CSC_sg.scala 260:26:@1652.4]
  assign _T_456 = io_reg2dp_weight_kernel[4:0]; // @[NV_NVDLA_CSC_sg.scala 260:87:@1653.4]
  assign _T_458 = _T_456 + 5'h1; // @[NV_NVDLA_CSC_sg.scala 260:110:@1654.4]
  assign _T_459 = _T_454 ? 6'h20 : _T_458; // @[NV_NVDLA_CSC_sg.scala 260:25:@1655.4]
  assign _GEN_63 = {{8'd0}, _T_459}; // @[NV_NVDLA_CSC_sg.scala 338:49:@1751.4]
  assign _T_601 = _T_596 + _GEN_63; // @[NV_NVDLA_CSC_sg.scala 338:49:@1751.4]
  assign _T_602 = _T_596 + _GEN_63; // @[NV_NVDLA_CSC_sg.scala 338:49:@1752.4]
  assign _GEN_64 = {{1'd0}, _T_602}; // @[NV_NVDLA_CSC_sg.scala 339:46:@1753.4]
  assign _T_603 = _GEN_64 <= _T_599; // @[NV_NVDLA_CSC_sg.scala 339:46:@1753.4]
  assign _T_615 = _T_600 & _T_603; // @[NV_NVDLA_CSC_sg.scala 350:37:@1765.4]
  assign _T_616 = _T_242 & _T_615; // @[NV_NVDLA_CSC_sg.scala 351:30:@1766.4]
  assign _T_617 = ~ _T_131; // @[NV_NVDLA_CSC_sg.scala 351:45:@1767.4]
  assign _T_618 = _T_616 & _T_617; // @[NV_NVDLA_CSC_sg.scala 351:43:@1768.4]
  assign _T_611 = NV_NVDLA_fifo_io_wr_prdy; // @[NV_NVDLA_CSC_sg.scala 346:30:@1762.4 NV_NVDLA_CSC_sg.scala 439:20:@1891.4]
  assign _T_613 = NV_NVDLA_fifo_1_io_wr_prdy; // @[NV_NVDLA_CSC_sg.scala 347:29:@1763.4 NV_NVDLA_CSC_sg.scala 452:19:@1902.4]
  assign _T_614 = _T_611 & _T_613; // @[NV_NVDLA_CSC_sg.scala 349:42:@1764.4]
  assign _T_620 = _T_150 | _T_614; // @[NV_NVDLA_CSC_sg.scala 351:69:@1770.4]
  assign _T_621 = _T_618 & _T_620; // @[NV_NVDLA_CSC_sg.scala 351:57:@1771.4]
  assign _T_570 = _T_554 == _T_347; // @[NV_NVDLA_CSC_sg.scala 315:38:@1729.4]
  assign _GEN_65 = {{2'd0}, _T_371}; // @[NV_NVDLA_CSC_sg.scala 314:47:@1728.4]
  assign _T_569 = _T_561 + _GEN_65; // @[NV_NVDLA_CSC_sg.scala 314:47:@1728.4]
  assign _GEN_66 = {{1'd0}, _T_354}; // @[NV_NVDLA_CSC_sg.scala 316:42:@1730.4]
  assign _T_571 = _T_569 > _GEN_66; // @[NV_NVDLA_CSC_sg.scala 316:42:@1730.4]
  assign _T_580 = _T_570 & _T_571; // @[NV_NVDLA_CSC_sg.scala 322:35:@1736.4]
  assign _T_634 = _T_621 & _T_580; // @[NV_NVDLA_CSC_sg.scala 358:28:@1790.4]
  assign _T_526 = _T_524 + 14'h40; // @[NV_NVDLA_CSC_sg.scala 298:45:@1705.4]
  assign _T_527 = _T_524 + 14'h40; // @[NV_NVDLA_CSC_sg.scala 298:45:@1706.4]
  assign _T_528 = _T_527 >= _T_361; // @[NV_NVDLA_CSC_sg.scala 299:47:@1707.4]
  assign _T_635 = _T_634 & _T_528; // @[NV_NVDLA_CSC_sg.scala 358:44:@1791.4]
  assign _GEN_67 = {{15'd0}, _T_390}; // @[NV_NVDLA_CSC_sg.scala 280:47:@1680.4]
  assign _T_494 = _T_489 + _GEN_67; // @[NV_NVDLA_CSC_sg.scala 280:47:@1680.4]
  assign _T_495 = _T_489 + _GEN_67; // @[NV_NVDLA_CSC_sg.scala 280:47:@1681.4]
  assign _T_497 = _T_495 >= _T_333; // @[NV_NVDLA_CSC_sg.scala 282:49:@1683.4]
  assign _T_636 = _T_635 & _T_497; // @[NV_NVDLA_CSC_sg.scala 358:62:@1792.4]
  assign _T_472 = ~ _T_384; // @[NV_NVDLA_CSC_sg.scala 270:24:@1664.4]
  assign _T_473 = _T_469 == io_reg2dp_dataout_height; // @[NV_NVDLA_CSC_sg.scala 270:55:@1665.4]
  assign _T_474 = _T_472 | _T_473; // @[NV_NVDLA_CSC_sg.scala 270:35:@1666.4]
  assign _T_637 = _T_636 & _T_474; // @[NV_NVDLA_CSC_sg.scala 358:79:@1793.4]
  assign _T_638 = _T_637 & _T_453; // @[NV_NVDLA_CSC_sg.scala 358:94:@1794.4]
  assign _T_436 = _T_239 | _T_638; // @[NV_NVDLA_CSC_sg.scala 251:19:@1639.4]
  assign _T_439 = _T_453 ? 1'h1 : _T_131; // @[NV_NVDLA_CSC_sg.scala 252:48:@1641.6]
  assign _T_440 = _T_239 ? 1'h0 : _T_439; // @[NV_NVDLA_CSC_sg.scala 252:25:@1642.6]
  assign _GEN_31 = _T_436 ? _T_440 : _T_131; // @[NV_NVDLA_CSC_sg.scala 251:33:@1640.4]
  assign _T_460 = _T_239 | _T_637; // @[NV_NVDLA_CSC_sg.scala 262:19:@1656.4]
  assign _T_462 = _T_239 ? 10'h0 : _T_452; // @[NV_NVDLA_CSC_sg.scala 263:27:@1658.6]
  assign _GEN_32 = _T_460 ? _T_462 : _T_449; // @[NV_NVDLA_CSC_sg.scala 262:33:@1657.4]
  assign _T_626 = _T_384 & _T_621; // @[NV_NVDLA_CSC_sg.scala 356:29:@1780.4]
  assign _T_627 = _T_626 & _T_580; // @[NV_NVDLA_CSC_sg.scala 356:39:@1781.4]
  assign _T_628 = _T_627 & _T_528; // @[NV_NVDLA_CSC_sg.scala 356:55:@1782.4]
  assign _T_629 = _T_628 & _T_497; // @[NV_NVDLA_CSC_sg.scala 356:73:@1783.4]
  assign _T_475 = _T_239 | _T_629; // @[NV_NVDLA_CSC_sg.scala 271:19:@1667.4]
  assign _T_479 = _T_469 + 13'h1; // @[NV_NVDLA_CSC_sg.scala 274:47:@1669.6]
  assign _T_480 = _T_469 + 13'h1; // @[NV_NVDLA_CSC_sg.scala 274:47:@1670.6]
  assign _T_481 = _T_474 ? 13'h0 : _T_480; // @[NV_NVDLA_CSC_sg.scala 273:32:@1671.6]
  assign _T_482 = _T_239 ? 13'h0 : _T_481; // @[NV_NVDLA_CSC_sg.scala 272:32:@1672.6]
  assign _GEN_33 = _T_475 ? _T_482 : _T_469; // @[NV_NVDLA_CSC_sg.scala 271:32:@1668.4]
  assign _T_491 = {_T_390,1'h0}; // @[Cat.scala 30:58:@1677.4]
  assign _GEN_68 = {{14'd0}, _T_491}; // @[NV_NVDLA_CSC_sg.scala 279:46:@1678.4]
  assign _T_492 = _T_489 + _GEN_68; // @[NV_NVDLA_CSC_sg.scala 279:46:@1678.4]
  assign _T_493 = _T_489 + _GEN_68; // @[NV_NVDLA_CSC_sg.scala 279:46:@1679.4]
  assign _T_496 = _T_493 <= _T_333; // @[NV_NVDLA_CSC_sg.scala 281:49:@1682.4]
  assign _T_498 = _T_333 - _T_489; // @[NV_NVDLA_CSC_sg.scala 284:43:@1684.4]
  assign _T_499 = $unsigned(_T_498); // @[NV_NVDLA_CSC_sg.scala 284:43:@1685.4]
  assign _T_500 = _T_499[21:0]; // @[NV_NVDLA_CSC_sg.scala 284:43:@1686.4]
  assign _T_501 = _T_500[6:0]; // @[NV_NVDLA_CSC_sg.scala 284:60:@1687.4]
  assign _T_502 = _T_497 ? _T_501 : {{1'd0}, _T_387}; // @[NV_NVDLA_CSC_sg.scala 285:59:@1688.4]
  assign _T_503 = _T_496 ? _T_390 : _T_502; // @[NV_NVDLA_CSC_sg.scala 285:25:@1689.4]
  assign _T_506 = _T_239 | _T_635; // @[NV_NVDLA_CSC_sg.scala 288:19:@1691.4]
  assign _GEN_70 = {{16'd0}, _T_387}; // @[NV_NVDLA_CSC_sg.scala 292:41:@1695.6]
  assign _T_511 = _T_489 + _GEN_70; // @[NV_NVDLA_CSC_sg.scala 292:41:@1695.6]
  assign _T_512 = _T_489 + _GEN_70; // @[NV_NVDLA_CSC_sg.scala 292:41:@1696.6]
  assign _T_513 = _T_496 ? _T_495 : _T_512; // @[NV_NVDLA_CSC_sg.scala 291:29:@1697.6]
  assign _T_514 = _T_497 ? 22'h0 : _T_513; // @[NV_NVDLA_CSC_sg.scala 290:29:@1698.6]
  assign _T_515 = _T_239 ? 22'h0 : _T_514; // @[NV_NVDLA_CSC_sg.scala 289:29:@1699.6]
  assign _GEN_34 = _T_506 ? _T_515 : _T_489; // @[NV_NVDLA_CSC_sg.scala 288:34:@1692.4]
  assign _T_529 = ~ _T_528; // @[NV_NVDLA_CSC_sg.scala 301:27:@1708.4]
  assign _T_531 = io_reg2dp_weight_channel_ext[5:0]; // @[NV_NVDLA_CSC_sg.scala 301:93:@1709.4]
  assign _T_533 = _T_531 + 6'h1; // @[NV_NVDLA_CSC_sg.scala 301:117:@1710.4]
  assign _T_534 = _T_529 ? 7'h40 : _T_533; // @[NV_NVDLA_CSC_sg.scala 301:26:@1711.4]
  assign _T_535 = _T_239 | _T_634; // @[NV_NVDLA_CSC_sg.scala 303:19:@1712.4]
  assign _T_546 = _T_528 ? 14'h0 : _T_527; // @[NV_NVDLA_CSC_sg.scala 304:63:@1716.6]
  assign _T_547 = _T_239 ? 14'h0 : _T_546; // @[NV_NVDLA_CSC_sg.scala 304:30:@1717.6]
  assign _GEN_35 = _T_535 ? _T_547 : _T_524; // @[NV_NVDLA_CSC_sg.scala 303:35:@1713.4]
  assign _T_567 = _T_554 + 5'h1; // @[NV_NVDLA_CSC_sg.scala 313:47:@1726.4]
  assign _T_568 = _T_554 + 5'h1; // @[NV_NVDLA_CSC_sg.scala 313:47:@1727.4]
  assign _T_572 = _T_371[2]; // @[NV_NVDLA_CSC_sg.scala 318:33:@1731.4]
  assign _T_574 = _T_371[1]; // @[NV_NVDLA_CSC_sg.scala 319:33:@1732.4]
  assign _T_577 = _T_574 ? 2'h1 : 2'h0; // @[NV_NVDLA_CSC_sg.scala 319:20:@1733.4]
  assign _T_578 = _T_572 ? 2'h3 : _T_577; // @[NV_NVDLA_CSC_sg.scala 318:20:@1734.4]
  assign _T_579 = _T_571 ? _T_374 : {{1'd0}, _T_578}; // @[NV_NVDLA_CSC_sg.scala 317:20:@1735.4]
  assign _T_581 = _T_239 | _T_621; // @[NV_NVDLA_CSC_sg.scala 324:19:@1737.4]
  assign _T_584 = _T_570 ? 5'h0 : _T_568; // @[NV_NVDLA_CSC_sg.scala 326:32:@1739.6]
  assign _T_585 = _T_239 ? 5'h0 : _T_584; // @[NV_NVDLA_CSC_sg.scala 325:31:@1740.6]
  assign _T_588 = _T_569[4:0]; // @[NV_NVDLA_CSC_sg.scala 330:48:@1742.6]
  assign _T_589 = _T_571 ? 5'h0 : _T_588; // @[NV_NVDLA_CSC_sg.scala 329:32:@1743.6]
  assign _T_590 = _T_239 ? 5'h0 : _T_589; // @[NV_NVDLA_CSC_sg.scala 328:31:@1744.6]
  assign _GEN_36 = _T_581 ? _T_585 : _T_554; // @[NV_NVDLA_CSC_sg.scala 324:29:@1738.4]
  assign _GEN_37 = _T_581 ? _T_590 : _T_561; // @[NV_NVDLA_CSC_sg.scala 324:29:@1738.4]
  assign _T_605 = _T_239 | _T_453; // @[NV_NVDLA_CSC_sg.scala 342:43:@1756.6]
  assign _T_606 = ~ io_reg2dp_skip_weight_rls; // @[NV_NVDLA_CSC_sg.scala 342:61:@1757.6]
  assign _T_607 = _T_605 | _T_606; // @[NV_NVDLA_CSC_sg.scala 342:59:@1758.6]
  assign _T_609 = _T_607 ? 14'h0 : _T_602; // @[NV_NVDLA_CSC_sg.scala 342:32:@1759.6]
  assign _GEN_38 = _T_460 ? _T_609 : _T_596; // @[NV_NVDLA_CSC_sg.scala 341:33:@1755.4]
  assign _T_639 = ~ _T_242; // @[NV_NVDLA_CSC_sg.scala 360:20:@1796.4]
  assign _T_642 = _T_615 & _T_617; // @[NV_NVDLA_CSC_sg.scala 360:57:@1798.4]
  assign _T_645 = _T_614 ? 1'h0 : _T_136; // @[NV_NVDLA_CSC_sg.scala 360:83:@1799.4]
  assign _T_646 = _T_642 ? 1'h1 : _T_645; // @[NV_NVDLA_CSC_sg.scala 360:45:@1800.4]
  assign _T_647 = _T_639 ? 1'h0 : _T_646; // @[NV_NVDLA_CSC_sg.scala 360:19:@1801.4]
  assign _T_687 = _T_654 + 2'h1; // @[NV_NVDLA_CSC_sg.scala 375:61:@1815.4]
  assign _T_688 = _T_654 + 2'h1; // @[NV_NVDLA_CSC_sg.scala 375:61:@1816.4]
  assign _T_689 = _T_239 ? 2'h3 : _T_688; // @[NV_NVDLA_CSC_sg.scala 375:24:@1817.4]
  assign _T_690 = _T_580 & _T_528; // @[NV_NVDLA_CSC_sg.scala 379:43:@1818.4]
  assign _T_692 = _T_690 & _T_497; // @[NV_NVDLA_CSC_sg.scala 380:59:@1820.4]
  assign _T_693 = _T_692 & _T_474; // @[NV_NVDLA_CSC_sg.scala 380:76:@1821.4]
  assign _T_697 = _T_693 & _T_453; // @[NV_NVDLA_CSC_sg.scala 381:91:@1825.4]
  assign _GEN_39 = _T_581 ? _T_689 : _T_654; // @[NV_NVDLA_CSC_sg.scala 383:29:@1827.4]
  assign _T_704 = ~ io_reg2dp_skip_data_rls; // @[NV_NVDLA_CSC_sg.scala 396:32:@1843.6]
  assign _T_705 = _T_704 & _T_697; // @[NV_NVDLA_CSC_sg.scala 396:57:@1844.6]
  assign _GEN_40 = _T_621 ? _T_554 : _T_657; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  assign _GEN_41 = _T_621 ? _T_561 : _T_660; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  assign _GEN_42 = _T_621 ? _T_534 : _T_663; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  assign _GEN_43 = _T_621 ? _T_503 : _T_666; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  assign _GEN_44 = _T_621 ? _T_579 : _T_669; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  assign _GEN_45 = _T_621 ? _T_580 : _T_672; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  assign _GEN_46 = _T_621 ? _T_690 : _T_675; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  assign _GEN_47 = _T_621 ? _T_693 : _T_678; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  assign _GEN_48 = _T_621 ? _T_697 : _T_681; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  assign _GEN_49 = _T_621 ? _T_705 : _T_684; // @[NV_NVDLA_CSC_sg.scala 386:18:@1833.4]
  assign _T_718 = _T_669[1:0]; // @[NV_NVDLA_CSC_sg.scala 406:42:@1851.4]
  assign _T_731 = {_T_684,_T_681,_T_678,_T_675,_T_672,_T_718,_T_666,_T_663,_T_660,_T_657}; // @[Cat.scala 30:58:@1864.4]
  assign _T_734 = _T_606 & _T_693; // @[NV_NVDLA_CSC_sg.scala 415:57:@1871.6]
  assign _GEN_50 = _T_621 ? {{1'd0}, _T_459} : _T_708; // @[NV_NVDLA_CSC_sg.scala 411:18:@1866.4]
  assign _GEN_51 = _T_621 ? _T_534 : _T_711; // @[NV_NVDLA_CSC_sg.scala 411:18:@1866.4]
  assign _GEN_52 = _T_621 ? _T_579 : _T_714; // @[NV_NVDLA_CSC_sg.scala 411:18:@1866.4]
  assign _GEN_53 = _T_621 ? _T_734 : _T_717; // @[NV_NVDLA_CSC_sg.scala 411:18:@1866.4]
  assign _T_735 = _T_714[1:0]; // @[NV_NVDLA_CSC_sg.scala 423:41:@1874.4]
  assign _T_736 = _T_708[5:0]; // @[NV_NVDLA_CSC_sg.scala 423:67:@1875.4]
  assign _T_741 = {_T_717,_T_678,_T_675,_T_735,_T_736,_T_711}; // @[Cat.scala 30:58:@1880.4]
  assign _T_750 = NV_NVDLA_fifo_1_io_rd_pd[17:0]; // @[NV_NVDLA_CSC_sg.scala 465:32:@1910.4]
  assign _T_754 = _T_748[23:17]; // @[NV_NVDLA_CSC_sg.scala 471:42:@1914.4]
  assign _T_762 = _T_750[12:7]; // @[NV_NVDLA_CSC_sg.scala 481:38:@1923.4]
  assign _T_774 = io_reg2dp_y_extension == 2'h2; // @[NV_NVDLA_CSC_sg.scala 492:61:@1932.4]
  assign _T_776 = _T_754 + 7'h3; // @[NV_NVDLA_CSC_sg.scala 492:106:@1933.4]
  assign _T_778 = _T_776 & 8'hfc; // @[NV_NVDLA_CSC_sg.scala 492:127:@1934.4]
  assign _T_779 = _T_778[6:0]; // @[NV_NVDLA_CSC_sg.scala 492:147:@1935.4]
  assign _T_781 = io_reg2dp_y_extension == 2'h1; // @[NV_NVDLA_CSC_sg.scala 493:61:@1936.4]
  assign _T_783 = _T_754 + 7'h1; // @[NV_NVDLA_CSC_sg.scala 493:106:@1937.4]
  assign _T_785 = _T_783 & 8'hfe; // @[NV_NVDLA_CSC_sg.scala 493:127:@1938.4]
  assign _T_786 = _T_785[6:0]; // @[NV_NVDLA_CSC_sg.scala 493:147:@1939.4]
  assign _T_787 = _T_781 ? _T_786 : _T_754; // @[NV_NVDLA_CSC_sg.scala 493:38:@1940.4]
  assign _T_788 = _T_774 ? _T_779 : _T_787; // @[NV_NVDLA_CSC_sg.scala 492:38:@1941.4]
  assign _T_789 = _T_472 ? 7'h0 : _T_788; // @[NV_NVDLA_CSC_sg.scala 491:38:@1942.4]
  assign _T_790 = _T_384 ? _T_789 : _T_754; // @[NV_NVDLA_CSC_sg.scala 496:34:@1943.4]
  assign _T_814 = ~ _T_867; // @[NV_NVDLA_CSC_sg.scala 508:30:@1952.4]
  assign _T_817 = _T_796 < 7'h20; // @[NV_NVDLA_CSC_sg.scala 509:49:@1953.4]
  assign _T_819 = _T_817 ? 7'h20 : _T_796; // @[NV_NVDLA_CSC_sg.scala 509:29:@1954.4]
  assign _T_820 = _T_814 ? 7'h0 : _T_819; // @[NV_NVDLA_CSC_sg.scala 508:29:@1955.4]
  assign _T_856 = _T_861 & _T_885; // @[NV_NVDLA_CSC_sg.scala 520:54:@1981.4]
  assign _T_857 = _T_747 == _T_749; // @[NV_NVDLA_CSC_sg.scala 520:85:@1982.4]
  assign _T_858 = _T_856 | _T_857; // @[NV_NVDLA_CSC_sg.scala 520:70:@1983.4]
  assign _T_859 = _T_160 & _T_858; // @[NV_NVDLA_CSC_sg.scala 520:32:@1984.4]
  assign _T_821 = ~ _T_859; // @[NV_NVDLA_CSC_sg.scala 513:29:@1956.4]
  assign _T_824 = _T_762 <= 6'h1; // @[NV_NVDLA_CSC_sg.scala 514:41:@1957.4]
  assign _T_826 = _T_799 <= 6'h1; // @[NV_NVDLA_CSC_sg.scala 514:73:@1958.4]
  assign _T_827 = _T_824 & _T_826; // @[NV_NVDLA_CSC_sg.scala 514:62:@1959.4]
  assign _T_829 = _T_762 > _T_799; // @[NV_NVDLA_CSC_sg.scala 515:41:@1960.4]
  assign _T_830 = _T_829 ? _T_762 : _T_799; // @[NV_NVDLA_CSC_sg.scala 515:29:@1961.4]
  assign _T_831 = _T_827 ? 6'h2 : _T_830; // @[NV_NVDLA_CSC_sg.scala 514:29:@1962.4]
  assign _T_832 = _T_821 ? 6'h0 : _T_831; // @[NV_NVDLA_CSC_sg.scala 513:28:@1963.4]
  assign _GEN_71 = {{1'd0}, _T_832}; // @[NV_NVDLA_CSC_sg.scala 517:41:@1964.4]
  assign _T_833 = _T_820 >= _GEN_71; // @[NV_NVDLA_CSC_sg.scala 517:41:@1964.4]
  assign _T_835 = _T_820 - 7'h1; // @[NV_NVDLA_CSC_sg.scala 517:76:@1965.4]
  assign _T_836 = $unsigned(_T_835); // @[NV_NVDLA_CSC_sg.scala 517:76:@1966.4]
  assign _T_837 = _T_836[6:0]; // @[NV_NVDLA_CSC_sg.scala 517:76:@1967.4]
  assign _T_839 = _T_832 - 6'h1; // @[NV_NVDLA_CSC_sg.scala 517:99:@1968.4]
  assign _T_840 = $unsigned(_T_839); // @[NV_NVDLA_CSC_sg.scala 517:99:@1969.4]
  assign _T_841 = _T_840[5:0]; // @[NV_NVDLA_CSC_sg.scala 517:99:@1970.4]
  assign _T_842 = _T_833 ? _T_837 : {{1'd0}, _T_841}; // @[NV_NVDLA_CSC_sg.scala 517:25:@1971.4]
  assign _T_843 = _T_842[5:0]; // @[NV_NVDLA_CSC_sg.scala 517:106:@1972.4]
  assign _T_845 = _T_799 - 6'h1; // @[NV_NVDLA_CSC_sg.scala 518:31:@1973.4]
  assign _T_846 = $unsigned(_T_845); // @[NV_NVDLA_CSC_sg.scala 518:31:@1974.4]
  assign _T_847 = _T_846[5:0]; // @[NV_NVDLA_CSC_sg.scala 518:31:@1975.4]
  assign _T_848 = _T_867 | _T_859; // @[NV_NVDLA_CSC_sg.scala 519:39:@1976.4]
  assign _T_852 = _T_861 ? 6'h0 : _T_847; // @[NV_NVDLA_CSC_sg.scala 519:70:@1978.4]
  assign _T_853 = _T_848 ? _T_843 : _T_852; // @[NV_NVDLA_CSC_sg.scala 519:24:@1979.4]
  assign _GEN_54 = _T_793 ? _T_754 : _T_191; // @[NV_NVDLA_CSC_sg.scala 525:26:@1995.4]
  assign _GEN_55 = _T_793 ? _T_790 : _T_796; // @[NV_NVDLA_CSC_sg.scala 525:26:@1995.4]
  assign _GEN_57 = _T_859 ? _T_750 : _T_811; // @[NV_NVDLA_CSC_sg.scala 535:23:@2005.4]
  assign _T_879 = _T_873 ? {{1'd0}, _T_875} : 4'h0; // @[NV_NVDLA_CSC_sg.scala 559:29:@2020.4]
  assign _T_880 = _T_867 & _T_757; // @[NV_NVDLA_CSC_sg.scala 560:43:@2021.4]
  assign _T_882 = _T_880 ? _T_877 : 9'h0; // @[NV_NVDLA_CSC_sg.scala 560:29:@2022.4]
  assign _T_886 = _T_867 | _T_873; // @[NV_NVDLA_CSC_sg.scala 563:24:@2027.4]
  assign _GEN_72 = {{5'd0}, _T_879}; // @[NV_NVDLA_CSC_sg.scala 564:34:@2029.6]
  assign _T_887 = _T_870 + _GEN_72; // @[NV_NVDLA_CSC_sg.scala 564:34:@2029.6]
  assign _T_888 = _T_870 + _GEN_72; // @[NV_NVDLA_CSC_sg.scala 564:34:@2030.6]
  assign _T_889 = _T_888 - _T_882; // @[NV_NVDLA_CSC_sg.scala 564:51:@2031.6]
  assign _T_890 = $unsigned(_T_889); // @[NV_NVDLA_CSC_sg.scala 564:51:@2032.6]
  assign _T_891 = _T_890[8:0]; // @[NV_NVDLA_CSC_sg.scala 564:51:@2033.6]
  assign _GEN_59 = _T_886 ? _T_891 : _T_870; // @[NV_NVDLA_CSC_sg.scala 563:37:@2028.4]
  assign _T_892 = _T_621 & _T_697; // @[NV_NVDLA_CSC_sg.scala 570:31:@2036.4]
  assign _T_894 = _T_892 & _T_704; // @[NV_NVDLA_CSC_sg.scala 570:49:@2038.4]
  assign _T_895 = _T_238 & io_reg2dp_op_en; // @[NV_NVDLA_CSC_sg.scala 571:37:@2039.4]
  assign _T_896 = ~ io_reg2dp_data_reuse; // @[NV_NVDLA_CSC_sg.scala 571:58:@2040.4]
  assign _T_897 = _T_896 | _T_253; // @[NV_NVDLA_CSC_sg.scala 571:80:@2041.4]
  assign _T_898 = _T_895 & _T_897; // @[NV_NVDLA_CSC_sg.scala 571:55:@2042.4]
  assign _T_900 = _T_289 != 14'h0; // @[NV_NVDLA_CSC_sg.scala 571:113:@2043.4]
  assign _T_901 = _T_898 & _T_900; // @[NV_NVDLA_CSC_sg.scala 571:98:@2044.4]
  assign _T_903 = io_cdma2sc_dat_updt_valid ? io_cdma2sc_dat_updt_bits_slices : 14'h0; // @[NV_NVDLA_CSC_sg.scala 572:29:@2045.4]
  assign _T_905 = _T_901 ? _T_289 : 14'h0; // @[NV_NVDLA_CSC_sg.scala 573:58:@2046.4]
  assign _T_906 = _T_894 ? _T_381 : _T_905; // @[NV_NVDLA_CSC_sg.scala 573:29:@2047.4]
  assign _T_908 = _T_621 & _T_606; // @[NV_NVDLA_CSC_sg.scala 574:30:@2049.4]
  assign _T_909 = _T_908 & _T_693; // @[NV_NVDLA_CSC_sg.scala 574:59:@2050.4]
  assign _T_911 = ~ io_reg2dp_weight_reuse; // @[NV_NVDLA_CSC_sg.scala 575:56:@2052.4]
  assign _T_912 = _T_895 & _T_911; // @[NV_NVDLA_CSC_sg.scala 575:54:@2053.4]
  assign _T_913 = _T_912 & _T_306; // @[NV_NVDLA_CSC_sg.scala 575:80:@2054.4]
  assign _T_915 = io_cdma2sc_wt_updt_valid ? io_cdma2sc_wt_updt_bits_kernels : 14'h0; // @[NV_NVDLA_CSC_sg.scala 576:30:@2055.4]
  assign _T_917 = {7'h0,_T_459}; // @[Cat.scala 30:58:@2056.4]
  assign _T_919 = _T_913 ? _T_303 : 14'h0; // @[NV_NVDLA_CSC_sg.scala 577:81:@2057.4]
  assign _T_920 = _T_909 ? {{1'd0}, _T_917} : _T_919; // @[NV_NVDLA_CSC_sg.scala 577:30:@2058.4]
  assign _T_921 = _T_174 | _T_894; // @[NV_NVDLA_CSC_sg.scala 579:26:@2059.4]
  assign _T_922 = _T_921 | _T_901; // @[NV_NVDLA_CSC_sg.scala 579:40:@2060.4]
  assign _T_923 = _T_922 | io_cdma2sc_dat_updt_valid; // @[NV_NVDLA_CSC_sg.scala 579:60:@2061.4]
  assign _T_925 = _T_593 + _T_903; // @[NV_NVDLA_CSC_sg.scala 580:75:@2063.6]
  assign _T_926 = _T_593 + _T_903; // @[NV_NVDLA_CSC_sg.scala 580:75:@2064.6]
  assign _T_927 = _T_926 - _T_906; // @[NV_NVDLA_CSC_sg.scala 580:92:@2065.6]
  assign _T_928 = $unsigned(_T_927); // @[NV_NVDLA_CSC_sg.scala 580:92:@2066.6]
  assign _T_929 = _T_928[13:0]; // @[NV_NVDLA_CSC_sg.scala 580:92:@2067.6]
  assign _T_930 = _T_174 ? 14'h0 : _T_929; // @[NV_NVDLA_CSC_sg.scala 580:26:@2068.6]
  assign _GEN_60 = _T_923 ? _T_930 : _T_593; // @[NV_NVDLA_CSC_sg.scala 579:88:@2062.4]
  assign _T_931 = _T_183 | _T_909; // @[NV_NVDLA_CSC_sg.scala 582:25:@2071.4]
  assign _T_932 = _T_931 | _T_913; // @[NV_NVDLA_CSC_sg.scala 582:38:@2072.4]
  assign _T_933 = _T_932 | io_cdma2sc_wt_updt_valid; // @[NV_NVDLA_CSC_sg.scala 582:57:@2073.4]
  assign _GEN_73 = {{1'd0}, _T_915}; // @[NV_NVDLA_CSC_sg.scala 583:75:@2075.6]
  assign _T_935 = _T_599 + _GEN_73; // @[NV_NVDLA_CSC_sg.scala 583:75:@2075.6]
  assign _T_936 = _T_599 + _GEN_73; // @[NV_NVDLA_CSC_sg.scala 583:75:@2076.6]
  assign _GEN_74 = {{1'd0}, _T_920}; // @[NV_NVDLA_CSC_sg.scala 583:93:@2077.6]
  assign _T_937 = _T_936 - _GEN_74; // @[NV_NVDLA_CSC_sg.scala 583:93:@2077.6]
  assign _T_938 = $unsigned(_T_937); // @[NV_NVDLA_CSC_sg.scala 583:93:@2078.6]
  assign _T_939 = _T_938[14:0]; // @[NV_NVDLA_CSC_sg.scala 583:93:@2079.6]
  assign _T_940 = _T_183 ? 15'h0 : _T_939; // @[NV_NVDLA_CSC_sg.scala 583:27:@2080.6]
  assign _GEN_61 = _T_933 ? _T_940 : _T_599; // @[NV_NVDLA_CSC_sg.scala 582:84:@2074.4]
  assign io_sc2cdma_dat_pending_req = _T_174; // @[NV_NVDLA_CSC_sg.scala 175:32:@1549.4]
  assign io_sc2cdma_wt_pending_req = _T_183; // @[NV_NVDLA_CSC_sg.scala 176:31:@1550.4]
  assign io_sc_state = _T_238 ? 2'h0 : _T_251; // @[NV_NVDLA_CSC_sg.scala 165:17:@1523.4]
  assign io_sg2dl_pd_valid = _T_802; // @[NV_NVDLA_CSC_sg.scala 539:23:@2008.4]
  assign io_sg2dl_reuse_rls = _T_943; // @[NV_NVDLA_CSC_sg.scala 586:24:@2085.4]
  assign io_sg2wl_pd_valid = _T_808; // @[NV_NVDLA_CSC_sg.scala 541:23:@2010.4]
  assign io_sg2wl_pd_bits = _T_811; // @[NV_NVDLA_CSC_sg.scala 542:22:@2011.4]
  assign io_sg2wl_reuse_rls = _T_946; // @[NV_NVDLA_CSC_sg.scala 587:24:@2088.4]
  assign io_dp2reg_done = _T_259; // @[NV_NVDLA_CSC_sg.scala 168:20:@1529.4]
  assign NV_NVDLA_fifo_clock = io_nvdla_core_clk; // @[:@1886.4]
  assign NV_NVDLA_fifo_reset = reset; // @[:@1887.4]
  assign NV_NVDLA_fifo_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CSC_sg.scala 436:23:@1888.4]
  assign NV_NVDLA_fifo_io_wr_pvld = _T_136 & _T_613; // @[NV_NVDLA_CSC_sg.scala 438:27:@1890.4]
  assign NV_NVDLA_fifo_io_wr_pd = {_T_654,_T_731}; // @[NV_NVDLA_CSC_sg.scala 440:25:@1892.4]
  assign NV_NVDLA_fifo_io_rd_prdy = _T_863 & _T_866; // @[NV_NVDLA_CSC_sg.scala 442:27:@1894.4]
  assign NV_NVDLA_fifo_1_clock = io_nvdla_core_clk; // @[:@1897.4]
  assign NV_NVDLA_fifo_1_reset = reset; // @[:@1898.4]
  assign NV_NVDLA_fifo_1_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CSC_sg.scala 449:22:@1899.4]
  assign NV_NVDLA_fifo_1_io_wr_pvld = _T_136 & _T_611; // @[NV_NVDLA_CSC_sg.scala 451:26:@1901.4]
  assign NV_NVDLA_fifo_1_io_wr_pd = {_T_654,_T_741}; // @[NV_NVDLA_CSC_sg.scala 453:24:@1903.4]
  assign NV_NVDLA_fifo_1_io_rd_prdy = _T_160 & _T_858; // @[NV_NVDLA_CSC_sg.scala 455:26:@1905.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_131 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_136 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_165 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_168 = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_171 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_174 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_180 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_183 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_177 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_186 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_191 = _RAND_11[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_198 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_201 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_799 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_870 = _RAND_15[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_237 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_259 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_289 = _RAND_18[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_296 = _RAND_19[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_303 = _RAND_20[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_306 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_326 = _RAND_22[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_333 = _RAND_23[21:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_347 = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_354 = _RAND_25[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_361 = _RAND_26[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_368 = _RAND_27[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_371 = _RAND_28[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_374 = _RAND_29[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_381 = _RAND_30[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_384 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_387 = _RAND_32[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_390 = _RAND_33[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_593 = _RAND_34[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_596 = _RAND_35[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_449 = _RAND_36[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_599 = _RAND_37[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_554 = _RAND_38[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_561 = _RAND_39[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_524 = _RAND_40[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_489 = _RAND_41[21:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_469 = _RAND_42[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_654 = _RAND_43[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_657 = _RAND_44[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_660 = _RAND_45[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_663 = _RAND_46[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_666 = _RAND_47[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_669 = _RAND_48[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_672 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_675 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_678 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_681 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_684 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_708 = _RAND_54[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_711 = _RAND_55[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_714 = _RAND_56[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_717 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_793 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_796 = _RAND_59[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_802 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_808 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_811 = _RAND_62[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_873 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_875 = _RAND_64[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_943 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_946 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_131 <= 1'h0;
    end else begin
      if (_T_436) begin
        if (_T_239) begin
          _T_131 <= 1'h0;
        end else begin
          if (_T_453) begin
            _T_131 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_136 <= 1'h0;
    end else begin
      if (_T_639) begin
        _T_136 <= 1'h0;
      end else begin
        if (_T_642) begin
          _T_136 <= 1'h1;
        end else begin
          if (_T_614) begin
            _T_136 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_142 <= 2'h0;
    end else begin
      if (_T_145) begin
        if (_T_146) begin
          _T_142 <= 2'h1;
        end else begin
          if (io_reg2dp_op_en) begin
            _T_142 <= 2'h2;
          end else begin
            _T_142 <= 2'h0;
          end
        end
      end else begin
        if (_T_147) begin
          if (_T_217) begin
            _T_142 <= 2'h2;
          end else begin
            _T_142 <= 2'h0;
          end
        end else begin
          if (_T_148) begin
            if (_T_151) begin
              _T_142 <= 2'h3;
            end else begin
              _T_142 <= 2'h0;
            end
          end else begin
            _T_142 <= 2'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_165 <= 5'h1f;
    end else begin
      if (io_dp2reg_done) begin
        _T_165 <= io_reg2dp_data_bank;
      end
    end
    if (reset) begin
      _T_168 <= 5'h1f;
    end else begin
      if (io_dp2reg_done) begin
        _T_168 <= io_reg2dp_weight_bank;
      end
    end
    if (reset) begin
      _T_171 <= 1'h0;
    end else begin
      if (_T_271) begin
        _T_171 <= 1'h1;
      end else begin
        if (_T_262) begin
          _T_171 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_174 <= 1'h0;
    end else begin
      if (_T_260) begin
        _T_174 <= 1'h1;
      end else begin
        if (_T_262) begin
          _T_174 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      if (_T_277) begin
        _T_180 <= 1'h1;
      end else begin
        if (_T_262) begin
          _T_180 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_183 <= 1'h0;
    end else begin
      if (_T_245) begin
        _T_183 <= 1'h1;
      end else begin
        if (_T_262) begin
          _T_183 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_177 <= 1'h0;
    end else begin
      _T_177 <= io_cdma2sc_dat_pending_ack;
    end
    if (reset) begin
      _T_186 <= 1'h0;
    end else begin
      _T_186 <= io_cdma2sc_wt_pending_ack;
    end
    if (reset) begin
      _T_191 <= 7'h0;
    end else begin
      if (_T_793) begin
        _T_191 <= _T_754;
      end
    end
    if (reset) begin
      _T_198 <= 8'h0;
    end else begin
      if (_T_226) begin
        _T_198 <= _T_228;
      end
    end
    if (reset) begin
      _T_201 <= 8'h0;
    end else begin
      if (_T_244) begin
        if (_T_219) begin
          _T_201 <= _T_198;
        end else begin
          _T_201 <= _T_223;
        end
      end
    end
    if (reset) begin
      _T_799 <= 6'h0;
    end else begin
      if (_T_848) begin
        _T_799 <= _T_843;
      end else begin
        if (_T_861) begin
          _T_799 <= 6'h0;
        end else begin
          _T_799 <= _T_847;
        end
      end
    end
    if (reset) begin
      _T_237 <= 3'h0;
    end else begin
      if (io_dp2reg_done) begin
        _T_237 <= _T_318;
      end
    end
    if (reset) begin
      _T_259 <= 1'h0;
    end else begin
      _T_259 <= _T_256;
    end
    if (reset) begin
      _T_289 <= 14'h0;
    end else begin
      if (io_dp2reg_done) begin
        _T_289 <= _T_296;
      end
    end
    if (reset) begin
      _T_296 <= 14'h0;
    end else begin
      if (_T_239) begin
        if (io_reg2dp_skip_data_rls) begin
          _T_296 <= _T_395;
        end else begin
          _T_296 <= _T_424;
        end
      end
    end
    if (reset) begin
      _T_303 <= 14'h0;
    end else begin
      if (io_dp2reg_done) begin
        _T_303 <= _T_308;
      end
    end
    if (reset) begin
      _T_306 <= 1'h0;
    end else begin
      if (io_dp2reg_done) begin
        _T_306 <= io_reg2dp_skip_weight_rls;
      end
    end
    if (reset) begin
      _T_326 <= 14'h0;
    end else begin
      if (_T_239) begin
        _T_326 <= _T_395;
      end
    end
    if (reset) begin
      _T_333 <= 22'h0;
    end else begin
      if (_T_239) begin
        if (_T_313) begin
          _T_333 <= {{8'd0}, _T_397};
        end else begin
          _T_333 <= _T_399;
        end
      end
    end
    if (reset) begin
      _T_347 <= 5'h0;
    end else begin
      if (_T_239) begin
        if (_T_313) begin
          _T_347 <= 5'h0;
        end else begin
          _T_347 <= io_reg2dp_weight_width_ext;
        end
      end
    end
    if (reset) begin
      _T_354 <= 5'h0;
    end else begin
      if (_T_239) begin
        _T_354 <= io_reg2dp_weight_height_ext;
      end
    end
    if (reset) begin
      _T_361 <= 14'h0;
    end else begin
      if (_T_239) begin
        _T_361 <= _T_405;
      end
    end
    if (reset) begin
      _T_368 <= 10'h0;
    end else begin
      if (_T_239) begin
        _T_368 <= {{1'd0}, _T_408};
      end
    end
    if (reset) begin
      _T_371 <= 3'h1;
    end else begin
      if (_T_239) begin
        _T_371 <= _T_393;
      end
    end
    if (reset) begin
      _T_374 <= 3'h1;
    end else begin
      if (_T_239) begin
        _T_374 <= {{1'd0}, _T_417};
      end
    end
    if (reset) begin
      _T_381 <= 14'h0;
    end else begin
      if (_T_239) begin
        _T_381 <= {{2'd0}, _T_420};
      end
    end
    if (reset) begin
      _T_384 <= 1'h0;
    end else begin
      if (_T_239) begin
        _T_384 <= _T_313;
      end
    end
    if (reset) begin
      _T_387 <= 6'h20;
    end else begin
      _T_387 <= _GEN_29[5:0];
    end
    if (reset) begin
      _T_390 <= 7'h40;
    end else begin
      if (_T_239) begin
        _T_390 <= 7'h40;
      end
    end
    if (reset) begin
      _T_593 <= 14'h0;
    end else begin
      if (_T_923) begin
        if (_T_174) begin
          _T_593 <= 14'h0;
        end else begin
          _T_593 <= _T_929;
        end
      end
    end
    if (reset) begin
      _T_596 <= 14'h0;
    end else begin
      if (_T_460) begin
        if (_T_607) begin
          _T_596 <= 14'h0;
        end else begin
          _T_596 <= _T_602;
        end
      end
    end
    if (reset) begin
      _T_449 <= 10'h0;
    end else begin
      if (_T_460) begin
        if (_T_239) begin
          _T_449 <= 10'h0;
        end else begin
          _T_449 <= _T_452;
        end
      end
    end
    if (reset) begin
      _T_599 <= 15'h0;
    end else begin
      if (_T_933) begin
        if (_T_183) begin
          _T_599 <= 15'h0;
        end else begin
          _T_599 <= _T_939;
        end
      end
    end
    if (reset) begin
      _T_554 <= 5'h0;
    end else begin
      if (_T_581) begin
        if (_T_239) begin
          _T_554 <= 5'h0;
        end else begin
          if (_T_570) begin
            _T_554 <= 5'h0;
          end else begin
            _T_554 <= _T_568;
          end
        end
      end
    end
    if (reset) begin
      _T_561 <= 5'h0;
    end else begin
      if (_T_581) begin
        if (_T_239) begin
          _T_561 <= 5'h0;
        end else begin
          if (_T_571) begin
            _T_561 <= 5'h0;
          end else begin
            _T_561 <= _T_588;
          end
        end
      end
    end
    if (reset) begin
      _T_524 <= 14'h0;
    end else begin
      if (_T_535) begin
        if (_T_239) begin
          _T_524 <= 14'h0;
        end else begin
          if (_T_528) begin
            _T_524 <= 14'h0;
          end else begin
            _T_524 <= _T_527;
          end
        end
      end
    end
    if (reset) begin
      _T_489 <= 22'h0;
    end else begin
      if (_T_506) begin
        if (_T_239) begin
          _T_489 <= 22'h0;
        end else begin
          if (_T_497) begin
            _T_489 <= 22'h0;
          end else begin
            if (_T_496) begin
              _T_489 <= _T_495;
            end else begin
              _T_489 <= _T_512;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_469 <= 13'h0;
    end else begin
      if (_T_475) begin
        if (_T_239) begin
          _T_469 <= 13'h0;
        end else begin
          if (_T_474) begin
            _T_469 <= 13'h0;
          end else begin
            _T_469 <= _T_480;
          end
        end
      end
    end
    if (reset) begin
      _T_654 <= 2'h3;
    end else begin
      if (_T_581) begin
        if (_T_239) begin
          _T_654 <= 2'h3;
        end else begin
          _T_654 <= _T_688;
        end
      end
    end
    if (reset) begin
      _T_657 <= 5'h0;
    end else begin
      if (_T_621) begin
        _T_657 <= _T_554;
      end
    end
    if (reset) begin
      _T_660 <= 5'h0;
    end else begin
      if (_T_621) begin
        _T_660 <= _T_561;
      end
    end
    if (reset) begin
      _T_663 <= 7'h0;
    end else begin
      if (_T_621) begin
        if (_T_529) begin
          _T_663 <= 7'h40;
        end else begin
          _T_663 <= _T_533;
        end
      end
    end
    if (reset) begin
      _T_666 <= 7'h0;
    end else begin
      if (_T_621) begin
        if (_T_496) begin
          _T_666 <= _T_390;
        end else begin
          if (_T_497) begin
            _T_666 <= _T_501;
          end else begin
            _T_666 <= {{1'd0}, _T_387};
          end
        end
      end
    end
    if (reset) begin
      _T_669 <= 3'h0;
    end else begin
      if (_T_621) begin
        if (_T_571) begin
          _T_669 <= _T_374;
        end else begin
          _T_669 <= {{1'd0}, _T_578};
        end
      end
    end
    if (reset) begin
      _T_672 <= 1'h0;
    end else begin
      if (_T_621) begin
        _T_672 <= _T_580;
      end
    end
    if (reset) begin
      _T_675 <= 1'h0;
    end else begin
      if (_T_621) begin
        _T_675 <= _T_690;
      end
    end
    if (reset) begin
      _T_678 <= 1'h0;
    end else begin
      if (_T_621) begin
        _T_678 <= _T_693;
      end
    end
    if (reset) begin
      _T_681 <= 1'h0;
    end else begin
      if (_T_621) begin
        _T_681 <= _T_697;
      end
    end
    if (reset) begin
      _T_684 <= 1'h0;
    end else begin
      if (_T_621) begin
        _T_684 <= _T_705;
      end
    end
    if (reset) begin
      _T_708 <= 7'h0;
    end else begin
      if (_T_621) begin
        _T_708 <= {{1'd0}, _T_459};
      end
    end
    if (reset) begin
      _T_711 <= 7'h0;
    end else begin
      if (_T_621) begin
        if (_T_529) begin
          _T_711 <= 7'h40;
        end else begin
          _T_711 <= _T_533;
        end
      end
    end
    if (reset) begin
      _T_714 <= 3'h0;
    end else begin
      if (_T_621) begin
        if (_T_571) begin
          _T_714 <= _T_374;
        end else begin
          _T_714 <= {{1'd0}, _T_578};
        end
      end
    end
    if (reset) begin
      _T_717 <= 1'h0;
    end else begin
      if (_T_621) begin
        _T_717 <= _T_734;
      end
    end
    if (reset) begin
      _T_793 <= 1'h0;
    end else begin
      _T_793 <= _T_859;
    end
    if (reset) begin
      _T_796 <= 7'h0;
    end else begin
      if (_T_793) begin
        if (_T_384) begin
          if (_T_472) begin
            _T_796 <= 7'h0;
          end else begin
            if (_T_774) begin
              _T_796 <= _T_779;
            end else begin
              if (_T_781) begin
                _T_796 <= _T_786;
              end else begin
                _T_796 <= _T_754;
              end
            end
          end
        end else begin
          _T_796 <= _T_754;
        end
      end
    end
    if (reset) begin
      _T_802 <= 1'h0;
    end else begin
      _T_802 <= _T_867;
    end
    if (reset) begin
      _T_808 <= 1'h0;
    end else begin
      _T_808 <= _T_859;
    end
    if (reset) begin
      _T_811 <= 18'h0;
    end else begin
      if (_T_859) begin
        _T_811 <= _T_750;
      end
    end
  end
  always @(posedge io_nvdla_core_ng_clk) begin
    if (reset) begin
      _T_870 <= 9'h40;
    end else begin
      if (_T_886) begin
        _T_870 <= _T_891;
      end
    end
    if (reset) begin
      _T_873 <= 1'h0;
    end else begin
      _T_873 <= io_accu2sc_credit_size_valid;
    end
    if (io_accu2sc_credit_size_valid) begin
      _T_875 <= io_accu2sc_credit_size_bits;
    end
    if (reset) begin
      _T_943 <= 1'h0;
    end else begin
      _T_943 <= _T_901;
    end
    if (reset) begin
      _T_946 <= 1'h0;
    end else begin
      _T_946 <= _T_913;
    end
  end
endmodule
module NV_NVDLA_CSC_WL_dec( // @[:@2090.2]
  input        reset, // @[:@2092.4]
  input        io_nvdla_core_clk, // @[:@2093.4]
  input        io_input_valid, // @[:@2093.4]
  input        io_input_bits_mask_0, // @[:@2093.4]
  input        io_input_bits_mask_1, // @[:@2093.4]
  input        io_input_bits_mask_2, // @[:@2093.4]
  input        io_input_bits_mask_3, // @[:@2093.4]
  input        io_input_bits_mask_4, // @[:@2093.4]
  input        io_input_bits_mask_5, // @[:@2093.4]
  input        io_input_bits_mask_6, // @[:@2093.4]
  input        io_input_bits_mask_7, // @[:@2093.4]
  input        io_input_bits_mask_8, // @[:@2093.4]
  input        io_input_bits_mask_9, // @[:@2093.4]
  input        io_input_bits_mask_10, // @[:@2093.4]
  input        io_input_bits_mask_11, // @[:@2093.4]
  input        io_input_bits_mask_12, // @[:@2093.4]
  input        io_input_bits_mask_13, // @[:@2093.4]
  input        io_input_bits_mask_14, // @[:@2093.4]
  input        io_input_bits_mask_15, // @[:@2093.4]
  input        io_input_bits_mask_16, // @[:@2093.4]
  input        io_input_bits_mask_17, // @[:@2093.4]
  input        io_input_bits_mask_18, // @[:@2093.4]
  input        io_input_bits_mask_19, // @[:@2093.4]
  input        io_input_bits_mask_20, // @[:@2093.4]
  input        io_input_bits_mask_21, // @[:@2093.4]
  input        io_input_bits_mask_22, // @[:@2093.4]
  input        io_input_bits_mask_23, // @[:@2093.4]
  input        io_input_bits_mask_24, // @[:@2093.4]
  input        io_input_bits_mask_25, // @[:@2093.4]
  input        io_input_bits_mask_26, // @[:@2093.4]
  input        io_input_bits_mask_27, // @[:@2093.4]
  input        io_input_bits_mask_28, // @[:@2093.4]
  input        io_input_bits_mask_29, // @[:@2093.4]
  input        io_input_bits_mask_30, // @[:@2093.4]
  input        io_input_bits_mask_31, // @[:@2093.4]
  input        io_input_bits_mask_32, // @[:@2093.4]
  input        io_input_bits_mask_33, // @[:@2093.4]
  input        io_input_bits_mask_34, // @[:@2093.4]
  input        io_input_bits_mask_35, // @[:@2093.4]
  input        io_input_bits_mask_36, // @[:@2093.4]
  input        io_input_bits_mask_37, // @[:@2093.4]
  input        io_input_bits_mask_38, // @[:@2093.4]
  input        io_input_bits_mask_39, // @[:@2093.4]
  input        io_input_bits_mask_40, // @[:@2093.4]
  input        io_input_bits_mask_41, // @[:@2093.4]
  input        io_input_bits_mask_42, // @[:@2093.4]
  input        io_input_bits_mask_43, // @[:@2093.4]
  input        io_input_bits_mask_44, // @[:@2093.4]
  input        io_input_bits_mask_45, // @[:@2093.4]
  input        io_input_bits_mask_46, // @[:@2093.4]
  input        io_input_bits_mask_47, // @[:@2093.4]
  input        io_input_bits_mask_48, // @[:@2093.4]
  input        io_input_bits_mask_49, // @[:@2093.4]
  input        io_input_bits_mask_50, // @[:@2093.4]
  input        io_input_bits_mask_51, // @[:@2093.4]
  input        io_input_bits_mask_52, // @[:@2093.4]
  input        io_input_bits_mask_53, // @[:@2093.4]
  input        io_input_bits_mask_54, // @[:@2093.4]
  input        io_input_bits_mask_55, // @[:@2093.4]
  input        io_input_bits_mask_56, // @[:@2093.4]
  input        io_input_bits_mask_57, // @[:@2093.4]
  input        io_input_bits_mask_58, // @[:@2093.4]
  input        io_input_bits_mask_59, // @[:@2093.4]
  input        io_input_bits_mask_60, // @[:@2093.4]
  input        io_input_bits_mask_61, // @[:@2093.4]
  input        io_input_bits_mask_62, // @[:@2093.4]
  input        io_input_bits_mask_63, // @[:@2093.4]
  input  [7:0] io_input_bits_data_0, // @[:@2093.4]
  input  [7:0] io_input_bits_data_1, // @[:@2093.4]
  input  [7:0] io_input_bits_data_2, // @[:@2093.4]
  input  [7:0] io_input_bits_data_3, // @[:@2093.4]
  input  [7:0] io_input_bits_data_4, // @[:@2093.4]
  input  [7:0] io_input_bits_data_5, // @[:@2093.4]
  input  [7:0] io_input_bits_data_6, // @[:@2093.4]
  input  [7:0] io_input_bits_data_7, // @[:@2093.4]
  input  [7:0] io_input_bits_data_8, // @[:@2093.4]
  input  [7:0] io_input_bits_data_9, // @[:@2093.4]
  input  [7:0] io_input_bits_data_10, // @[:@2093.4]
  input  [7:0] io_input_bits_data_11, // @[:@2093.4]
  input  [7:0] io_input_bits_data_12, // @[:@2093.4]
  input  [7:0] io_input_bits_data_13, // @[:@2093.4]
  input  [7:0] io_input_bits_data_14, // @[:@2093.4]
  input  [7:0] io_input_bits_data_15, // @[:@2093.4]
  input  [7:0] io_input_bits_data_16, // @[:@2093.4]
  input  [7:0] io_input_bits_data_17, // @[:@2093.4]
  input  [7:0] io_input_bits_data_18, // @[:@2093.4]
  input  [7:0] io_input_bits_data_19, // @[:@2093.4]
  input  [7:0] io_input_bits_data_20, // @[:@2093.4]
  input  [7:0] io_input_bits_data_21, // @[:@2093.4]
  input  [7:0] io_input_bits_data_22, // @[:@2093.4]
  input  [7:0] io_input_bits_data_23, // @[:@2093.4]
  input  [7:0] io_input_bits_data_24, // @[:@2093.4]
  input  [7:0] io_input_bits_data_25, // @[:@2093.4]
  input  [7:0] io_input_bits_data_26, // @[:@2093.4]
  input  [7:0] io_input_bits_data_27, // @[:@2093.4]
  input  [7:0] io_input_bits_data_28, // @[:@2093.4]
  input  [7:0] io_input_bits_data_29, // @[:@2093.4]
  input  [7:0] io_input_bits_data_30, // @[:@2093.4]
  input  [7:0] io_input_bits_data_31, // @[:@2093.4]
  input  [7:0] io_input_bits_data_32, // @[:@2093.4]
  input  [7:0] io_input_bits_data_33, // @[:@2093.4]
  input  [7:0] io_input_bits_data_34, // @[:@2093.4]
  input  [7:0] io_input_bits_data_35, // @[:@2093.4]
  input  [7:0] io_input_bits_data_36, // @[:@2093.4]
  input  [7:0] io_input_bits_data_37, // @[:@2093.4]
  input  [7:0] io_input_bits_data_38, // @[:@2093.4]
  input  [7:0] io_input_bits_data_39, // @[:@2093.4]
  input  [7:0] io_input_bits_data_40, // @[:@2093.4]
  input  [7:0] io_input_bits_data_41, // @[:@2093.4]
  input  [7:0] io_input_bits_data_42, // @[:@2093.4]
  input  [7:0] io_input_bits_data_43, // @[:@2093.4]
  input  [7:0] io_input_bits_data_44, // @[:@2093.4]
  input  [7:0] io_input_bits_data_45, // @[:@2093.4]
  input  [7:0] io_input_bits_data_46, // @[:@2093.4]
  input  [7:0] io_input_bits_data_47, // @[:@2093.4]
  input  [7:0] io_input_bits_data_48, // @[:@2093.4]
  input  [7:0] io_input_bits_data_49, // @[:@2093.4]
  input  [7:0] io_input_bits_data_50, // @[:@2093.4]
  input  [7:0] io_input_bits_data_51, // @[:@2093.4]
  input  [7:0] io_input_bits_data_52, // @[:@2093.4]
  input  [7:0] io_input_bits_data_53, // @[:@2093.4]
  input  [7:0] io_input_bits_data_54, // @[:@2093.4]
  input  [7:0] io_input_bits_data_55, // @[:@2093.4]
  input  [7:0] io_input_bits_data_56, // @[:@2093.4]
  input  [7:0] io_input_bits_data_57, // @[:@2093.4]
  input  [7:0] io_input_bits_data_58, // @[:@2093.4]
  input  [7:0] io_input_bits_data_59, // @[:@2093.4]
  input  [7:0] io_input_bits_data_60, // @[:@2093.4]
  input  [7:0] io_input_bits_data_61, // @[:@2093.4]
  input  [7:0] io_input_bits_data_62, // @[:@2093.4]
  input  [7:0] io_input_bits_data_63, // @[:@2093.4]
  input        io_input_bits_sel_0, // @[:@2093.4]
  input        io_input_bits_sel_1, // @[:@2093.4]
  input        io_input_bits_sel_2, // @[:@2093.4]
  input        io_input_bits_sel_3, // @[:@2093.4]
  input        io_input_bits_sel_4, // @[:@2093.4]
  input        io_input_bits_sel_5, // @[:@2093.4]
  input        io_input_bits_sel_6, // @[:@2093.4]
  input        io_input_bits_sel_7, // @[:@2093.4]
  input        io_input_bits_sel_8, // @[:@2093.4]
  input        io_input_bits_sel_9, // @[:@2093.4]
  input        io_input_bits_sel_10, // @[:@2093.4]
  input        io_input_bits_sel_11, // @[:@2093.4]
  input        io_input_bits_sel_12, // @[:@2093.4]
  input        io_input_bits_sel_13, // @[:@2093.4]
  input        io_input_bits_sel_14, // @[:@2093.4]
  input        io_input_bits_sel_15, // @[:@2093.4]
  input        io_input_bits_sel_16, // @[:@2093.4]
  input        io_input_bits_sel_17, // @[:@2093.4]
  input        io_input_bits_sel_18, // @[:@2093.4]
  input        io_input_bits_sel_19, // @[:@2093.4]
  input        io_input_bits_sel_20, // @[:@2093.4]
  input        io_input_bits_sel_21, // @[:@2093.4]
  input        io_input_bits_sel_22, // @[:@2093.4]
  input        io_input_bits_sel_23, // @[:@2093.4]
  input        io_input_bits_sel_24, // @[:@2093.4]
  input        io_input_bits_sel_25, // @[:@2093.4]
  input        io_input_bits_sel_26, // @[:@2093.4]
  input        io_input_bits_sel_27, // @[:@2093.4]
  input        io_input_bits_sel_28, // @[:@2093.4]
  input        io_input_bits_sel_29, // @[:@2093.4]
  input        io_input_bits_sel_30, // @[:@2093.4]
  input        io_input_bits_sel_31, // @[:@2093.4]
  input  [9:0] io_input_mask_en, // @[:@2093.4]
  output       io_output_valid, // @[:@2093.4]
  output       io_output_bits_mask_0, // @[:@2093.4]
  output       io_output_bits_mask_1, // @[:@2093.4]
  output       io_output_bits_mask_2, // @[:@2093.4]
  output       io_output_bits_mask_3, // @[:@2093.4]
  output       io_output_bits_mask_4, // @[:@2093.4]
  output       io_output_bits_mask_5, // @[:@2093.4]
  output       io_output_bits_mask_6, // @[:@2093.4]
  output       io_output_bits_mask_7, // @[:@2093.4]
  output       io_output_bits_mask_8, // @[:@2093.4]
  output       io_output_bits_mask_9, // @[:@2093.4]
  output       io_output_bits_mask_10, // @[:@2093.4]
  output       io_output_bits_mask_11, // @[:@2093.4]
  output       io_output_bits_mask_12, // @[:@2093.4]
  output       io_output_bits_mask_13, // @[:@2093.4]
  output       io_output_bits_mask_14, // @[:@2093.4]
  output       io_output_bits_mask_15, // @[:@2093.4]
  output       io_output_bits_mask_16, // @[:@2093.4]
  output       io_output_bits_mask_17, // @[:@2093.4]
  output       io_output_bits_mask_18, // @[:@2093.4]
  output       io_output_bits_mask_19, // @[:@2093.4]
  output       io_output_bits_mask_20, // @[:@2093.4]
  output       io_output_bits_mask_21, // @[:@2093.4]
  output       io_output_bits_mask_22, // @[:@2093.4]
  output       io_output_bits_mask_23, // @[:@2093.4]
  output       io_output_bits_mask_24, // @[:@2093.4]
  output       io_output_bits_mask_25, // @[:@2093.4]
  output       io_output_bits_mask_26, // @[:@2093.4]
  output       io_output_bits_mask_27, // @[:@2093.4]
  output       io_output_bits_mask_28, // @[:@2093.4]
  output       io_output_bits_mask_29, // @[:@2093.4]
  output       io_output_bits_mask_30, // @[:@2093.4]
  output       io_output_bits_mask_31, // @[:@2093.4]
  output       io_output_bits_mask_32, // @[:@2093.4]
  output       io_output_bits_mask_33, // @[:@2093.4]
  output       io_output_bits_mask_34, // @[:@2093.4]
  output       io_output_bits_mask_35, // @[:@2093.4]
  output       io_output_bits_mask_36, // @[:@2093.4]
  output       io_output_bits_mask_37, // @[:@2093.4]
  output       io_output_bits_mask_38, // @[:@2093.4]
  output       io_output_bits_mask_39, // @[:@2093.4]
  output       io_output_bits_mask_40, // @[:@2093.4]
  output       io_output_bits_mask_41, // @[:@2093.4]
  output       io_output_bits_mask_42, // @[:@2093.4]
  output       io_output_bits_mask_43, // @[:@2093.4]
  output       io_output_bits_mask_44, // @[:@2093.4]
  output       io_output_bits_mask_45, // @[:@2093.4]
  output       io_output_bits_mask_46, // @[:@2093.4]
  output       io_output_bits_mask_47, // @[:@2093.4]
  output       io_output_bits_mask_48, // @[:@2093.4]
  output       io_output_bits_mask_49, // @[:@2093.4]
  output       io_output_bits_mask_50, // @[:@2093.4]
  output       io_output_bits_mask_51, // @[:@2093.4]
  output       io_output_bits_mask_52, // @[:@2093.4]
  output       io_output_bits_mask_53, // @[:@2093.4]
  output       io_output_bits_mask_54, // @[:@2093.4]
  output       io_output_bits_mask_55, // @[:@2093.4]
  output       io_output_bits_mask_56, // @[:@2093.4]
  output       io_output_bits_mask_57, // @[:@2093.4]
  output       io_output_bits_mask_58, // @[:@2093.4]
  output       io_output_bits_mask_59, // @[:@2093.4]
  output       io_output_bits_mask_60, // @[:@2093.4]
  output       io_output_bits_mask_61, // @[:@2093.4]
  output       io_output_bits_mask_62, // @[:@2093.4]
  output       io_output_bits_mask_63, // @[:@2093.4]
  output [7:0] io_output_bits_data_0, // @[:@2093.4]
  output [7:0] io_output_bits_data_1, // @[:@2093.4]
  output [7:0] io_output_bits_data_2, // @[:@2093.4]
  output [7:0] io_output_bits_data_3, // @[:@2093.4]
  output [7:0] io_output_bits_data_4, // @[:@2093.4]
  output [7:0] io_output_bits_data_5, // @[:@2093.4]
  output [7:0] io_output_bits_data_6, // @[:@2093.4]
  output [7:0] io_output_bits_data_7, // @[:@2093.4]
  output [7:0] io_output_bits_data_8, // @[:@2093.4]
  output [7:0] io_output_bits_data_9, // @[:@2093.4]
  output [7:0] io_output_bits_data_10, // @[:@2093.4]
  output [7:0] io_output_bits_data_11, // @[:@2093.4]
  output [7:0] io_output_bits_data_12, // @[:@2093.4]
  output [7:0] io_output_bits_data_13, // @[:@2093.4]
  output [7:0] io_output_bits_data_14, // @[:@2093.4]
  output [7:0] io_output_bits_data_15, // @[:@2093.4]
  output [7:0] io_output_bits_data_16, // @[:@2093.4]
  output [7:0] io_output_bits_data_17, // @[:@2093.4]
  output [7:0] io_output_bits_data_18, // @[:@2093.4]
  output [7:0] io_output_bits_data_19, // @[:@2093.4]
  output [7:0] io_output_bits_data_20, // @[:@2093.4]
  output [7:0] io_output_bits_data_21, // @[:@2093.4]
  output [7:0] io_output_bits_data_22, // @[:@2093.4]
  output [7:0] io_output_bits_data_23, // @[:@2093.4]
  output [7:0] io_output_bits_data_24, // @[:@2093.4]
  output [7:0] io_output_bits_data_25, // @[:@2093.4]
  output [7:0] io_output_bits_data_26, // @[:@2093.4]
  output [7:0] io_output_bits_data_27, // @[:@2093.4]
  output [7:0] io_output_bits_data_28, // @[:@2093.4]
  output [7:0] io_output_bits_data_29, // @[:@2093.4]
  output [7:0] io_output_bits_data_30, // @[:@2093.4]
  output [7:0] io_output_bits_data_31, // @[:@2093.4]
  output [7:0] io_output_bits_data_32, // @[:@2093.4]
  output [7:0] io_output_bits_data_33, // @[:@2093.4]
  output [7:0] io_output_bits_data_34, // @[:@2093.4]
  output [7:0] io_output_bits_data_35, // @[:@2093.4]
  output [7:0] io_output_bits_data_36, // @[:@2093.4]
  output [7:0] io_output_bits_data_37, // @[:@2093.4]
  output [7:0] io_output_bits_data_38, // @[:@2093.4]
  output [7:0] io_output_bits_data_39, // @[:@2093.4]
  output [7:0] io_output_bits_data_40, // @[:@2093.4]
  output [7:0] io_output_bits_data_41, // @[:@2093.4]
  output [7:0] io_output_bits_data_42, // @[:@2093.4]
  output [7:0] io_output_bits_data_43, // @[:@2093.4]
  output [7:0] io_output_bits_data_44, // @[:@2093.4]
  output [7:0] io_output_bits_data_45, // @[:@2093.4]
  output [7:0] io_output_bits_data_46, // @[:@2093.4]
  output [7:0] io_output_bits_data_47, // @[:@2093.4]
  output [7:0] io_output_bits_data_48, // @[:@2093.4]
  output [7:0] io_output_bits_data_49, // @[:@2093.4]
  output [7:0] io_output_bits_data_50, // @[:@2093.4]
  output [7:0] io_output_bits_data_51, // @[:@2093.4]
  output [7:0] io_output_bits_data_52, // @[:@2093.4]
  output [7:0] io_output_bits_data_53, // @[:@2093.4]
  output [7:0] io_output_bits_data_54, // @[:@2093.4]
  output [7:0] io_output_bits_data_55, // @[:@2093.4]
  output [7:0] io_output_bits_data_56, // @[:@2093.4]
  output [7:0] io_output_bits_data_57, // @[:@2093.4]
  output [7:0] io_output_bits_data_58, // @[:@2093.4]
  output [7:0] io_output_bits_data_59, // @[:@2093.4]
  output [7:0] io_output_bits_data_60, // @[:@2093.4]
  output [7:0] io_output_bits_data_61, // @[:@2093.4]
  output [7:0] io_output_bits_data_62, // @[:@2093.4]
  output [7:0] io_output_bits_data_63, // @[:@2093.4]
  output       io_output_bits_sel_0, // @[:@2093.4]
  output       io_output_bits_sel_1, // @[:@2093.4]
  output       io_output_bits_sel_2, // @[:@2093.4]
  output       io_output_bits_sel_3, // @[:@2093.4]
  output       io_output_bits_sel_4, // @[:@2093.4]
  output       io_output_bits_sel_5, // @[:@2093.4]
  output       io_output_bits_sel_6, // @[:@2093.4]
  output       io_output_bits_sel_7, // @[:@2093.4]
  output       io_output_bits_sel_8, // @[:@2093.4]
  output       io_output_bits_sel_9, // @[:@2093.4]
  output       io_output_bits_sel_10, // @[:@2093.4]
  output       io_output_bits_sel_11, // @[:@2093.4]
  output       io_output_bits_sel_12, // @[:@2093.4]
  output       io_output_bits_sel_13, // @[:@2093.4]
  output       io_output_bits_sel_14, // @[:@2093.4]
  output       io_output_bits_sel_15, // @[:@2093.4]
  output       io_output_bits_sel_16, // @[:@2093.4]
  output       io_output_bits_sel_17, // @[:@2093.4]
  output       io_output_bits_sel_18, // @[:@2093.4]
  output       io_output_bits_sel_19, // @[:@2093.4]
  output       io_output_bits_sel_20, // @[:@2093.4]
  output       io_output_bits_sel_21, // @[:@2093.4]
  output       io_output_bits_sel_22, // @[:@2093.4]
  output       io_output_bits_sel_23, // @[:@2093.4]
  output       io_output_bits_sel_24, // @[:@2093.4]
  output       io_output_bits_sel_25, // @[:@2093.4]
  output       io_output_bits_sel_26, // @[:@2093.4]
  output       io_output_bits_sel_27, // @[:@2093.4]
  output       io_output_bits_sel_28, // @[:@2093.4]
  output       io_output_bits_sel_29, // @[:@2093.4]
  output       io_output_bits_sel_30, // @[:@2093.4]
  output       io_output_bits_sel_31 // @[:@2093.4]
);
  wire  _T_1771; // @[NV_NVDLA_CSC_WL_dec.scala 56:48:@2095.4]
  wire  _T_1906_0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_1; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_2; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_3; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_4; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_5; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_6; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_7; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_8; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_9; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_10; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_11; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_12; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_13; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_14; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_15; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_16; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_17; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_18; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_19; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_20; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_21; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_22; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_23; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_24; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_25; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_26; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_27; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_28; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_29; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_30; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_31; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_32; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_33; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_34; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_35; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_36; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_37; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_38; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_39; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_40; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_41; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_42; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_43; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_44; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_45; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_46; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_47; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_48; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_49; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_50; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_51; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_52; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_53; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_54; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_55; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_56; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_57; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_58; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_59; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_60; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_61; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_62; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire  _T_1906_63; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  wire [7:0] _T_2174; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2169.4]
  wire [15:0] _T_2182; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2177.4]
  wire [7:0] _T_2189; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2184.4]
  wire [31:0] _T_2198; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2193.4]
  wire [7:0] _T_2205; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2200.4]
  wire [15:0] _T_2213; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2208.4]
  wire [7:0] _T_2220; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2215.4]
  wire [31:0] _T_2229; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2224.4]
  wire [63:0] _T_2230; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2225.4]
  wire  _T_2231; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2226.4]
  wire [1:0] _T_2296; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2292.4]
  wire  _T_2297; // @[Bitwise.scala 50:65:@2293.4]
  wire  _T_2298; // @[Bitwise.scala 50:65:@2294.4]
  wire [1:0] _T_2299; // @[Bitwise.scala 48:55:@2295.4]
  wire [2:0] _T_2363; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2360.4]
  wire  _T_2364; // @[Bitwise.scala 50:65:@2361.4]
  wire  _T_2365; // @[Bitwise.scala 50:65:@2362.4]
  wire  _T_2366; // @[Bitwise.scala 50:65:@2363.4]
  wire [1:0] _T_2367; // @[Bitwise.scala 48:55:@2364.4]
  wire [1:0] _GEN_544; // @[Bitwise.scala 48:55:@2365.4]
  wire [2:0] _T_2368; // @[Bitwise.scala 48:55:@2365.4]
  wire [3:0] _T_2432; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2430.4]
  wire  _T_2433; // @[Bitwise.scala 50:65:@2431.4]
  wire  _T_2434; // @[Bitwise.scala 50:65:@2432.4]
  wire  _T_2435; // @[Bitwise.scala 50:65:@2433.4]
  wire  _T_2436; // @[Bitwise.scala 50:65:@2434.4]
  wire [1:0] _T_2437; // @[Bitwise.scala 48:55:@2435.4]
  wire [1:0] _T_2438; // @[Bitwise.scala 48:55:@2436.4]
  wire [2:0] _T_2439; // @[Bitwise.scala 48:55:@2437.4]
  wire [4:0] _T_2503; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2502.4]
  wire  _T_2504; // @[Bitwise.scala 50:65:@2503.4]
  wire  _T_2505; // @[Bitwise.scala 50:65:@2504.4]
  wire  _T_2506; // @[Bitwise.scala 50:65:@2505.4]
  wire  _T_2507; // @[Bitwise.scala 50:65:@2506.4]
  wire  _T_2508; // @[Bitwise.scala 50:65:@2507.4]
  wire [1:0] _T_2509; // @[Bitwise.scala 48:55:@2508.4]
  wire [1:0] _T_2510; // @[Bitwise.scala 48:55:@2509.4]
  wire [1:0] _GEN_545; // @[Bitwise.scala 48:55:@2510.4]
  wire [2:0] _T_2511; // @[Bitwise.scala 48:55:@2510.4]
  wire [2:0] _GEN_546; // @[Bitwise.scala 48:55:@2511.4]
  wire [3:0] _T_2512; // @[Bitwise.scala 48:55:@2511.4]
  wire [5:0] _T_2576; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2576.4]
  wire  _T_2577; // @[Bitwise.scala 50:65:@2577.4]
  wire  _T_2578; // @[Bitwise.scala 50:65:@2578.4]
  wire  _T_2579; // @[Bitwise.scala 50:65:@2579.4]
  wire  _T_2580; // @[Bitwise.scala 50:65:@2580.4]
  wire  _T_2581; // @[Bitwise.scala 50:65:@2581.4]
  wire  _T_2582; // @[Bitwise.scala 50:65:@2582.4]
  wire [1:0] _T_2583; // @[Bitwise.scala 48:55:@2583.4]
  wire [1:0] _GEN_547; // @[Bitwise.scala 48:55:@2584.4]
  wire [2:0] _T_2584; // @[Bitwise.scala 48:55:@2584.4]
  wire [1:0] _T_2585; // @[Bitwise.scala 48:55:@2585.4]
  wire [1:0] _GEN_548; // @[Bitwise.scala 48:55:@2586.4]
  wire [2:0] _T_2586; // @[Bitwise.scala 48:55:@2586.4]
  wire [3:0] _T_2587; // @[Bitwise.scala 48:55:@2587.4]
  wire [6:0] _T_2651; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2652.4]
  wire  _T_2652; // @[Bitwise.scala 50:65:@2653.4]
  wire  _T_2653; // @[Bitwise.scala 50:65:@2654.4]
  wire  _T_2654; // @[Bitwise.scala 50:65:@2655.4]
  wire  _T_2655; // @[Bitwise.scala 50:65:@2656.4]
  wire  _T_2656; // @[Bitwise.scala 50:65:@2657.4]
  wire  _T_2657; // @[Bitwise.scala 50:65:@2658.4]
  wire  _T_2658; // @[Bitwise.scala 50:65:@2659.4]
  wire [1:0] _T_2659; // @[Bitwise.scala 48:55:@2660.4]
  wire [1:0] _GEN_549; // @[Bitwise.scala 48:55:@2661.4]
  wire [2:0] _T_2660; // @[Bitwise.scala 48:55:@2661.4]
  wire [1:0] _T_2661; // @[Bitwise.scala 48:55:@2662.4]
  wire [1:0] _T_2662; // @[Bitwise.scala 48:55:@2663.4]
  wire [2:0] _T_2663; // @[Bitwise.scala 48:55:@2664.4]
  wire [3:0] _T_2664; // @[Bitwise.scala 48:55:@2665.4]
  wire [7:0] _T_2728; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2730.4]
  wire  _T_2729; // @[Bitwise.scala 50:65:@2731.4]
  wire  _T_2730; // @[Bitwise.scala 50:65:@2732.4]
  wire  _T_2731; // @[Bitwise.scala 50:65:@2733.4]
  wire  _T_2732; // @[Bitwise.scala 50:65:@2734.4]
  wire  _T_2733; // @[Bitwise.scala 50:65:@2735.4]
  wire  _T_2734; // @[Bitwise.scala 50:65:@2736.4]
  wire  _T_2735; // @[Bitwise.scala 50:65:@2737.4]
  wire  _T_2736; // @[Bitwise.scala 50:65:@2738.4]
  wire [1:0] _T_2737; // @[Bitwise.scala 48:55:@2739.4]
  wire [1:0] _T_2738; // @[Bitwise.scala 48:55:@2740.4]
  wire [2:0] _T_2739; // @[Bitwise.scala 48:55:@2741.4]
  wire [1:0] _T_2740; // @[Bitwise.scala 48:55:@2742.4]
  wire [1:0] _T_2741; // @[Bitwise.scala 48:55:@2743.4]
  wire [2:0] _T_2742; // @[Bitwise.scala 48:55:@2744.4]
  wire [3:0] _T_2743; // @[Bitwise.scala 48:55:@2745.4]
  wire [8:0] _T_2807; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2810.4]
  wire  _T_2808; // @[Bitwise.scala 50:65:@2811.4]
  wire  _T_2809; // @[Bitwise.scala 50:65:@2812.4]
  wire  _T_2810; // @[Bitwise.scala 50:65:@2813.4]
  wire  _T_2811; // @[Bitwise.scala 50:65:@2814.4]
  wire  _T_2812; // @[Bitwise.scala 50:65:@2815.4]
  wire  _T_2813; // @[Bitwise.scala 50:65:@2816.4]
  wire  _T_2814; // @[Bitwise.scala 50:65:@2817.4]
  wire  _T_2815; // @[Bitwise.scala 50:65:@2818.4]
  wire  _T_2816; // @[Bitwise.scala 50:65:@2819.4]
  wire [1:0] _T_2817; // @[Bitwise.scala 48:55:@2820.4]
  wire [1:0] _T_2818; // @[Bitwise.scala 48:55:@2821.4]
  wire [2:0] _T_2819; // @[Bitwise.scala 48:55:@2822.4]
  wire [1:0] _T_2820; // @[Bitwise.scala 48:55:@2823.4]
  wire [1:0] _T_2821; // @[Bitwise.scala 48:55:@2824.4]
  wire [1:0] _GEN_550; // @[Bitwise.scala 48:55:@2825.4]
  wire [2:0] _T_2822; // @[Bitwise.scala 48:55:@2825.4]
  wire [2:0] _GEN_551; // @[Bitwise.scala 48:55:@2826.4]
  wire [3:0] _T_2823; // @[Bitwise.scala 48:55:@2826.4]
  wire [3:0] _GEN_552; // @[Bitwise.scala 48:55:@2827.4]
  wire [4:0] _T_2824; // @[Bitwise.scala 48:55:@2827.4]
  wire [9:0] _T_2888; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2892.4]
  wire  _T_2889; // @[Bitwise.scala 50:65:@2893.4]
  wire  _T_2890; // @[Bitwise.scala 50:65:@2894.4]
  wire  _T_2891; // @[Bitwise.scala 50:65:@2895.4]
  wire  _T_2892; // @[Bitwise.scala 50:65:@2896.4]
  wire  _T_2893; // @[Bitwise.scala 50:65:@2897.4]
  wire  _T_2894; // @[Bitwise.scala 50:65:@2898.4]
  wire  _T_2895; // @[Bitwise.scala 50:65:@2899.4]
  wire  _T_2896; // @[Bitwise.scala 50:65:@2900.4]
  wire  _T_2897; // @[Bitwise.scala 50:65:@2901.4]
  wire  _T_2898; // @[Bitwise.scala 50:65:@2902.4]
  wire [1:0] _T_2899; // @[Bitwise.scala 48:55:@2903.4]
  wire [1:0] _T_2900; // @[Bitwise.scala 48:55:@2904.4]
  wire [1:0] _GEN_553; // @[Bitwise.scala 48:55:@2905.4]
  wire [2:0] _T_2901; // @[Bitwise.scala 48:55:@2905.4]
  wire [2:0] _GEN_554; // @[Bitwise.scala 48:55:@2906.4]
  wire [3:0] _T_2902; // @[Bitwise.scala 48:55:@2906.4]
  wire [1:0] _T_2903; // @[Bitwise.scala 48:55:@2907.4]
  wire [1:0] _T_2904; // @[Bitwise.scala 48:55:@2908.4]
  wire [1:0] _GEN_555; // @[Bitwise.scala 48:55:@2909.4]
  wire [2:0] _T_2905; // @[Bitwise.scala 48:55:@2909.4]
  wire [2:0] _GEN_556; // @[Bitwise.scala 48:55:@2910.4]
  wire [3:0] _T_2906; // @[Bitwise.scala 48:55:@2910.4]
  wire [4:0] _T_2907; // @[Bitwise.scala 48:55:@2911.4]
  wire [10:0] _T_2971; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2976.4]
  wire  _T_2972; // @[Bitwise.scala 50:65:@2977.4]
  wire  _T_2973; // @[Bitwise.scala 50:65:@2978.4]
  wire  _T_2974; // @[Bitwise.scala 50:65:@2979.4]
  wire  _T_2975; // @[Bitwise.scala 50:65:@2980.4]
  wire  _T_2976; // @[Bitwise.scala 50:65:@2981.4]
  wire  _T_2977; // @[Bitwise.scala 50:65:@2982.4]
  wire  _T_2978; // @[Bitwise.scala 50:65:@2983.4]
  wire  _T_2979; // @[Bitwise.scala 50:65:@2984.4]
  wire  _T_2980; // @[Bitwise.scala 50:65:@2985.4]
  wire  _T_2981; // @[Bitwise.scala 50:65:@2986.4]
  wire  _T_2982; // @[Bitwise.scala 50:65:@2987.4]
  wire [1:0] _T_2983; // @[Bitwise.scala 48:55:@2988.4]
  wire [1:0] _T_2984; // @[Bitwise.scala 48:55:@2989.4]
  wire [1:0] _GEN_557; // @[Bitwise.scala 48:55:@2990.4]
  wire [2:0] _T_2985; // @[Bitwise.scala 48:55:@2990.4]
  wire [2:0] _GEN_558; // @[Bitwise.scala 48:55:@2991.4]
  wire [3:0] _T_2986; // @[Bitwise.scala 48:55:@2991.4]
  wire [1:0] _T_2987; // @[Bitwise.scala 48:55:@2992.4]
  wire [1:0] _GEN_559; // @[Bitwise.scala 48:55:@2993.4]
  wire [2:0] _T_2988; // @[Bitwise.scala 48:55:@2993.4]
  wire [1:0] _T_2989; // @[Bitwise.scala 48:55:@2994.4]
  wire [1:0] _GEN_560; // @[Bitwise.scala 48:55:@2995.4]
  wire [2:0] _T_2990; // @[Bitwise.scala 48:55:@2995.4]
  wire [3:0] _T_2991; // @[Bitwise.scala 48:55:@2996.4]
  wire [4:0] _T_2992; // @[Bitwise.scala 48:55:@2997.4]
  wire [11:0] _T_3056; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3062.4]
  wire  _T_3057; // @[Bitwise.scala 50:65:@3063.4]
  wire  _T_3058; // @[Bitwise.scala 50:65:@3064.4]
  wire  _T_3059; // @[Bitwise.scala 50:65:@3065.4]
  wire  _T_3060; // @[Bitwise.scala 50:65:@3066.4]
  wire  _T_3061; // @[Bitwise.scala 50:65:@3067.4]
  wire  _T_3062; // @[Bitwise.scala 50:65:@3068.4]
  wire  _T_3063; // @[Bitwise.scala 50:65:@3069.4]
  wire  _T_3064; // @[Bitwise.scala 50:65:@3070.4]
  wire  _T_3065; // @[Bitwise.scala 50:65:@3071.4]
  wire  _T_3066; // @[Bitwise.scala 50:65:@3072.4]
  wire  _T_3067; // @[Bitwise.scala 50:65:@3073.4]
  wire  _T_3068; // @[Bitwise.scala 50:65:@3074.4]
  wire [1:0] _T_3069; // @[Bitwise.scala 48:55:@3075.4]
  wire [1:0] _GEN_561; // @[Bitwise.scala 48:55:@3076.4]
  wire [2:0] _T_3070; // @[Bitwise.scala 48:55:@3076.4]
  wire [1:0] _T_3071; // @[Bitwise.scala 48:55:@3077.4]
  wire [1:0] _GEN_562; // @[Bitwise.scala 48:55:@3078.4]
  wire [2:0] _T_3072; // @[Bitwise.scala 48:55:@3078.4]
  wire [3:0] _T_3073; // @[Bitwise.scala 48:55:@3079.4]
  wire [1:0] _T_3074; // @[Bitwise.scala 48:55:@3080.4]
  wire [1:0] _GEN_563; // @[Bitwise.scala 48:55:@3081.4]
  wire [2:0] _T_3075; // @[Bitwise.scala 48:55:@3081.4]
  wire [1:0] _T_3076; // @[Bitwise.scala 48:55:@3082.4]
  wire [1:0] _GEN_564; // @[Bitwise.scala 48:55:@3083.4]
  wire [2:0] _T_3077; // @[Bitwise.scala 48:55:@3083.4]
  wire [3:0] _T_3078; // @[Bitwise.scala 48:55:@3084.4]
  wire [4:0] _T_3079; // @[Bitwise.scala 48:55:@3085.4]
  wire [12:0] _T_3143; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3150.4]
  wire  _T_3144; // @[Bitwise.scala 50:65:@3151.4]
  wire  _T_3145; // @[Bitwise.scala 50:65:@3152.4]
  wire  _T_3146; // @[Bitwise.scala 50:65:@3153.4]
  wire  _T_3147; // @[Bitwise.scala 50:65:@3154.4]
  wire  _T_3148; // @[Bitwise.scala 50:65:@3155.4]
  wire  _T_3149; // @[Bitwise.scala 50:65:@3156.4]
  wire  _T_3150; // @[Bitwise.scala 50:65:@3157.4]
  wire  _T_3151; // @[Bitwise.scala 50:65:@3158.4]
  wire  _T_3152; // @[Bitwise.scala 50:65:@3159.4]
  wire  _T_3153; // @[Bitwise.scala 50:65:@3160.4]
  wire  _T_3154; // @[Bitwise.scala 50:65:@3161.4]
  wire  _T_3155; // @[Bitwise.scala 50:65:@3162.4]
  wire  _T_3156; // @[Bitwise.scala 50:65:@3163.4]
  wire [1:0] _T_3157; // @[Bitwise.scala 48:55:@3164.4]
  wire [1:0] _GEN_565; // @[Bitwise.scala 48:55:@3165.4]
  wire [2:0] _T_3158; // @[Bitwise.scala 48:55:@3165.4]
  wire [1:0] _T_3159; // @[Bitwise.scala 48:55:@3166.4]
  wire [1:0] _GEN_566; // @[Bitwise.scala 48:55:@3167.4]
  wire [2:0] _T_3160; // @[Bitwise.scala 48:55:@3167.4]
  wire [3:0] _T_3161; // @[Bitwise.scala 48:55:@3168.4]
  wire [1:0] _T_3162; // @[Bitwise.scala 48:55:@3169.4]
  wire [1:0] _GEN_567; // @[Bitwise.scala 48:55:@3170.4]
  wire [2:0] _T_3163; // @[Bitwise.scala 48:55:@3170.4]
  wire [1:0] _T_3164; // @[Bitwise.scala 48:55:@3171.4]
  wire [1:0] _T_3165; // @[Bitwise.scala 48:55:@3172.4]
  wire [2:0] _T_3166; // @[Bitwise.scala 48:55:@3173.4]
  wire [3:0] _T_3167; // @[Bitwise.scala 48:55:@3174.4]
  wire [4:0] _T_3168; // @[Bitwise.scala 48:55:@3175.4]
  wire [13:0] _T_3232; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3240.4]
  wire  _T_3233; // @[Bitwise.scala 50:65:@3241.4]
  wire  _T_3234; // @[Bitwise.scala 50:65:@3242.4]
  wire  _T_3235; // @[Bitwise.scala 50:65:@3243.4]
  wire  _T_3236; // @[Bitwise.scala 50:65:@3244.4]
  wire  _T_3237; // @[Bitwise.scala 50:65:@3245.4]
  wire  _T_3238; // @[Bitwise.scala 50:65:@3246.4]
  wire  _T_3239; // @[Bitwise.scala 50:65:@3247.4]
  wire  _T_3240; // @[Bitwise.scala 50:65:@3248.4]
  wire  _T_3241; // @[Bitwise.scala 50:65:@3249.4]
  wire  _T_3242; // @[Bitwise.scala 50:65:@3250.4]
  wire  _T_3243; // @[Bitwise.scala 50:65:@3251.4]
  wire  _T_3244; // @[Bitwise.scala 50:65:@3252.4]
  wire  _T_3245; // @[Bitwise.scala 50:65:@3253.4]
  wire  _T_3246; // @[Bitwise.scala 50:65:@3254.4]
  wire [1:0] _T_3247; // @[Bitwise.scala 48:55:@3255.4]
  wire [1:0] _GEN_568; // @[Bitwise.scala 48:55:@3256.4]
  wire [2:0] _T_3248; // @[Bitwise.scala 48:55:@3256.4]
  wire [1:0] _T_3249; // @[Bitwise.scala 48:55:@3257.4]
  wire [1:0] _T_3250; // @[Bitwise.scala 48:55:@3258.4]
  wire [2:0] _T_3251; // @[Bitwise.scala 48:55:@3259.4]
  wire [3:0] _T_3252; // @[Bitwise.scala 48:55:@3260.4]
  wire [1:0] _T_3253; // @[Bitwise.scala 48:55:@3261.4]
  wire [1:0] _GEN_569; // @[Bitwise.scala 48:55:@3262.4]
  wire [2:0] _T_3254; // @[Bitwise.scala 48:55:@3262.4]
  wire [1:0] _T_3255; // @[Bitwise.scala 48:55:@3263.4]
  wire [1:0] _T_3256; // @[Bitwise.scala 48:55:@3264.4]
  wire [2:0] _T_3257; // @[Bitwise.scala 48:55:@3265.4]
  wire [3:0] _T_3258; // @[Bitwise.scala 48:55:@3266.4]
  wire [4:0] _T_3259; // @[Bitwise.scala 48:55:@3267.4]
  wire [14:0] _T_3323; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3332.4]
  wire  _T_3324; // @[Bitwise.scala 50:65:@3333.4]
  wire  _T_3325; // @[Bitwise.scala 50:65:@3334.4]
  wire  _T_3326; // @[Bitwise.scala 50:65:@3335.4]
  wire  _T_3327; // @[Bitwise.scala 50:65:@3336.4]
  wire  _T_3328; // @[Bitwise.scala 50:65:@3337.4]
  wire  _T_3329; // @[Bitwise.scala 50:65:@3338.4]
  wire  _T_3330; // @[Bitwise.scala 50:65:@3339.4]
  wire  _T_3331; // @[Bitwise.scala 50:65:@3340.4]
  wire  _T_3332; // @[Bitwise.scala 50:65:@3341.4]
  wire  _T_3333; // @[Bitwise.scala 50:65:@3342.4]
  wire  _T_3334; // @[Bitwise.scala 50:65:@3343.4]
  wire  _T_3335; // @[Bitwise.scala 50:65:@3344.4]
  wire  _T_3336; // @[Bitwise.scala 50:65:@3345.4]
  wire  _T_3337; // @[Bitwise.scala 50:65:@3346.4]
  wire  _T_3338; // @[Bitwise.scala 50:65:@3347.4]
  wire [1:0] _T_3339; // @[Bitwise.scala 48:55:@3348.4]
  wire [1:0] _GEN_570; // @[Bitwise.scala 48:55:@3349.4]
  wire [2:0] _T_3340; // @[Bitwise.scala 48:55:@3349.4]
  wire [1:0] _T_3341; // @[Bitwise.scala 48:55:@3350.4]
  wire [1:0] _T_3342; // @[Bitwise.scala 48:55:@3351.4]
  wire [2:0] _T_3343; // @[Bitwise.scala 48:55:@3352.4]
  wire [3:0] _T_3344; // @[Bitwise.scala 48:55:@3353.4]
  wire [1:0] _T_3345; // @[Bitwise.scala 48:55:@3354.4]
  wire [1:0] _T_3346; // @[Bitwise.scala 48:55:@3355.4]
  wire [2:0] _T_3347; // @[Bitwise.scala 48:55:@3356.4]
  wire [1:0] _T_3348; // @[Bitwise.scala 48:55:@3357.4]
  wire [1:0] _T_3349; // @[Bitwise.scala 48:55:@3358.4]
  wire [2:0] _T_3350; // @[Bitwise.scala 48:55:@3359.4]
  wire [3:0] _T_3351; // @[Bitwise.scala 48:55:@3360.4]
  wire [4:0] _T_3352; // @[Bitwise.scala 48:55:@3361.4]
  wire [15:0] _T_3416; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3426.4]
  wire  _T_3417; // @[Bitwise.scala 50:65:@3427.4]
  wire  _T_3418; // @[Bitwise.scala 50:65:@3428.4]
  wire  _T_3419; // @[Bitwise.scala 50:65:@3429.4]
  wire  _T_3420; // @[Bitwise.scala 50:65:@3430.4]
  wire  _T_3421; // @[Bitwise.scala 50:65:@3431.4]
  wire  _T_3422; // @[Bitwise.scala 50:65:@3432.4]
  wire  _T_3423; // @[Bitwise.scala 50:65:@3433.4]
  wire  _T_3424; // @[Bitwise.scala 50:65:@3434.4]
  wire  _T_3425; // @[Bitwise.scala 50:65:@3435.4]
  wire  _T_3426; // @[Bitwise.scala 50:65:@3436.4]
  wire  _T_3427; // @[Bitwise.scala 50:65:@3437.4]
  wire  _T_3428; // @[Bitwise.scala 50:65:@3438.4]
  wire  _T_3429; // @[Bitwise.scala 50:65:@3439.4]
  wire  _T_3430; // @[Bitwise.scala 50:65:@3440.4]
  wire  _T_3431; // @[Bitwise.scala 50:65:@3441.4]
  wire  _T_3432; // @[Bitwise.scala 50:65:@3442.4]
  wire [1:0] _T_3433; // @[Bitwise.scala 48:55:@3443.4]
  wire [1:0] _T_3434; // @[Bitwise.scala 48:55:@3444.4]
  wire [2:0] _T_3435; // @[Bitwise.scala 48:55:@3445.4]
  wire [1:0] _T_3436; // @[Bitwise.scala 48:55:@3446.4]
  wire [1:0] _T_3437; // @[Bitwise.scala 48:55:@3447.4]
  wire [2:0] _T_3438; // @[Bitwise.scala 48:55:@3448.4]
  wire [3:0] _T_3439; // @[Bitwise.scala 48:55:@3449.4]
  wire [1:0] _T_3440; // @[Bitwise.scala 48:55:@3450.4]
  wire [1:0] _T_3441; // @[Bitwise.scala 48:55:@3451.4]
  wire [2:0] _T_3442; // @[Bitwise.scala 48:55:@3452.4]
  wire [1:0] _T_3443; // @[Bitwise.scala 48:55:@3453.4]
  wire [1:0] _T_3444; // @[Bitwise.scala 48:55:@3454.4]
  wire [2:0] _T_3445; // @[Bitwise.scala 48:55:@3455.4]
  wire [3:0] _T_3446; // @[Bitwise.scala 48:55:@3456.4]
  wire [4:0] _T_3447; // @[Bitwise.scala 48:55:@3457.4]
  wire [16:0] _T_3511; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3522.4]
  wire  _T_3512; // @[Bitwise.scala 50:65:@3523.4]
  wire  _T_3513; // @[Bitwise.scala 50:65:@3524.4]
  wire  _T_3514; // @[Bitwise.scala 50:65:@3525.4]
  wire  _T_3515; // @[Bitwise.scala 50:65:@3526.4]
  wire  _T_3516; // @[Bitwise.scala 50:65:@3527.4]
  wire  _T_3517; // @[Bitwise.scala 50:65:@3528.4]
  wire  _T_3518; // @[Bitwise.scala 50:65:@3529.4]
  wire  _T_3519; // @[Bitwise.scala 50:65:@3530.4]
  wire  _T_3520; // @[Bitwise.scala 50:65:@3531.4]
  wire  _T_3521; // @[Bitwise.scala 50:65:@3532.4]
  wire  _T_3522; // @[Bitwise.scala 50:65:@3533.4]
  wire  _T_3523; // @[Bitwise.scala 50:65:@3534.4]
  wire  _T_3524; // @[Bitwise.scala 50:65:@3535.4]
  wire  _T_3525; // @[Bitwise.scala 50:65:@3536.4]
  wire  _T_3526; // @[Bitwise.scala 50:65:@3537.4]
  wire  _T_3527; // @[Bitwise.scala 50:65:@3538.4]
  wire  _T_3528; // @[Bitwise.scala 50:65:@3539.4]
  wire [1:0] _T_3529; // @[Bitwise.scala 48:55:@3540.4]
  wire [1:0] _T_3530; // @[Bitwise.scala 48:55:@3541.4]
  wire [2:0] _T_3531; // @[Bitwise.scala 48:55:@3542.4]
  wire [1:0] _T_3532; // @[Bitwise.scala 48:55:@3543.4]
  wire [1:0] _T_3533; // @[Bitwise.scala 48:55:@3544.4]
  wire [2:0] _T_3534; // @[Bitwise.scala 48:55:@3545.4]
  wire [3:0] _T_3535; // @[Bitwise.scala 48:55:@3546.4]
  wire [1:0] _T_3536; // @[Bitwise.scala 48:55:@3547.4]
  wire [1:0] _T_3537; // @[Bitwise.scala 48:55:@3548.4]
  wire [2:0] _T_3538; // @[Bitwise.scala 48:55:@3549.4]
  wire [1:0] _T_3539; // @[Bitwise.scala 48:55:@3550.4]
  wire [1:0] _T_3540; // @[Bitwise.scala 48:55:@3551.4]
  wire [1:0] _GEN_571; // @[Bitwise.scala 48:55:@3552.4]
  wire [2:0] _T_3541; // @[Bitwise.scala 48:55:@3552.4]
  wire [2:0] _GEN_572; // @[Bitwise.scala 48:55:@3553.4]
  wire [3:0] _T_3542; // @[Bitwise.scala 48:55:@3553.4]
  wire [3:0] _GEN_573; // @[Bitwise.scala 48:55:@3554.4]
  wire [4:0] _T_3543; // @[Bitwise.scala 48:55:@3554.4]
  wire [4:0] _GEN_574; // @[Bitwise.scala 48:55:@3555.4]
  wire [5:0] _T_3544; // @[Bitwise.scala 48:55:@3555.4]
  wire [17:0] _T_3608; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3620.4]
  wire  _T_3609; // @[Bitwise.scala 50:65:@3621.4]
  wire  _T_3610; // @[Bitwise.scala 50:65:@3622.4]
  wire  _T_3611; // @[Bitwise.scala 50:65:@3623.4]
  wire  _T_3612; // @[Bitwise.scala 50:65:@3624.4]
  wire  _T_3613; // @[Bitwise.scala 50:65:@3625.4]
  wire  _T_3614; // @[Bitwise.scala 50:65:@3626.4]
  wire  _T_3615; // @[Bitwise.scala 50:65:@3627.4]
  wire  _T_3616; // @[Bitwise.scala 50:65:@3628.4]
  wire  _T_3617; // @[Bitwise.scala 50:65:@3629.4]
  wire  _T_3618; // @[Bitwise.scala 50:65:@3630.4]
  wire  _T_3619; // @[Bitwise.scala 50:65:@3631.4]
  wire  _T_3620; // @[Bitwise.scala 50:65:@3632.4]
  wire  _T_3621; // @[Bitwise.scala 50:65:@3633.4]
  wire  _T_3622; // @[Bitwise.scala 50:65:@3634.4]
  wire  _T_3623; // @[Bitwise.scala 50:65:@3635.4]
  wire  _T_3624; // @[Bitwise.scala 50:65:@3636.4]
  wire  _T_3625; // @[Bitwise.scala 50:65:@3637.4]
  wire  _T_3626; // @[Bitwise.scala 50:65:@3638.4]
  wire [1:0] _T_3627; // @[Bitwise.scala 48:55:@3639.4]
  wire [1:0] _T_3628; // @[Bitwise.scala 48:55:@3640.4]
  wire [2:0] _T_3629; // @[Bitwise.scala 48:55:@3641.4]
  wire [1:0] _T_3630; // @[Bitwise.scala 48:55:@3642.4]
  wire [1:0] _T_3631; // @[Bitwise.scala 48:55:@3643.4]
  wire [1:0] _GEN_575; // @[Bitwise.scala 48:55:@3644.4]
  wire [2:0] _T_3632; // @[Bitwise.scala 48:55:@3644.4]
  wire [2:0] _GEN_576; // @[Bitwise.scala 48:55:@3645.4]
  wire [3:0] _T_3633; // @[Bitwise.scala 48:55:@3645.4]
  wire [3:0] _GEN_577; // @[Bitwise.scala 48:55:@3646.4]
  wire [4:0] _T_3634; // @[Bitwise.scala 48:55:@3646.4]
  wire [1:0] _T_3635; // @[Bitwise.scala 48:55:@3647.4]
  wire [1:0] _T_3636; // @[Bitwise.scala 48:55:@3648.4]
  wire [2:0] _T_3637; // @[Bitwise.scala 48:55:@3649.4]
  wire [1:0] _T_3638; // @[Bitwise.scala 48:55:@3650.4]
  wire [1:0] _T_3639; // @[Bitwise.scala 48:55:@3651.4]
  wire [1:0] _GEN_578; // @[Bitwise.scala 48:55:@3652.4]
  wire [2:0] _T_3640; // @[Bitwise.scala 48:55:@3652.4]
  wire [2:0] _GEN_579; // @[Bitwise.scala 48:55:@3653.4]
  wire [3:0] _T_3641; // @[Bitwise.scala 48:55:@3653.4]
  wire [3:0] _GEN_580; // @[Bitwise.scala 48:55:@3654.4]
  wire [4:0] _T_3642; // @[Bitwise.scala 48:55:@3654.4]
  wire [5:0] _T_3643; // @[Bitwise.scala 48:55:@3655.4]
  wire [18:0] _T_3707; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3720.4]
  wire  _T_3708; // @[Bitwise.scala 50:65:@3721.4]
  wire  _T_3709; // @[Bitwise.scala 50:65:@3722.4]
  wire  _T_3710; // @[Bitwise.scala 50:65:@3723.4]
  wire  _T_3711; // @[Bitwise.scala 50:65:@3724.4]
  wire  _T_3712; // @[Bitwise.scala 50:65:@3725.4]
  wire  _T_3713; // @[Bitwise.scala 50:65:@3726.4]
  wire  _T_3714; // @[Bitwise.scala 50:65:@3727.4]
  wire  _T_3715; // @[Bitwise.scala 50:65:@3728.4]
  wire  _T_3716; // @[Bitwise.scala 50:65:@3729.4]
  wire  _T_3717; // @[Bitwise.scala 50:65:@3730.4]
  wire  _T_3718; // @[Bitwise.scala 50:65:@3731.4]
  wire  _T_3719; // @[Bitwise.scala 50:65:@3732.4]
  wire  _T_3720; // @[Bitwise.scala 50:65:@3733.4]
  wire  _T_3721; // @[Bitwise.scala 50:65:@3734.4]
  wire  _T_3722; // @[Bitwise.scala 50:65:@3735.4]
  wire  _T_3723; // @[Bitwise.scala 50:65:@3736.4]
  wire  _T_3724; // @[Bitwise.scala 50:65:@3737.4]
  wire  _T_3725; // @[Bitwise.scala 50:65:@3738.4]
  wire  _T_3726; // @[Bitwise.scala 50:65:@3739.4]
  wire [1:0] _T_3727; // @[Bitwise.scala 48:55:@3740.4]
  wire [1:0] _T_3728; // @[Bitwise.scala 48:55:@3741.4]
  wire [2:0] _T_3729; // @[Bitwise.scala 48:55:@3742.4]
  wire [1:0] _T_3730; // @[Bitwise.scala 48:55:@3743.4]
  wire [1:0] _T_3731; // @[Bitwise.scala 48:55:@3744.4]
  wire [1:0] _GEN_581; // @[Bitwise.scala 48:55:@3745.4]
  wire [2:0] _T_3732; // @[Bitwise.scala 48:55:@3745.4]
  wire [2:0] _GEN_582; // @[Bitwise.scala 48:55:@3746.4]
  wire [3:0] _T_3733; // @[Bitwise.scala 48:55:@3746.4]
  wire [3:0] _GEN_583; // @[Bitwise.scala 48:55:@3747.4]
  wire [4:0] _T_3734; // @[Bitwise.scala 48:55:@3747.4]
  wire [1:0] _T_3735; // @[Bitwise.scala 48:55:@3748.4]
  wire [1:0] _T_3736; // @[Bitwise.scala 48:55:@3749.4]
  wire [1:0] _GEN_584; // @[Bitwise.scala 48:55:@3750.4]
  wire [2:0] _T_3737; // @[Bitwise.scala 48:55:@3750.4]
  wire [2:0] _GEN_585; // @[Bitwise.scala 48:55:@3751.4]
  wire [3:0] _T_3738; // @[Bitwise.scala 48:55:@3751.4]
  wire [1:0] _T_3739; // @[Bitwise.scala 48:55:@3752.4]
  wire [1:0] _T_3740; // @[Bitwise.scala 48:55:@3753.4]
  wire [1:0] _GEN_586; // @[Bitwise.scala 48:55:@3754.4]
  wire [2:0] _T_3741; // @[Bitwise.scala 48:55:@3754.4]
  wire [2:0] _GEN_587; // @[Bitwise.scala 48:55:@3755.4]
  wire [3:0] _T_3742; // @[Bitwise.scala 48:55:@3755.4]
  wire [4:0] _T_3743; // @[Bitwise.scala 48:55:@3756.4]
  wire [5:0] _T_3744; // @[Bitwise.scala 48:55:@3757.4]
  wire [19:0] _T_3808; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3822.4]
  wire  _T_3809; // @[Bitwise.scala 50:65:@3823.4]
  wire  _T_3810; // @[Bitwise.scala 50:65:@3824.4]
  wire  _T_3811; // @[Bitwise.scala 50:65:@3825.4]
  wire  _T_3812; // @[Bitwise.scala 50:65:@3826.4]
  wire  _T_3813; // @[Bitwise.scala 50:65:@3827.4]
  wire  _T_3814; // @[Bitwise.scala 50:65:@3828.4]
  wire  _T_3815; // @[Bitwise.scala 50:65:@3829.4]
  wire  _T_3816; // @[Bitwise.scala 50:65:@3830.4]
  wire  _T_3817; // @[Bitwise.scala 50:65:@3831.4]
  wire  _T_3818; // @[Bitwise.scala 50:65:@3832.4]
  wire  _T_3819; // @[Bitwise.scala 50:65:@3833.4]
  wire  _T_3820; // @[Bitwise.scala 50:65:@3834.4]
  wire  _T_3821; // @[Bitwise.scala 50:65:@3835.4]
  wire  _T_3822; // @[Bitwise.scala 50:65:@3836.4]
  wire  _T_3823; // @[Bitwise.scala 50:65:@3837.4]
  wire  _T_3824; // @[Bitwise.scala 50:65:@3838.4]
  wire  _T_3825; // @[Bitwise.scala 50:65:@3839.4]
  wire  _T_3826; // @[Bitwise.scala 50:65:@3840.4]
  wire  _T_3827; // @[Bitwise.scala 50:65:@3841.4]
  wire  _T_3828; // @[Bitwise.scala 50:65:@3842.4]
  wire [1:0] _T_3829; // @[Bitwise.scala 48:55:@3843.4]
  wire [1:0] _T_3830; // @[Bitwise.scala 48:55:@3844.4]
  wire [1:0] _GEN_588; // @[Bitwise.scala 48:55:@3845.4]
  wire [2:0] _T_3831; // @[Bitwise.scala 48:55:@3845.4]
  wire [2:0] _GEN_589; // @[Bitwise.scala 48:55:@3846.4]
  wire [3:0] _T_3832; // @[Bitwise.scala 48:55:@3846.4]
  wire [1:0] _T_3833; // @[Bitwise.scala 48:55:@3847.4]
  wire [1:0] _T_3834; // @[Bitwise.scala 48:55:@3848.4]
  wire [1:0] _GEN_590; // @[Bitwise.scala 48:55:@3849.4]
  wire [2:0] _T_3835; // @[Bitwise.scala 48:55:@3849.4]
  wire [2:0] _GEN_591; // @[Bitwise.scala 48:55:@3850.4]
  wire [3:0] _T_3836; // @[Bitwise.scala 48:55:@3850.4]
  wire [4:0] _T_3837; // @[Bitwise.scala 48:55:@3851.4]
  wire [1:0] _T_3838; // @[Bitwise.scala 48:55:@3852.4]
  wire [1:0] _T_3839; // @[Bitwise.scala 48:55:@3853.4]
  wire [1:0] _GEN_592; // @[Bitwise.scala 48:55:@3854.4]
  wire [2:0] _T_3840; // @[Bitwise.scala 48:55:@3854.4]
  wire [2:0] _GEN_593; // @[Bitwise.scala 48:55:@3855.4]
  wire [3:0] _T_3841; // @[Bitwise.scala 48:55:@3855.4]
  wire [1:0] _T_3842; // @[Bitwise.scala 48:55:@3856.4]
  wire [1:0] _T_3843; // @[Bitwise.scala 48:55:@3857.4]
  wire [1:0] _GEN_594; // @[Bitwise.scala 48:55:@3858.4]
  wire [2:0] _T_3844; // @[Bitwise.scala 48:55:@3858.4]
  wire [2:0] _GEN_595; // @[Bitwise.scala 48:55:@3859.4]
  wire [3:0] _T_3845; // @[Bitwise.scala 48:55:@3859.4]
  wire [4:0] _T_3846; // @[Bitwise.scala 48:55:@3860.4]
  wire [5:0] _T_3847; // @[Bitwise.scala 48:55:@3861.4]
  wire [20:0] _T_3911; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3926.4]
  wire  _T_3912; // @[Bitwise.scala 50:65:@3927.4]
  wire  _T_3913; // @[Bitwise.scala 50:65:@3928.4]
  wire  _T_3914; // @[Bitwise.scala 50:65:@3929.4]
  wire  _T_3915; // @[Bitwise.scala 50:65:@3930.4]
  wire  _T_3916; // @[Bitwise.scala 50:65:@3931.4]
  wire  _T_3917; // @[Bitwise.scala 50:65:@3932.4]
  wire  _T_3918; // @[Bitwise.scala 50:65:@3933.4]
  wire  _T_3919; // @[Bitwise.scala 50:65:@3934.4]
  wire  _T_3920; // @[Bitwise.scala 50:65:@3935.4]
  wire  _T_3921; // @[Bitwise.scala 50:65:@3936.4]
  wire  _T_3922; // @[Bitwise.scala 50:65:@3937.4]
  wire  _T_3923; // @[Bitwise.scala 50:65:@3938.4]
  wire  _T_3924; // @[Bitwise.scala 50:65:@3939.4]
  wire  _T_3925; // @[Bitwise.scala 50:65:@3940.4]
  wire  _T_3926; // @[Bitwise.scala 50:65:@3941.4]
  wire  _T_3927; // @[Bitwise.scala 50:65:@3942.4]
  wire  _T_3928; // @[Bitwise.scala 50:65:@3943.4]
  wire  _T_3929; // @[Bitwise.scala 50:65:@3944.4]
  wire  _T_3930; // @[Bitwise.scala 50:65:@3945.4]
  wire  _T_3931; // @[Bitwise.scala 50:65:@3946.4]
  wire  _T_3932; // @[Bitwise.scala 50:65:@3947.4]
  wire [1:0] _T_3933; // @[Bitwise.scala 48:55:@3948.4]
  wire [1:0] _T_3934; // @[Bitwise.scala 48:55:@3949.4]
  wire [1:0] _GEN_596; // @[Bitwise.scala 48:55:@3950.4]
  wire [2:0] _T_3935; // @[Bitwise.scala 48:55:@3950.4]
  wire [2:0] _GEN_597; // @[Bitwise.scala 48:55:@3951.4]
  wire [3:0] _T_3936; // @[Bitwise.scala 48:55:@3951.4]
  wire [1:0] _T_3937; // @[Bitwise.scala 48:55:@3952.4]
  wire [1:0] _T_3938; // @[Bitwise.scala 48:55:@3953.4]
  wire [1:0] _GEN_598; // @[Bitwise.scala 48:55:@3954.4]
  wire [2:0] _T_3939; // @[Bitwise.scala 48:55:@3954.4]
  wire [2:0] _GEN_599; // @[Bitwise.scala 48:55:@3955.4]
  wire [3:0] _T_3940; // @[Bitwise.scala 48:55:@3955.4]
  wire [4:0] _T_3941; // @[Bitwise.scala 48:55:@3956.4]
  wire [1:0] _T_3942; // @[Bitwise.scala 48:55:@3957.4]
  wire [1:0] _T_3943; // @[Bitwise.scala 48:55:@3958.4]
  wire [1:0] _GEN_600; // @[Bitwise.scala 48:55:@3959.4]
  wire [2:0] _T_3944; // @[Bitwise.scala 48:55:@3959.4]
  wire [2:0] _GEN_601; // @[Bitwise.scala 48:55:@3960.4]
  wire [3:0] _T_3945; // @[Bitwise.scala 48:55:@3960.4]
  wire [1:0] _T_3946; // @[Bitwise.scala 48:55:@3961.4]
  wire [1:0] _GEN_602; // @[Bitwise.scala 48:55:@3962.4]
  wire [2:0] _T_3947; // @[Bitwise.scala 48:55:@3962.4]
  wire [1:0] _T_3948; // @[Bitwise.scala 48:55:@3963.4]
  wire [1:0] _GEN_603; // @[Bitwise.scala 48:55:@3964.4]
  wire [2:0] _T_3949; // @[Bitwise.scala 48:55:@3964.4]
  wire [3:0] _T_3950; // @[Bitwise.scala 48:55:@3965.4]
  wire [4:0] _T_3951; // @[Bitwise.scala 48:55:@3966.4]
  wire [5:0] _T_3952; // @[Bitwise.scala 48:55:@3967.4]
  wire [21:0] _T_4016; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4032.4]
  wire  _T_4017; // @[Bitwise.scala 50:65:@4033.4]
  wire  _T_4018; // @[Bitwise.scala 50:65:@4034.4]
  wire  _T_4019; // @[Bitwise.scala 50:65:@4035.4]
  wire  _T_4020; // @[Bitwise.scala 50:65:@4036.4]
  wire  _T_4021; // @[Bitwise.scala 50:65:@4037.4]
  wire  _T_4022; // @[Bitwise.scala 50:65:@4038.4]
  wire  _T_4023; // @[Bitwise.scala 50:65:@4039.4]
  wire  _T_4024; // @[Bitwise.scala 50:65:@4040.4]
  wire  _T_4025; // @[Bitwise.scala 50:65:@4041.4]
  wire  _T_4026; // @[Bitwise.scala 50:65:@4042.4]
  wire  _T_4027; // @[Bitwise.scala 50:65:@4043.4]
  wire  _T_4028; // @[Bitwise.scala 50:65:@4044.4]
  wire  _T_4029; // @[Bitwise.scala 50:65:@4045.4]
  wire  _T_4030; // @[Bitwise.scala 50:65:@4046.4]
  wire  _T_4031; // @[Bitwise.scala 50:65:@4047.4]
  wire  _T_4032; // @[Bitwise.scala 50:65:@4048.4]
  wire  _T_4033; // @[Bitwise.scala 50:65:@4049.4]
  wire  _T_4034; // @[Bitwise.scala 50:65:@4050.4]
  wire  _T_4035; // @[Bitwise.scala 50:65:@4051.4]
  wire  _T_4036; // @[Bitwise.scala 50:65:@4052.4]
  wire  _T_4037; // @[Bitwise.scala 50:65:@4053.4]
  wire  _T_4038; // @[Bitwise.scala 50:65:@4054.4]
  wire [1:0] _T_4039; // @[Bitwise.scala 48:55:@4055.4]
  wire [1:0] _T_4040; // @[Bitwise.scala 48:55:@4056.4]
  wire [1:0] _GEN_604; // @[Bitwise.scala 48:55:@4057.4]
  wire [2:0] _T_4041; // @[Bitwise.scala 48:55:@4057.4]
  wire [2:0] _GEN_605; // @[Bitwise.scala 48:55:@4058.4]
  wire [3:0] _T_4042; // @[Bitwise.scala 48:55:@4058.4]
  wire [1:0] _T_4043; // @[Bitwise.scala 48:55:@4059.4]
  wire [1:0] _GEN_606; // @[Bitwise.scala 48:55:@4060.4]
  wire [2:0] _T_4044; // @[Bitwise.scala 48:55:@4060.4]
  wire [1:0] _T_4045; // @[Bitwise.scala 48:55:@4061.4]
  wire [1:0] _GEN_607; // @[Bitwise.scala 48:55:@4062.4]
  wire [2:0] _T_4046; // @[Bitwise.scala 48:55:@4062.4]
  wire [3:0] _T_4047; // @[Bitwise.scala 48:55:@4063.4]
  wire [4:0] _T_4048; // @[Bitwise.scala 48:55:@4064.4]
  wire [1:0] _T_4049; // @[Bitwise.scala 48:55:@4065.4]
  wire [1:0] _T_4050; // @[Bitwise.scala 48:55:@4066.4]
  wire [1:0] _GEN_608; // @[Bitwise.scala 48:55:@4067.4]
  wire [2:0] _T_4051; // @[Bitwise.scala 48:55:@4067.4]
  wire [2:0] _GEN_609; // @[Bitwise.scala 48:55:@4068.4]
  wire [3:0] _T_4052; // @[Bitwise.scala 48:55:@4068.4]
  wire [1:0] _T_4053; // @[Bitwise.scala 48:55:@4069.4]
  wire [1:0] _GEN_610; // @[Bitwise.scala 48:55:@4070.4]
  wire [2:0] _T_4054; // @[Bitwise.scala 48:55:@4070.4]
  wire [1:0] _T_4055; // @[Bitwise.scala 48:55:@4071.4]
  wire [1:0] _GEN_611; // @[Bitwise.scala 48:55:@4072.4]
  wire [2:0] _T_4056; // @[Bitwise.scala 48:55:@4072.4]
  wire [3:0] _T_4057; // @[Bitwise.scala 48:55:@4073.4]
  wire [4:0] _T_4058; // @[Bitwise.scala 48:55:@4074.4]
  wire [5:0] _T_4059; // @[Bitwise.scala 48:55:@4075.4]
  wire [22:0] _T_4123; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4140.4]
  wire  _T_4124; // @[Bitwise.scala 50:65:@4141.4]
  wire  _T_4125; // @[Bitwise.scala 50:65:@4142.4]
  wire  _T_4126; // @[Bitwise.scala 50:65:@4143.4]
  wire  _T_4127; // @[Bitwise.scala 50:65:@4144.4]
  wire  _T_4128; // @[Bitwise.scala 50:65:@4145.4]
  wire  _T_4129; // @[Bitwise.scala 50:65:@4146.4]
  wire  _T_4130; // @[Bitwise.scala 50:65:@4147.4]
  wire  _T_4131; // @[Bitwise.scala 50:65:@4148.4]
  wire  _T_4132; // @[Bitwise.scala 50:65:@4149.4]
  wire  _T_4133; // @[Bitwise.scala 50:65:@4150.4]
  wire  _T_4134; // @[Bitwise.scala 50:65:@4151.4]
  wire  _T_4135; // @[Bitwise.scala 50:65:@4152.4]
  wire  _T_4136; // @[Bitwise.scala 50:65:@4153.4]
  wire  _T_4137; // @[Bitwise.scala 50:65:@4154.4]
  wire  _T_4138; // @[Bitwise.scala 50:65:@4155.4]
  wire  _T_4139; // @[Bitwise.scala 50:65:@4156.4]
  wire  _T_4140; // @[Bitwise.scala 50:65:@4157.4]
  wire  _T_4141; // @[Bitwise.scala 50:65:@4158.4]
  wire  _T_4142; // @[Bitwise.scala 50:65:@4159.4]
  wire  _T_4143; // @[Bitwise.scala 50:65:@4160.4]
  wire  _T_4144; // @[Bitwise.scala 50:65:@4161.4]
  wire  _T_4145; // @[Bitwise.scala 50:65:@4162.4]
  wire  _T_4146; // @[Bitwise.scala 50:65:@4163.4]
  wire [1:0] _T_4147; // @[Bitwise.scala 48:55:@4164.4]
  wire [1:0] _T_4148; // @[Bitwise.scala 48:55:@4165.4]
  wire [1:0] _GEN_612; // @[Bitwise.scala 48:55:@4166.4]
  wire [2:0] _T_4149; // @[Bitwise.scala 48:55:@4166.4]
  wire [2:0] _GEN_613; // @[Bitwise.scala 48:55:@4167.4]
  wire [3:0] _T_4150; // @[Bitwise.scala 48:55:@4167.4]
  wire [1:0] _T_4151; // @[Bitwise.scala 48:55:@4168.4]
  wire [1:0] _GEN_614; // @[Bitwise.scala 48:55:@4169.4]
  wire [2:0] _T_4152; // @[Bitwise.scala 48:55:@4169.4]
  wire [1:0] _T_4153; // @[Bitwise.scala 48:55:@4170.4]
  wire [1:0] _GEN_615; // @[Bitwise.scala 48:55:@4171.4]
  wire [2:0] _T_4154; // @[Bitwise.scala 48:55:@4171.4]
  wire [3:0] _T_4155; // @[Bitwise.scala 48:55:@4172.4]
  wire [4:0] _T_4156; // @[Bitwise.scala 48:55:@4173.4]
  wire [1:0] _T_4157; // @[Bitwise.scala 48:55:@4174.4]
  wire [1:0] _GEN_616; // @[Bitwise.scala 48:55:@4175.4]
  wire [2:0] _T_4158; // @[Bitwise.scala 48:55:@4175.4]
  wire [1:0] _T_4159; // @[Bitwise.scala 48:55:@4176.4]
  wire [1:0] _GEN_617; // @[Bitwise.scala 48:55:@4177.4]
  wire [2:0] _T_4160; // @[Bitwise.scala 48:55:@4177.4]
  wire [3:0] _T_4161; // @[Bitwise.scala 48:55:@4178.4]
  wire [1:0] _T_4162; // @[Bitwise.scala 48:55:@4179.4]
  wire [1:0] _GEN_618; // @[Bitwise.scala 48:55:@4180.4]
  wire [2:0] _T_4163; // @[Bitwise.scala 48:55:@4180.4]
  wire [1:0] _T_4164; // @[Bitwise.scala 48:55:@4181.4]
  wire [1:0] _GEN_619; // @[Bitwise.scala 48:55:@4182.4]
  wire [2:0] _T_4165; // @[Bitwise.scala 48:55:@4182.4]
  wire [3:0] _T_4166; // @[Bitwise.scala 48:55:@4183.4]
  wire [4:0] _T_4167; // @[Bitwise.scala 48:55:@4184.4]
  wire [5:0] _T_4168; // @[Bitwise.scala 48:55:@4185.4]
  wire [23:0] _T_4232; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4250.4]
  wire  _T_4233; // @[Bitwise.scala 50:65:@4251.4]
  wire  _T_4234; // @[Bitwise.scala 50:65:@4252.4]
  wire  _T_4235; // @[Bitwise.scala 50:65:@4253.4]
  wire  _T_4236; // @[Bitwise.scala 50:65:@4254.4]
  wire  _T_4237; // @[Bitwise.scala 50:65:@4255.4]
  wire  _T_4238; // @[Bitwise.scala 50:65:@4256.4]
  wire  _T_4239; // @[Bitwise.scala 50:65:@4257.4]
  wire  _T_4240; // @[Bitwise.scala 50:65:@4258.4]
  wire  _T_4241; // @[Bitwise.scala 50:65:@4259.4]
  wire  _T_4242; // @[Bitwise.scala 50:65:@4260.4]
  wire  _T_4243; // @[Bitwise.scala 50:65:@4261.4]
  wire  _T_4244; // @[Bitwise.scala 50:65:@4262.4]
  wire  _T_4245; // @[Bitwise.scala 50:65:@4263.4]
  wire  _T_4246; // @[Bitwise.scala 50:65:@4264.4]
  wire  _T_4247; // @[Bitwise.scala 50:65:@4265.4]
  wire  _T_4248; // @[Bitwise.scala 50:65:@4266.4]
  wire  _T_4249; // @[Bitwise.scala 50:65:@4267.4]
  wire  _T_4250; // @[Bitwise.scala 50:65:@4268.4]
  wire  _T_4251; // @[Bitwise.scala 50:65:@4269.4]
  wire  _T_4252; // @[Bitwise.scala 50:65:@4270.4]
  wire  _T_4253; // @[Bitwise.scala 50:65:@4271.4]
  wire  _T_4254; // @[Bitwise.scala 50:65:@4272.4]
  wire  _T_4255; // @[Bitwise.scala 50:65:@4273.4]
  wire  _T_4256; // @[Bitwise.scala 50:65:@4274.4]
  wire [1:0] _T_4257; // @[Bitwise.scala 48:55:@4275.4]
  wire [1:0] _GEN_620; // @[Bitwise.scala 48:55:@4276.4]
  wire [2:0] _T_4258; // @[Bitwise.scala 48:55:@4276.4]
  wire [1:0] _T_4259; // @[Bitwise.scala 48:55:@4277.4]
  wire [1:0] _GEN_621; // @[Bitwise.scala 48:55:@4278.4]
  wire [2:0] _T_4260; // @[Bitwise.scala 48:55:@4278.4]
  wire [3:0] _T_4261; // @[Bitwise.scala 48:55:@4279.4]
  wire [1:0] _T_4262; // @[Bitwise.scala 48:55:@4280.4]
  wire [1:0] _GEN_622; // @[Bitwise.scala 48:55:@4281.4]
  wire [2:0] _T_4263; // @[Bitwise.scala 48:55:@4281.4]
  wire [1:0] _T_4264; // @[Bitwise.scala 48:55:@4282.4]
  wire [1:0] _GEN_623; // @[Bitwise.scala 48:55:@4283.4]
  wire [2:0] _T_4265; // @[Bitwise.scala 48:55:@4283.4]
  wire [3:0] _T_4266; // @[Bitwise.scala 48:55:@4284.4]
  wire [4:0] _T_4267; // @[Bitwise.scala 48:55:@4285.4]
  wire [1:0] _T_4268; // @[Bitwise.scala 48:55:@4286.4]
  wire [1:0] _GEN_624; // @[Bitwise.scala 48:55:@4287.4]
  wire [2:0] _T_4269; // @[Bitwise.scala 48:55:@4287.4]
  wire [1:0] _T_4270; // @[Bitwise.scala 48:55:@4288.4]
  wire [1:0] _GEN_625; // @[Bitwise.scala 48:55:@4289.4]
  wire [2:0] _T_4271; // @[Bitwise.scala 48:55:@4289.4]
  wire [3:0] _T_4272; // @[Bitwise.scala 48:55:@4290.4]
  wire [1:0] _T_4273; // @[Bitwise.scala 48:55:@4291.4]
  wire [1:0] _GEN_626; // @[Bitwise.scala 48:55:@4292.4]
  wire [2:0] _T_4274; // @[Bitwise.scala 48:55:@4292.4]
  wire [1:0] _T_4275; // @[Bitwise.scala 48:55:@4293.4]
  wire [1:0] _GEN_627; // @[Bitwise.scala 48:55:@4294.4]
  wire [2:0] _T_4276; // @[Bitwise.scala 48:55:@4294.4]
  wire [3:0] _T_4277; // @[Bitwise.scala 48:55:@4295.4]
  wire [4:0] _T_4278; // @[Bitwise.scala 48:55:@4296.4]
  wire [5:0] _T_4279; // @[Bitwise.scala 48:55:@4297.4]
  wire [24:0] _T_4343; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4362.4]
  wire  _T_4344; // @[Bitwise.scala 50:65:@4363.4]
  wire  _T_4345; // @[Bitwise.scala 50:65:@4364.4]
  wire  _T_4346; // @[Bitwise.scala 50:65:@4365.4]
  wire  _T_4347; // @[Bitwise.scala 50:65:@4366.4]
  wire  _T_4348; // @[Bitwise.scala 50:65:@4367.4]
  wire  _T_4349; // @[Bitwise.scala 50:65:@4368.4]
  wire  _T_4350; // @[Bitwise.scala 50:65:@4369.4]
  wire  _T_4351; // @[Bitwise.scala 50:65:@4370.4]
  wire  _T_4352; // @[Bitwise.scala 50:65:@4371.4]
  wire  _T_4353; // @[Bitwise.scala 50:65:@4372.4]
  wire  _T_4354; // @[Bitwise.scala 50:65:@4373.4]
  wire  _T_4355; // @[Bitwise.scala 50:65:@4374.4]
  wire  _T_4356; // @[Bitwise.scala 50:65:@4375.4]
  wire  _T_4357; // @[Bitwise.scala 50:65:@4376.4]
  wire  _T_4358; // @[Bitwise.scala 50:65:@4377.4]
  wire  _T_4359; // @[Bitwise.scala 50:65:@4378.4]
  wire  _T_4360; // @[Bitwise.scala 50:65:@4379.4]
  wire  _T_4361; // @[Bitwise.scala 50:65:@4380.4]
  wire  _T_4362; // @[Bitwise.scala 50:65:@4381.4]
  wire  _T_4363; // @[Bitwise.scala 50:65:@4382.4]
  wire  _T_4364; // @[Bitwise.scala 50:65:@4383.4]
  wire  _T_4365; // @[Bitwise.scala 50:65:@4384.4]
  wire  _T_4366; // @[Bitwise.scala 50:65:@4385.4]
  wire  _T_4367; // @[Bitwise.scala 50:65:@4386.4]
  wire  _T_4368; // @[Bitwise.scala 50:65:@4387.4]
  wire [1:0] _T_4369; // @[Bitwise.scala 48:55:@4388.4]
  wire [1:0] _GEN_628; // @[Bitwise.scala 48:55:@4389.4]
  wire [2:0] _T_4370; // @[Bitwise.scala 48:55:@4389.4]
  wire [1:0] _T_4371; // @[Bitwise.scala 48:55:@4390.4]
  wire [1:0] _GEN_629; // @[Bitwise.scala 48:55:@4391.4]
  wire [2:0] _T_4372; // @[Bitwise.scala 48:55:@4391.4]
  wire [3:0] _T_4373; // @[Bitwise.scala 48:55:@4392.4]
  wire [1:0] _T_4374; // @[Bitwise.scala 48:55:@4393.4]
  wire [1:0] _GEN_630; // @[Bitwise.scala 48:55:@4394.4]
  wire [2:0] _T_4375; // @[Bitwise.scala 48:55:@4394.4]
  wire [1:0] _T_4376; // @[Bitwise.scala 48:55:@4395.4]
  wire [1:0] _GEN_631; // @[Bitwise.scala 48:55:@4396.4]
  wire [2:0] _T_4377; // @[Bitwise.scala 48:55:@4396.4]
  wire [3:0] _T_4378; // @[Bitwise.scala 48:55:@4397.4]
  wire [4:0] _T_4379; // @[Bitwise.scala 48:55:@4398.4]
  wire [1:0] _T_4380; // @[Bitwise.scala 48:55:@4399.4]
  wire [1:0] _GEN_632; // @[Bitwise.scala 48:55:@4400.4]
  wire [2:0] _T_4381; // @[Bitwise.scala 48:55:@4400.4]
  wire [1:0] _T_4382; // @[Bitwise.scala 48:55:@4401.4]
  wire [1:0] _GEN_633; // @[Bitwise.scala 48:55:@4402.4]
  wire [2:0] _T_4383; // @[Bitwise.scala 48:55:@4402.4]
  wire [3:0] _T_4384; // @[Bitwise.scala 48:55:@4403.4]
  wire [1:0] _T_4385; // @[Bitwise.scala 48:55:@4404.4]
  wire [1:0] _GEN_634; // @[Bitwise.scala 48:55:@4405.4]
  wire [2:0] _T_4386; // @[Bitwise.scala 48:55:@4405.4]
  wire [1:0] _T_4387; // @[Bitwise.scala 48:55:@4406.4]
  wire [1:0] _T_4388; // @[Bitwise.scala 48:55:@4407.4]
  wire [2:0] _T_4389; // @[Bitwise.scala 48:55:@4408.4]
  wire [3:0] _T_4390; // @[Bitwise.scala 48:55:@4409.4]
  wire [4:0] _T_4391; // @[Bitwise.scala 48:55:@4410.4]
  wire [5:0] _T_4392; // @[Bitwise.scala 48:55:@4411.4]
  wire [25:0] _T_4456; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4476.4]
  wire  _T_4457; // @[Bitwise.scala 50:65:@4477.4]
  wire  _T_4458; // @[Bitwise.scala 50:65:@4478.4]
  wire  _T_4459; // @[Bitwise.scala 50:65:@4479.4]
  wire  _T_4460; // @[Bitwise.scala 50:65:@4480.4]
  wire  _T_4461; // @[Bitwise.scala 50:65:@4481.4]
  wire  _T_4462; // @[Bitwise.scala 50:65:@4482.4]
  wire  _T_4463; // @[Bitwise.scala 50:65:@4483.4]
  wire  _T_4464; // @[Bitwise.scala 50:65:@4484.4]
  wire  _T_4465; // @[Bitwise.scala 50:65:@4485.4]
  wire  _T_4466; // @[Bitwise.scala 50:65:@4486.4]
  wire  _T_4467; // @[Bitwise.scala 50:65:@4487.4]
  wire  _T_4468; // @[Bitwise.scala 50:65:@4488.4]
  wire  _T_4469; // @[Bitwise.scala 50:65:@4489.4]
  wire  _T_4470; // @[Bitwise.scala 50:65:@4490.4]
  wire  _T_4471; // @[Bitwise.scala 50:65:@4491.4]
  wire  _T_4472; // @[Bitwise.scala 50:65:@4492.4]
  wire  _T_4473; // @[Bitwise.scala 50:65:@4493.4]
  wire  _T_4474; // @[Bitwise.scala 50:65:@4494.4]
  wire  _T_4475; // @[Bitwise.scala 50:65:@4495.4]
  wire  _T_4476; // @[Bitwise.scala 50:65:@4496.4]
  wire  _T_4477; // @[Bitwise.scala 50:65:@4497.4]
  wire  _T_4478; // @[Bitwise.scala 50:65:@4498.4]
  wire  _T_4479; // @[Bitwise.scala 50:65:@4499.4]
  wire  _T_4480; // @[Bitwise.scala 50:65:@4500.4]
  wire  _T_4481; // @[Bitwise.scala 50:65:@4501.4]
  wire  _T_4482; // @[Bitwise.scala 50:65:@4502.4]
  wire [1:0] _T_4483; // @[Bitwise.scala 48:55:@4503.4]
  wire [1:0] _GEN_635; // @[Bitwise.scala 48:55:@4504.4]
  wire [2:0] _T_4484; // @[Bitwise.scala 48:55:@4504.4]
  wire [1:0] _T_4485; // @[Bitwise.scala 48:55:@4505.4]
  wire [1:0] _GEN_636; // @[Bitwise.scala 48:55:@4506.4]
  wire [2:0] _T_4486; // @[Bitwise.scala 48:55:@4506.4]
  wire [3:0] _T_4487; // @[Bitwise.scala 48:55:@4507.4]
  wire [1:0] _T_4488; // @[Bitwise.scala 48:55:@4508.4]
  wire [1:0] _GEN_637; // @[Bitwise.scala 48:55:@4509.4]
  wire [2:0] _T_4489; // @[Bitwise.scala 48:55:@4509.4]
  wire [1:0] _T_4490; // @[Bitwise.scala 48:55:@4510.4]
  wire [1:0] _T_4491; // @[Bitwise.scala 48:55:@4511.4]
  wire [2:0] _T_4492; // @[Bitwise.scala 48:55:@4512.4]
  wire [3:0] _T_4493; // @[Bitwise.scala 48:55:@4513.4]
  wire [4:0] _T_4494; // @[Bitwise.scala 48:55:@4514.4]
  wire [1:0] _T_4495; // @[Bitwise.scala 48:55:@4515.4]
  wire [1:0] _GEN_638; // @[Bitwise.scala 48:55:@4516.4]
  wire [2:0] _T_4496; // @[Bitwise.scala 48:55:@4516.4]
  wire [1:0] _T_4497; // @[Bitwise.scala 48:55:@4517.4]
  wire [1:0] _GEN_639; // @[Bitwise.scala 48:55:@4518.4]
  wire [2:0] _T_4498; // @[Bitwise.scala 48:55:@4518.4]
  wire [3:0] _T_4499; // @[Bitwise.scala 48:55:@4519.4]
  wire [1:0] _T_4500; // @[Bitwise.scala 48:55:@4520.4]
  wire [1:0] _GEN_640; // @[Bitwise.scala 48:55:@4521.4]
  wire [2:0] _T_4501; // @[Bitwise.scala 48:55:@4521.4]
  wire [1:0] _T_4502; // @[Bitwise.scala 48:55:@4522.4]
  wire [1:0] _T_4503; // @[Bitwise.scala 48:55:@4523.4]
  wire [2:0] _T_4504; // @[Bitwise.scala 48:55:@4524.4]
  wire [3:0] _T_4505; // @[Bitwise.scala 48:55:@4525.4]
  wire [4:0] _T_4506; // @[Bitwise.scala 48:55:@4526.4]
  wire [5:0] _T_4507; // @[Bitwise.scala 48:55:@4527.4]
  wire [26:0] _T_4571; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4592.4]
  wire  _T_4572; // @[Bitwise.scala 50:65:@4593.4]
  wire  _T_4573; // @[Bitwise.scala 50:65:@4594.4]
  wire  _T_4574; // @[Bitwise.scala 50:65:@4595.4]
  wire  _T_4575; // @[Bitwise.scala 50:65:@4596.4]
  wire  _T_4576; // @[Bitwise.scala 50:65:@4597.4]
  wire  _T_4577; // @[Bitwise.scala 50:65:@4598.4]
  wire  _T_4578; // @[Bitwise.scala 50:65:@4599.4]
  wire  _T_4579; // @[Bitwise.scala 50:65:@4600.4]
  wire  _T_4580; // @[Bitwise.scala 50:65:@4601.4]
  wire  _T_4581; // @[Bitwise.scala 50:65:@4602.4]
  wire  _T_4582; // @[Bitwise.scala 50:65:@4603.4]
  wire  _T_4583; // @[Bitwise.scala 50:65:@4604.4]
  wire  _T_4584; // @[Bitwise.scala 50:65:@4605.4]
  wire  _T_4585; // @[Bitwise.scala 50:65:@4606.4]
  wire  _T_4586; // @[Bitwise.scala 50:65:@4607.4]
  wire  _T_4587; // @[Bitwise.scala 50:65:@4608.4]
  wire  _T_4588; // @[Bitwise.scala 50:65:@4609.4]
  wire  _T_4589; // @[Bitwise.scala 50:65:@4610.4]
  wire  _T_4590; // @[Bitwise.scala 50:65:@4611.4]
  wire  _T_4591; // @[Bitwise.scala 50:65:@4612.4]
  wire  _T_4592; // @[Bitwise.scala 50:65:@4613.4]
  wire  _T_4593; // @[Bitwise.scala 50:65:@4614.4]
  wire  _T_4594; // @[Bitwise.scala 50:65:@4615.4]
  wire  _T_4595; // @[Bitwise.scala 50:65:@4616.4]
  wire  _T_4596; // @[Bitwise.scala 50:65:@4617.4]
  wire  _T_4597; // @[Bitwise.scala 50:65:@4618.4]
  wire  _T_4598; // @[Bitwise.scala 50:65:@4619.4]
  wire [1:0] _T_4599; // @[Bitwise.scala 48:55:@4620.4]
  wire [1:0] _GEN_641; // @[Bitwise.scala 48:55:@4621.4]
  wire [2:0] _T_4600; // @[Bitwise.scala 48:55:@4621.4]
  wire [1:0] _T_4601; // @[Bitwise.scala 48:55:@4622.4]
  wire [1:0] _GEN_642; // @[Bitwise.scala 48:55:@4623.4]
  wire [2:0] _T_4602; // @[Bitwise.scala 48:55:@4623.4]
  wire [3:0] _T_4603; // @[Bitwise.scala 48:55:@4624.4]
  wire [1:0] _T_4604; // @[Bitwise.scala 48:55:@4625.4]
  wire [1:0] _GEN_643; // @[Bitwise.scala 48:55:@4626.4]
  wire [2:0] _T_4605; // @[Bitwise.scala 48:55:@4626.4]
  wire [1:0] _T_4606; // @[Bitwise.scala 48:55:@4627.4]
  wire [1:0] _T_4607; // @[Bitwise.scala 48:55:@4628.4]
  wire [2:0] _T_4608; // @[Bitwise.scala 48:55:@4629.4]
  wire [3:0] _T_4609; // @[Bitwise.scala 48:55:@4630.4]
  wire [4:0] _T_4610; // @[Bitwise.scala 48:55:@4631.4]
  wire [1:0] _T_4611; // @[Bitwise.scala 48:55:@4632.4]
  wire [1:0] _GEN_644; // @[Bitwise.scala 48:55:@4633.4]
  wire [2:0] _T_4612; // @[Bitwise.scala 48:55:@4633.4]
  wire [1:0] _T_4613; // @[Bitwise.scala 48:55:@4634.4]
  wire [1:0] _T_4614; // @[Bitwise.scala 48:55:@4635.4]
  wire [2:0] _T_4615; // @[Bitwise.scala 48:55:@4636.4]
  wire [3:0] _T_4616; // @[Bitwise.scala 48:55:@4637.4]
  wire [1:0] _T_4617; // @[Bitwise.scala 48:55:@4638.4]
  wire [1:0] _GEN_645; // @[Bitwise.scala 48:55:@4639.4]
  wire [2:0] _T_4618; // @[Bitwise.scala 48:55:@4639.4]
  wire [1:0] _T_4619; // @[Bitwise.scala 48:55:@4640.4]
  wire [1:0] _T_4620; // @[Bitwise.scala 48:55:@4641.4]
  wire [2:0] _T_4621; // @[Bitwise.scala 48:55:@4642.4]
  wire [3:0] _T_4622; // @[Bitwise.scala 48:55:@4643.4]
  wire [4:0] _T_4623; // @[Bitwise.scala 48:55:@4644.4]
  wire [5:0] _T_4624; // @[Bitwise.scala 48:55:@4645.4]
  wire [27:0] _T_4688; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4710.4]
  wire  _T_4689; // @[Bitwise.scala 50:65:@4711.4]
  wire  _T_4690; // @[Bitwise.scala 50:65:@4712.4]
  wire  _T_4691; // @[Bitwise.scala 50:65:@4713.4]
  wire  _T_4692; // @[Bitwise.scala 50:65:@4714.4]
  wire  _T_4693; // @[Bitwise.scala 50:65:@4715.4]
  wire  _T_4694; // @[Bitwise.scala 50:65:@4716.4]
  wire  _T_4695; // @[Bitwise.scala 50:65:@4717.4]
  wire  _T_4696; // @[Bitwise.scala 50:65:@4718.4]
  wire  _T_4697; // @[Bitwise.scala 50:65:@4719.4]
  wire  _T_4698; // @[Bitwise.scala 50:65:@4720.4]
  wire  _T_4699; // @[Bitwise.scala 50:65:@4721.4]
  wire  _T_4700; // @[Bitwise.scala 50:65:@4722.4]
  wire  _T_4701; // @[Bitwise.scala 50:65:@4723.4]
  wire  _T_4702; // @[Bitwise.scala 50:65:@4724.4]
  wire  _T_4703; // @[Bitwise.scala 50:65:@4725.4]
  wire  _T_4704; // @[Bitwise.scala 50:65:@4726.4]
  wire  _T_4705; // @[Bitwise.scala 50:65:@4727.4]
  wire  _T_4706; // @[Bitwise.scala 50:65:@4728.4]
  wire  _T_4707; // @[Bitwise.scala 50:65:@4729.4]
  wire  _T_4708; // @[Bitwise.scala 50:65:@4730.4]
  wire  _T_4709; // @[Bitwise.scala 50:65:@4731.4]
  wire  _T_4710; // @[Bitwise.scala 50:65:@4732.4]
  wire  _T_4711; // @[Bitwise.scala 50:65:@4733.4]
  wire  _T_4712; // @[Bitwise.scala 50:65:@4734.4]
  wire  _T_4713; // @[Bitwise.scala 50:65:@4735.4]
  wire  _T_4714; // @[Bitwise.scala 50:65:@4736.4]
  wire  _T_4715; // @[Bitwise.scala 50:65:@4737.4]
  wire  _T_4716; // @[Bitwise.scala 50:65:@4738.4]
  wire [1:0] _T_4717; // @[Bitwise.scala 48:55:@4739.4]
  wire [1:0] _GEN_646; // @[Bitwise.scala 48:55:@4740.4]
  wire [2:0] _T_4718; // @[Bitwise.scala 48:55:@4740.4]
  wire [1:0] _T_4719; // @[Bitwise.scala 48:55:@4741.4]
  wire [1:0] _T_4720; // @[Bitwise.scala 48:55:@4742.4]
  wire [2:0] _T_4721; // @[Bitwise.scala 48:55:@4743.4]
  wire [3:0] _T_4722; // @[Bitwise.scala 48:55:@4744.4]
  wire [1:0] _T_4723; // @[Bitwise.scala 48:55:@4745.4]
  wire [1:0] _GEN_647; // @[Bitwise.scala 48:55:@4746.4]
  wire [2:0] _T_4724; // @[Bitwise.scala 48:55:@4746.4]
  wire [1:0] _T_4725; // @[Bitwise.scala 48:55:@4747.4]
  wire [1:0] _T_4726; // @[Bitwise.scala 48:55:@4748.4]
  wire [2:0] _T_4727; // @[Bitwise.scala 48:55:@4749.4]
  wire [3:0] _T_4728; // @[Bitwise.scala 48:55:@4750.4]
  wire [4:0] _T_4729; // @[Bitwise.scala 48:55:@4751.4]
  wire [1:0] _T_4730; // @[Bitwise.scala 48:55:@4752.4]
  wire [1:0] _GEN_648; // @[Bitwise.scala 48:55:@4753.4]
  wire [2:0] _T_4731; // @[Bitwise.scala 48:55:@4753.4]
  wire [1:0] _T_4732; // @[Bitwise.scala 48:55:@4754.4]
  wire [1:0] _T_4733; // @[Bitwise.scala 48:55:@4755.4]
  wire [2:0] _T_4734; // @[Bitwise.scala 48:55:@4756.4]
  wire [3:0] _T_4735; // @[Bitwise.scala 48:55:@4757.4]
  wire [1:0] _T_4736; // @[Bitwise.scala 48:55:@4758.4]
  wire [1:0] _GEN_649; // @[Bitwise.scala 48:55:@4759.4]
  wire [2:0] _T_4737; // @[Bitwise.scala 48:55:@4759.4]
  wire [1:0] _T_4738; // @[Bitwise.scala 48:55:@4760.4]
  wire [1:0] _T_4739; // @[Bitwise.scala 48:55:@4761.4]
  wire [2:0] _T_4740; // @[Bitwise.scala 48:55:@4762.4]
  wire [3:0] _T_4741; // @[Bitwise.scala 48:55:@4763.4]
  wire [4:0] _T_4742; // @[Bitwise.scala 48:55:@4764.4]
  wire [5:0] _T_4743; // @[Bitwise.scala 48:55:@4765.4]
  wire [28:0] _T_4807; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4830.4]
  wire  _T_4808; // @[Bitwise.scala 50:65:@4831.4]
  wire  _T_4809; // @[Bitwise.scala 50:65:@4832.4]
  wire  _T_4810; // @[Bitwise.scala 50:65:@4833.4]
  wire  _T_4811; // @[Bitwise.scala 50:65:@4834.4]
  wire  _T_4812; // @[Bitwise.scala 50:65:@4835.4]
  wire  _T_4813; // @[Bitwise.scala 50:65:@4836.4]
  wire  _T_4814; // @[Bitwise.scala 50:65:@4837.4]
  wire  _T_4815; // @[Bitwise.scala 50:65:@4838.4]
  wire  _T_4816; // @[Bitwise.scala 50:65:@4839.4]
  wire  _T_4817; // @[Bitwise.scala 50:65:@4840.4]
  wire  _T_4818; // @[Bitwise.scala 50:65:@4841.4]
  wire  _T_4819; // @[Bitwise.scala 50:65:@4842.4]
  wire  _T_4820; // @[Bitwise.scala 50:65:@4843.4]
  wire  _T_4821; // @[Bitwise.scala 50:65:@4844.4]
  wire  _T_4822; // @[Bitwise.scala 50:65:@4845.4]
  wire  _T_4823; // @[Bitwise.scala 50:65:@4846.4]
  wire  _T_4824; // @[Bitwise.scala 50:65:@4847.4]
  wire  _T_4825; // @[Bitwise.scala 50:65:@4848.4]
  wire  _T_4826; // @[Bitwise.scala 50:65:@4849.4]
  wire  _T_4827; // @[Bitwise.scala 50:65:@4850.4]
  wire  _T_4828; // @[Bitwise.scala 50:65:@4851.4]
  wire  _T_4829; // @[Bitwise.scala 50:65:@4852.4]
  wire  _T_4830; // @[Bitwise.scala 50:65:@4853.4]
  wire  _T_4831; // @[Bitwise.scala 50:65:@4854.4]
  wire  _T_4832; // @[Bitwise.scala 50:65:@4855.4]
  wire  _T_4833; // @[Bitwise.scala 50:65:@4856.4]
  wire  _T_4834; // @[Bitwise.scala 50:65:@4857.4]
  wire  _T_4835; // @[Bitwise.scala 50:65:@4858.4]
  wire  _T_4836; // @[Bitwise.scala 50:65:@4859.4]
  wire [1:0] _T_4837; // @[Bitwise.scala 48:55:@4860.4]
  wire [1:0] _GEN_650; // @[Bitwise.scala 48:55:@4861.4]
  wire [2:0] _T_4838; // @[Bitwise.scala 48:55:@4861.4]
  wire [1:0] _T_4839; // @[Bitwise.scala 48:55:@4862.4]
  wire [1:0] _T_4840; // @[Bitwise.scala 48:55:@4863.4]
  wire [2:0] _T_4841; // @[Bitwise.scala 48:55:@4864.4]
  wire [3:0] _T_4842; // @[Bitwise.scala 48:55:@4865.4]
  wire [1:0] _T_4843; // @[Bitwise.scala 48:55:@4866.4]
  wire [1:0] _GEN_651; // @[Bitwise.scala 48:55:@4867.4]
  wire [2:0] _T_4844; // @[Bitwise.scala 48:55:@4867.4]
  wire [1:0] _T_4845; // @[Bitwise.scala 48:55:@4868.4]
  wire [1:0] _T_4846; // @[Bitwise.scala 48:55:@4869.4]
  wire [2:0] _T_4847; // @[Bitwise.scala 48:55:@4870.4]
  wire [3:0] _T_4848; // @[Bitwise.scala 48:55:@4871.4]
  wire [4:0] _T_4849; // @[Bitwise.scala 48:55:@4872.4]
  wire [1:0] _T_4850; // @[Bitwise.scala 48:55:@4873.4]
  wire [1:0] _GEN_652; // @[Bitwise.scala 48:55:@4874.4]
  wire [2:0] _T_4851; // @[Bitwise.scala 48:55:@4874.4]
  wire [1:0] _T_4852; // @[Bitwise.scala 48:55:@4875.4]
  wire [1:0] _T_4853; // @[Bitwise.scala 48:55:@4876.4]
  wire [2:0] _T_4854; // @[Bitwise.scala 48:55:@4877.4]
  wire [3:0] _T_4855; // @[Bitwise.scala 48:55:@4878.4]
  wire [1:0] _T_4856; // @[Bitwise.scala 48:55:@4879.4]
  wire [1:0] _T_4857; // @[Bitwise.scala 48:55:@4880.4]
  wire [2:0] _T_4858; // @[Bitwise.scala 48:55:@4881.4]
  wire [1:0] _T_4859; // @[Bitwise.scala 48:55:@4882.4]
  wire [1:0] _T_4860; // @[Bitwise.scala 48:55:@4883.4]
  wire [2:0] _T_4861; // @[Bitwise.scala 48:55:@4884.4]
  wire [3:0] _T_4862; // @[Bitwise.scala 48:55:@4885.4]
  wire [4:0] _T_4863; // @[Bitwise.scala 48:55:@4886.4]
  wire [5:0] _T_4864; // @[Bitwise.scala 48:55:@4887.4]
  wire [29:0] _T_4928; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4952.4]
  wire  _T_4929; // @[Bitwise.scala 50:65:@4953.4]
  wire  _T_4930; // @[Bitwise.scala 50:65:@4954.4]
  wire  _T_4931; // @[Bitwise.scala 50:65:@4955.4]
  wire  _T_4932; // @[Bitwise.scala 50:65:@4956.4]
  wire  _T_4933; // @[Bitwise.scala 50:65:@4957.4]
  wire  _T_4934; // @[Bitwise.scala 50:65:@4958.4]
  wire  _T_4935; // @[Bitwise.scala 50:65:@4959.4]
  wire  _T_4936; // @[Bitwise.scala 50:65:@4960.4]
  wire  _T_4937; // @[Bitwise.scala 50:65:@4961.4]
  wire  _T_4938; // @[Bitwise.scala 50:65:@4962.4]
  wire  _T_4939; // @[Bitwise.scala 50:65:@4963.4]
  wire  _T_4940; // @[Bitwise.scala 50:65:@4964.4]
  wire  _T_4941; // @[Bitwise.scala 50:65:@4965.4]
  wire  _T_4942; // @[Bitwise.scala 50:65:@4966.4]
  wire  _T_4943; // @[Bitwise.scala 50:65:@4967.4]
  wire  _T_4944; // @[Bitwise.scala 50:65:@4968.4]
  wire  _T_4945; // @[Bitwise.scala 50:65:@4969.4]
  wire  _T_4946; // @[Bitwise.scala 50:65:@4970.4]
  wire  _T_4947; // @[Bitwise.scala 50:65:@4971.4]
  wire  _T_4948; // @[Bitwise.scala 50:65:@4972.4]
  wire  _T_4949; // @[Bitwise.scala 50:65:@4973.4]
  wire  _T_4950; // @[Bitwise.scala 50:65:@4974.4]
  wire  _T_4951; // @[Bitwise.scala 50:65:@4975.4]
  wire  _T_4952; // @[Bitwise.scala 50:65:@4976.4]
  wire  _T_4953; // @[Bitwise.scala 50:65:@4977.4]
  wire  _T_4954; // @[Bitwise.scala 50:65:@4978.4]
  wire  _T_4955; // @[Bitwise.scala 50:65:@4979.4]
  wire  _T_4956; // @[Bitwise.scala 50:65:@4980.4]
  wire  _T_4957; // @[Bitwise.scala 50:65:@4981.4]
  wire  _T_4958; // @[Bitwise.scala 50:65:@4982.4]
  wire [1:0] _T_4959; // @[Bitwise.scala 48:55:@4983.4]
  wire [1:0] _GEN_653; // @[Bitwise.scala 48:55:@4984.4]
  wire [2:0] _T_4960; // @[Bitwise.scala 48:55:@4984.4]
  wire [1:0] _T_4961; // @[Bitwise.scala 48:55:@4985.4]
  wire [1:0] _T_4962; // @[Bitwise.scala 48:55:@4986.4]
  wire [2:0] _T_4963; // @[Bitwise.scala 48:55:@4987.4]
  wire [3:0] _T_4964; // @[Bitwise.scala 48:55:@4988.4]
  wire [1:0] _T_4965; // @[Bitwise.scala 48:55:@4989.4]
  wire [1:0] _T_4966; // @[Bitwise.scala 48:55:@4990.4]
  wire [2:0] _T_4967; // @[Bitwise.scala 48:55:@4991.4]
  wire [1:0] _T_4968; // @[Bitwise.scala 48:55:@4992.4]
  wire [1:0] _T_4969; // @[Bitwise.scala 48:55:@4993.4]
  wire [2:0] _T_4970; // @[Bitwise.scala 48:55:@4994.4]
  wire [3:0] _T_4971; // @[Bitwise.scala 48:55:@4995.4]
  wire [4:0] _T_4972; // @[Bitwise.scala 48:55:@4996.4]
  wire [1:0] _T_4973; // @[Bitwise.scala 48:55:@4997.4]
  wire [1:0] _GEN_654; // @[Bitwise.scala 48:55:@4998.4]
  wire [2:0] _T_4974; // @[Bitwise.scala 48:55:@4998.4]
  wire [1:0] _T_4975; // @[Bitwise.scala 48:55:@4999.4]
  wire [1:0] _T_4976; // @[Bitwise.scala 48:55:@5000.4]
  wire [2:0] _T_4977; // @[Bitwise.scala 48:55:@5001.4]
  wire [3:0] _T_4978; // @[Bitwise.scala 48:55:@5002.4]
  wire [1:0] _T_4979; // @[Bitwise.scala 48:55:@5003.4]
  wire [1:0] _T_4980; // @[Bitwise.scala 48:55:@5004.4]
  wire [2:0] _T_4981; // @[Bitwise.scala 48:55:@5005.4]
  wire [1:0] _T_4982; // @[Bitwise.scala 48:55:@5006.4]
  wire [1:0] _T_4983; // @[Bitwise.scala 48:55:@5007.4]
  wire [2:0] _T_4984; // @[Bitwise.scala 48:55:@5008.4]
  wire [3:0] _T_4985; // @[Bitwise.scala 48:55:@5009.4]
  wire [4:0] _T_4986; // @[Bitwise.scala 48:55:@5010.4]
  wire [5:0] _T_4987; // @[Bitwise.scala 48:55:@5011.4]
  wire [30:0] _T_5051; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5076.4]
  wire  _T_5052; // @[Bitwise.scala 50:65:@5077.4]
  wire  _T_5053; // @[Bitwise.scala 50:65:@5078.4]
  wire  _T_5054; // @[Bitwise.scala 50:65:@5079.4]
  wire  _T_5055; // @[Bitwise.scala 50:65:@5080.4]
  wire  _T_5056; // @[Bitwise.scala 50:65:@5081.4]
  wire  _T_5057; // @[Bitwise.scala 50:65:@5082.4]
  wire  _T_5058; // @[Bitwise.scala 50:65:@5083.4]
  wire  _T_5059; // @[Bitwise.scala 50:65:@5084.4]
  wire  _T_5060; // @[Bitwise.scala 50:65:@5085.4]
  wire  _T_5061; // @[Bitwise.scala 50:65:@5086.4]
  wire  _T_5062; // @[Bitwise.scala 50:65:@5087.4]
  wire  _T_5063; // @[Bitwise.scala 50:65:@5088.4]
  wire  _T_5064; // @[Bitwise.scala 50:65:@5089.4]
  wire  _T_5065; // @[Bitwise.scala 50:65:@5090.4]
  wire  _T_5066; // @[Bitwise.scala 50:65:@5091.4]
  wire  _T_5067; // @[Bitwise.scala 50:65:@5092.4]
  wire  _T_5068; // @[Bitwise.scala 50:65:@5093.4]
  wire  _T_5069; // @[Bitwise.scala 50:65:@5094.4]
  wire  _T_5070; // @[Bitwise.scala 50:65:@5095.4]
  wire  _T_5071; // @[Bitwise.scala 50:65:@5096.4]
  wire  _T_5072; // @[Bitwise.scala 50:65:@5097.4]
  wire  _T_5073; // @[Bitwise.scala 50:65:@5098.4]
  wire  _T_5074; // @[Bitwise.scala 50:65:@5099.4]
  wire  _T_5075; // @[Bitwise.scala 50:65:@5100.4]
  wire  _T_5076; // @[Bitwise.scala 50:65:@5101.4]
  wire  _T_5077; // @[Bitwise.scala 50:65:@5102.4]
  wire  _T_5078; // @[Bitwise.scala 50:65:@5103.4]
  wire  _T_5079; // @[Bitwise.scala 50:65:@5104.4]
  wire  _T_5080; // @[Bitwise.scala 50:65:@5105.4]
  wire  _T_5081; // @[Bitwise.scala 50:65:@5106.4]
  wire  _T_5082; // @[Bitwise.scala 50:65:@5107.4]
  wire [1:0] _T_5083; // @[Bitwise.scala 48:55:@5108.4]
  wire [1:0] _GEN_655; // @[Bitwise.scala 48:55:@5109.4]
  wire [2:0] _T_5084; // @[Bitwise.scala 48:55:@5109.4]
  wire [1:0] _T_5085; // @[Bitwise.scala 48:55:@5110.4]
  wire [1:0] _T_5086; // @[Bitwise.scala 48:55:@5111.4]
  wire [2:0] _T_5087; // @[Bitwise.scala 48:55:@5112.4]
  wire [3:0] _T_5088; // @[Bitwise.scala 48:55:@5113.4]
  wire [1:0] _T_5089; // @[Bitwise.scala 48:55:@5114.4]
  wire [1:0] _T_5090; // @[Bitwise.scala 48:55:@5115.4]
  wire [2:0] _T_5091; // @[Bitwise.scala 48:55:@5116.4]
  wire [1:0] _T_5092; // @[Bitwise.scala 48:55:@5117.4]
  wire [1:0] _T_5093; // @[Bitwise.scala 48:55:@5118.4]
  wire [2:0] _T_5094; // @[Bitwise.scala 48:55:@5119.4]
  wire [3:0] _T_5095; // @[Bitwise.scala 48:55:@5120.4]
  wire [4:0] _T_5096; // @[Bitwise.scala 48:55:@5121.4]
  wire [1:0] _T_5097; // @[Bitwise.scala 48:55:@5122.4]
  wire [1:0] _T_5098; // @[Bitwise.scala 48:55:@5123.4]
  wire [2:0] _T_5099; // @[Bitwise.scala 48:55:@5124.4]
  wire [1:0] _T_5100; // @[Bitwise.scala 48:55:@5125.4]
  wire [1:0] _T_5101; // @[Bitwise.scala 48:55:@5126.4]
  wire [2:0] _T_5102; // @[Bitwise.scala 48:55:@5127.4]
  wire [3:0] _T_5103; // @[Bitwise.scala 48:55:@5128.4]
  wire [1:0] _T_5104; // @[Bitwise.scala 48:55:@5129.4]
  wire [1:0] _T_5105; // @[Bitwise.scala 48:55:@5130.4]
  wire [2:0] _T_5106; // @[Bitwise.scala 48:55:@5131.4]
  wire [1:0] _T_5107; // @[Bitwise.scala 48:55:@5132.4]
  wire [1:0] _T_5108; // @[Bitwise.scala 48:55:@5133.4]
  wire [2:0] _T_5109; // @[Bitwise.scala 48:55:@5134.4]
  wire [3:0] _T_5110; // @[Bitwise.scala 48:55:@5135.4]
  wire [4:0] _T_5111; // @[Bitwise.scala 48:55:@5136.4]
  wire [5:0] _T_5112; // @[Bitwise.scala 48:55:@5137.4]
  wire [31:0] _T_5176; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5202.4]
  wire  _T_5177; // @[Bitwise.scala 50:65:@5203.4]
  wire  _T_5178; // @[Bitwise.scala 50:65:@5204.4]
  wire  _T_5179; // @[Bitwise.scala 50:65:@5205.4]
  wire  _T_5180; // @[Bitwise.scala 50:65:@5206.4]
  wire  _T_5181; // @[Bitwise.scala 50:65:@5207.4]
  wire  _T_5182; // @[Bitwise.scala 50:65:@5208.4]
  wire  _T_5183; // @[Bitwise.scala 50:65:@5209.4]
  wire  _T_5184; // @[Bitwise.scala 50:65:@5210.4]
  wire  _T_5185; // @[Bitwise.scala 50:65:@5211.4]
  wire  _T_5186; // @[Bitwise.scala 50:65:@5212.4]
  wire  _T_5187; // @[Bitwise.scala 50:65:@5213.4]
  wire  _T_5188; // @[Bitwise.scala 50:65:@5214.4]
  wire  _T_5189; // @[Bitwise.scala 50:65:@5215.4]
  wire  _T_5190; // @[Bitwise.scala 50:65:@5216.4]
  wire  _T_5191; // @[Bitwise.scala 50:65:@5217.4]
  wire  _T_5192; // @[Bitwise.scala 50:65:@5218.4]
  wire  _T_5193; // @[Bitwise.scala 50:65:@5219.4]
  wire  _T_5194; // @[Bitwise.scala 50:65:@5220.4]
  wire  _T_5195; // @[Bitwise.scala 50:65:@5221.4]
  wire  _T_5196; // @[Bitwise.scala 50:65:@5222.4]
  wire  _T_5197; // @[Bitwise.scala 50:65:@5223.4]
  wire  _T_5198; // @[Bitwise.scala 50:65:@5224.4]
  wire  _T_5199; // @[Bitwise.scala 50:65:@5225.4]
  wire  _T_5200; // @[Bitwise.scala 50:65:@5226.4]
  wire  _T_5201; // @[Bitwise.scala 50:65:@5227.4]
  wire  _T_5202; // @[Bitwise.scala 50:65:@5228.4]
  wire  _T_5203; // @[Bitwise.scala 50:65:@5229.4]
  wire  _T_5204; // @[Bitwise.scala 50:65:@5230.4]
  wire  _T_5205; // @[Bitwise.scala 50:65:@5231.4]
  wire  _T_5206; // @[Bitwise.scala 50:65:@5232.4]
  wire  _T_5207; // @[Bitwise.scala 50:65:@5233.4]
  wire  _T_5208; // @[Bitwise.scala 50:65:@5234.4]
  wire [1:0] _T_5209; // @[Bitwise.scala 48:55:@5235.4]
  wire [1:0] _T_5210; // @[Bitwise.scala 48:55:@5236.4]
  wire [2:0] _T_5211; // @[Bitwise.scala 48:55:@5237.4]
  wire [1:0] _T_5212; // @[Bitwise.scala 48:55:@5238.4]
  wire [1:0] _T_5213; // @[Bitwise.scala 48:55:@5239.4]
  wire [2:0] _T_5214; // @[Bitwise.scala 48:55:@5240.4]
  wire [3:0] _T_5215; // @[Bitwise.scala 48:55:@5241.4]
  wire [1:0] _T_5216; // @[Bitwise.scala 48:55:@5242.4]
  wire [1:0] _T_5217; // @[Bitwise.scala 48:55:@5243.4]
  wire [2:0] _T_5218; // @[Bitwise.scala 48:55:@5244.4]
  wire [1:0] _T_5219; // @[Bitwise.scala 48:55:@5245.4]
  wire [1:0] _T_5220; // @[Bitwise.scala 48:55:@5246.4]
  wire [2:0] _T_5221; // @[Bitwise.scala 48:55:@5247.4]
  wire [3:0] _T_5222; // @[Bitwise.scala 48:55:@5248.4]
  wire [4:0] _T_5223; // @[Bitwise.scala 48:55:@5249.4]
  wire [1:0] _T_5224; // @[Bitwise.scala 48:55:@5250.4]
  wire [1:0] _T_5225; // @[Bitwise.scala 48:55:@5251.4]
  wire [2:0] _T_5226; // @[Bitwise.scala 48:55:@5252.4]
  wire [1:0] _T_5227; // @[Bitwise.scala 48:55:@5253.4]
  wire [1:0] _T_5228; // @[Bitwise.scala 48:55:@5254.4]
  wire [2:0] _T_5229; // @[Bitwise.scala 48:55:@5255.4]
  wire [3:0] _T_5230; // @[Bitwise.scala 48:55:@5256.4]
  wire [1:0] _T_5231; // @[Bitwise.scala 48:55:@5257.4]
  wire [1:0] _T_5232; // @[Bitwise.scala 48:55:@5258.4]
  wire [2:0] _T_5233; // @[Bitwise.scala 48:55:@5259.4]
  wire [1:0] _T_5234; // @[Bitwise.scala 48:55:@5260.4]
  wire [1:0] _T_5235; // @[Bitwise.scala 48:55:@5261.4]
  wire [2:0] _T_5236; // @[Bitwise.scala 48:55:@5262.4]
  wire [3:0] _T_5237; // @[Bitwise.scala 48:55:@5263.4]
  wire [4:0] _T_5238; // @[Bitwise.scala 48:55:@5264.4]
  wire [5:0] _T_5239; // @[Bitwise.scala 48:55:@5265.4]
  wire [32:0] _T_5303; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5330.4]
  wire  _T_5304; // @[Bitwise.scala 50:65:@5331.4]
  wire  _T_5305; // @[Bitwise.scala 50:65:@5332.4]
  wire  _T_5306; // @[Bitwise.scala 50:65:@5333.4]
  wire  _T_5307; // @[Bitwise.scala 50:65:@5334.4]
  wire  _T_5308; // @[Bitwise.scala 50:65:@5335.4]
  wire  _T_5309; // @[Bitwise.scala 50:65:@5336.4]
  wire  _T_5310; // @[Bitwise.scala 50:65:@5337.4]
  wire  _T_5311; // @[Bitwise.scala 50:65:@5338.4]
  wire  _T_5312; // @[Bitwise.scala 50:65:@5339.4]
  wire  _T_5313; // @[Bitwise.scala 50:65:@5340.4]
  wire  _T_5314; // @[Bitwise.scala 50:65:@5341.4]
  wire  _T_5315; // @[Bitwise.scala 50:65:@5342.4]
  wire  _T_5316; // @[Bitwise.scala 50:65:@5343.4]
  wire  _T_5317; // @[Bitwise.scala 50:65:@5344.4]
  wire  _T_5318; // @[Bitwise.scala 50:65:@5345.4]
  wire  _T_5319; // @[Bitwise.scala 50:65:@5346.4]
  wire  _T_5320; // @[Bitwise.scala 50:65:@5347.4]
  wire  _T_5321; // @[Bitwise.scala 50:65:@5348.4]
  wire  _T_5322; // @[Bitwise.scala 50:65:@5349.4]
  wire  _T_5323; // @[Bitwise.scala 50:65:@5350.4]
  wire  _T_5324; // @[Bitwise.scala 50:65:@5351.4]
  wire  _T_5325; // @[Bitwise.scala 50:65:@5352.4]
  wire  _T_5326; // @[Bitwise.scala 50:65:@5353.4]
  wire  _T_5327; // @[Bitwise.scala 50:65:@5354.4]
  wire  _T_5328; // @[Bitwise.scala 50:65:@5355.4]
  wire  _T_5329; // @[Bitwise.scala 50:65:@5356.4]
  wire  _T_5330; // @[Bitwise.scala 50:65:@5357.4]
  wire  _T_5331; // @[Bitwise.scala 50:65:@5358.4]
  wire  _T_5332; // @[Bitwise.scala 50:65:@5359.4]
  wire  _T_5333; // @[Bitwise.scala 50:65:@5360.4]
  wire  _T_5334; // @[Bitwise.scala 50:65:@5361.4]
  wire  _T_5335; // @[Bitwise.scala 50:65:@5362.4]
  wire  _T_5336; // @[Bitwise.scala 50:65:@5363.4]
  wire [1:0] _T_5337; // @[Bitwise.scala 48:55:@5364.4]
  wire [1:0] _T_5338; // @[Bitwise.scala 48:55:@5365.4]
  wire [2:0] _T_5339; // @[Bitwise.scala 48:55:@5366.4]
  wire [1:0] _T_5340; // @[Bitwise.scala 48:55:@5367.4]
  wire [1:0] _T_5341; // @[Bitwise.scala 48:55:@5368.4]
  wire [2:0] _T_5342; // @[Bitwise.scala 48:55:@5369.4]
  wire [3:0] _T_5343; // @[Bitwise.scala 48:55:@5370.4]
  wire [1:0] _T_5344; // @[Bitwise.scala 48:55:@5371.4]
  wire [1:0] _T_5345; // @[Bitwise.scala 48:55:@5372.4]
  wire [2:0] _T_5346; // @[Bitwise.scala 48:55:@5373.4]
  wire [1:0] _T_5347; // @[Bitwise.scala 48:55:@5374.4]
  wire [1:0] _T_5348; // @[Bitwise.scala 48:55:@5375.4]
  wire [2:0] _T_5349; // @[Bitwise.scala 48:55:@5376.4]
  wire [3:0] _T_5350; // @[Bitwise.scala 48:55:@5377.4]
  wire [4:0] _T_5351; // @[Bitwise.scala 48:55:@5378.4]
  wire [1:0] _T_5352; // @[Bitwise.scala 48:55:@5379.4]
  wire [1:0] _T_5353; // @[Bitwise.scala 48:55:@5380.4]
  wire [2:0] _T_5354; // @[Bitwise.scala 48:55:@5381.4]
  wire [1:0] _T_5355; // @[Bitwise.scala 48:55:@5382.4]
  wire [1:0] _T_5356; // @[Bitwise.scala 48:55:@5383.4]
  wire [2:0] _T_5357; // @[Bitwise.scala 48:55:@5384.4]
  wire [3:0] _T_5358; // @[Bitwise.scala 48:55:@5385.4]
  wire [1:0] _T_5359; // @[Bitwise.scala 48:55:@5386.4]
  wire [1:0] _T_5360; // @[Bitwise.scala 48:55:@5387.4]
  wire [2:0] _T_5361; // @[Bitwise.scala 48:55:@5388.4]
  wire [1:0] _T_5362; // @[Bitwise.scala 48:55:@5389.4]
  wire [1:0] _T_5363; // @[Bitwise.scala 48:55:@5390.4]
  wire [1:0] _GEN_656; // @[Bitwise.scala 48:55:@5391.4]
  wire [2:0] _T_5364; // @[Bitwise.scala 48:55:@5391.4]
  wire [2:0] _GEN_657; // @[Bitwise.scala 48:55:@5392.4]
  wire [3:0] _T_5365; // @[Bitwise.scala 48:55:@5392.4]
  wire [3:0] _GEN_658; // @[Bitwise.scala 48:55:@5393.4]
  wire [4:0] _T_5366; // @[Bitwise.scala 48:55:@5393.4]
  wire [4:0] _GEN_659; // @[Bitwise.scala 48:55:@5394.4]
  wire [5:0] _T_5367; // @[Bitwise.scala 48:55:@5394.4]
  wire [5:0] _GEN_660; // @[Bitwise.scala 48:55:@5395.4]
  wire [6:0] _T_5368; // @[Bitwise.scala 48:55:@5395.4]
  wire [33:0] _T_5432; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5460.4]
  wire  _T_5433; // @[Bitwise.scala 50:65:@5461.4]
  wire  _T_5434; // @[Bitwise.scala 50:65:@5462.4]
  wire  _T_5435; // @[Bitwise.scala 50:65:@5463.4]
  wire  _T_5436; // @[Bitwise.scala 50:65:@5464.4]
  wire  _T_5437; // @[Bitwise.scala 50:65:@5465.4]
  wire  _T_5438; // @[Bitwise.scala 50:65:@5466.4]
  wire  _T_5439; // @[Bitwise.scala 50:65:@5467.4]
  wire  _T_5440; // @[Bitwise.scala 50:65:@5468.4]
  wire  _T_5441; // @[Bitwise.scala 50:65:@5469.4]
  wire  _T_5442; // @[Bitwise.scala 50:65:@5470.4]
  wire  _T_5443; // @[Bitwise.scala 50:65:@5471.4]
  wire  _T_5444; // @[Bitwise.scala 50:65:@5472.4]
  wire  _T_5445; // @[Bitwise.scala 50:65:@5473.4]
  wire  _T_5446; // @[Bitwise.scala 50:65:@5474.4]
  wire  _T_5447; // @[Bitwise.scala 50:65:@5475.4]
  wire  _T_5448; // @[Bitwise.scala 50:65:@5476.4]
  wire  _T_5449; // @[Bitwise.scala 50:65:@5477.4]
  wire  _T_5450; // @[Bitwise.scala 50:65:@5478.4]
  wire  _T_5451; // @[Bitwise.scala 50:65:@5479.4]
  wire  _T_5452; // @[Bitwise.scala 50:65:@5480.4]
  wire  _T_5453; // @[Bitwise.scala 50:65:@5481.4]
  wire  _T_5454; // @[Bitwise.scala 50:65:@5482.4]
  wire  _T_5455; // @[Bitwise.scala 50:65:@5483.4]
  wire  _T_5456; // @[Bitwise.scala 50:65:@5484.4]
  wire  _T_5457; // @[Bitwise.scala 50:65:@5485.4]
  wire  _T_5458; // @[Bitwise.scala 50:65:@5486.4]
  wire  _T_5459; // @[Bitwise.scala 50:65:@5487.4]
  wire  _T_5460; // @[Bitwise.scala 50:65:@5488.4]
  wire  _T_5461; // @[Bitwise.scala 50:65:@5489.4]
  wire  _T_5462; // @[Bitwise.scala 50:65:@5490.4]
  wire  _T_5463; // @[Bitwise.scala 50:65:@5491.4]
  wire  _T_5464; // @[Bitwise.scala 50:65:@5492.4]
  wire  _T_5465; // @[Bitwise.scala 50:65:@5493.4]
  wire  _T_5466; // @[Bitwise.scala 50:65:@5494.4]
  wire [1:0] _T_5467; // @[Bitwise.scala 48:55:@5495.4]
  wire [1:0] _T_5468; // @[Bitwise.scala 48:55:@5496.4]
  wire [2:0] _T_5469; // @[Bitwise.scala 48:55:@5497.4]
  wire [1:0] _T_5470; // @[Bitwise.scala 48:55:@5498.4]
  wire [1:0] _T_5471; // @[Bitwise.scala 48:55:@5499.4]
  wire [2:0] _T_5472; // @[Bitwise.scala 48:55:@5500.4]
  wire [3:0] _T_5473; // @[Bitwise.scala 48:55:@5501.4]
  wire [1:0] _T_5474; // @[Bitwise.scala 48:55:@5502.4]
  wire [1:0] _T_5475; // @[Bitwise.scala 48:55:@5503.4]
  wire [2:0] _T_5476; // @[Bitwise.scala 48:55:@5504.4]
  wire [1:0] _T_5477; // @[Bitwise.scala 48:55:@5505.4]
  wire [1:0] _T_5478; // @[Bitwise.scala 48:55:@5506.4]
  wire [1:0] _GEN_661; // @[Bitwise.scala 48:55:@5507.4]
  wire [2:0] _T_5479; // @[Bitwise.scala 48:55:@5507.4]
  wire [2:0] _GEN_662; // @[Bitwise.scala 48:55:@5508.4]
  wire [3:0] _T_5480; // @[Bitwise.scala 48:55:@5508.4]
  wire [3:0] _GEN_663; // @[Bitwise.scala 48:55:@5509.4]
  wire [4:0] _T_5481; // @[Bitwise.scala 48:55:@5509.4]
  wire [4:0] _GEN_664; // @[Bitwise.scala 48:55:@5510.4]
  wire [5:0] _T_5482; // @[Bitwise.scala 48:55:@5510.4]
  wire [1:0] _T_5483; // @[Bitwise.scala 48:55:@5511.4]
  wire [1:0] _T_5484; // @[Bitwise.scala 48:55:@5512.4]
  wire [2:0] _T_5485; // @[Bitwise.scala 48:55:@5513.4]
  wire [1:0] _T_5486; // @[Bitwise.scala 48:55:@5514.4]
  wire [1:0] _T_5487; // @[Bitwise.scala 48:55:@5515.4]
  wire [2:0] _T_5488; // @[Bitwise.scala 48:55:@5516.4]
  wire [3:0] _T_5489; // @[Bitwise.scala 48:55:@5517.4]
  wire [1:0] _T_5490; // @[Bitwise.scala 48:55:@5518.4]
  wire [1:0] _T_5491; // @[Bitwise.scala 48:55:@5519.4]
  wire [2:0] _T_5492; // @[Bitwise.scala 48:55:@5520.4]
  wire [1:0] _T_5493; // @[Bitwise.scala 48:55:@5521.4]
  wire [1:0] _T_5494; // @[Bitwise.scala 48:55:@5522.4]
  wire [1:0] _GEN_665; // @[Bitwise.scala 48:55:@5523.4]
  wire [2:0] _T_5495; // @[Bitwise.scala 48:55:@5523.4]
  wire [2:0] _GEN_666; // @[Bitwise.scala 48:55:@5524.4]
  wire [3:0] _T_5496; // @[Bitwise.scala 48:55:@5524.4]
  wire [3:0] _GEN_667; // @[Bitwise.scala 48:55:@5525.4]
  wire [4:0] _T_5497; // @[Bitwise.scala 48:55:@5525.4]
  wire [4:0] _GEN_668; // @[Bitwise.scala 48:55:@5526.4]
  wire [5:0] _T_5498; // @[Bitwise.scala 48:55:@5526.4]
  wire [6:0] _T_5499; // @[Bitwise.scala 48:55:@5527.4]
  wire [34:0] _T_5563; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5592.4]
  wire  _T_5564; // @[Bitwise.scala 50:65:@5593.4]
  wire  _T_5565; // @[Bitwise.scala 50:65:@5594.4]
  wire  _T_5566; // @[Bitwise.scala 50:65:@5595.4]
  wire  _T_5567; // @[Bitwise.scala 50:65:@5596.4]
  wire  _T_5568; // @[Bitwise.scala 50:65:@5597.4]
  wire  _T_5569; // @[Bitwise.scala 50:65:@5598.4]
  wire  _T_5570; // @[Bitwise.scala 50:65:@5599.4]
  wire  _T_5571; // @[Bitwise.scala 50:65:@5600.4]
  wire  _T_5572; // @[Bitwise.scala 50:65:@5601.4]
  wire  _T_5573; // @[Bitwise.scala 50:65:@5602.4]
  wire  _T_5574; // @[Bitwise.scala 50:65:@5603.4]
  wire  _T_5575; // @[Bitwise.scala 50:65:@5604.4]
  wire  _T_5576; // @[Bitwise.scala 50:65:@5605.4]
  wire  _T_5577; // @[Bitwise.scala 50:65:@5606.4]
  wire  _T_5578; // @[Bitwise.scala 50:65:@5607.4]
  wire  _T_5579; // @[Bitwise.scala 50:65:@5608.4]
  wire  _T_5580; // @[Bitwise.scala 50:65:@5609.4]
  wire  _T_5581; // @[Bitwise.scala 50:65:@5610.4]
  wire  _T_5582; // @[Bitwise.scala 50:65:@5611.4]
  wire  _T_5583; // @[Bitwise.scala 50:65:@5612.4]
  wire  _T_5584; // @[Bitwise.scala 50:65:@5613.4]
  wire  _T_5585; // @[Bitwise.scala 50:65:@5614.4]
  wire  _T_5586; // @[Bitwise.scala 50:65:@5615.4]
  wire  _T_5587; // @[Bitwise.scala 50:65:@5616.4]
  wire  _T_5588; // @[Bitwise.scala 50:65:@5617.4]
  wire  _T_5589; // @[Bitwise.scala 50:65:@5618.4]
  wire  _T_5590; // @[Bitwise.scala 50:65:@5619.4]
  wire  _T_5591; // @[Bitwise.scala 50:65:@5620.4]
  wire  _T_5592; // @[Bitwise.scala 50:65:@5621.4]
  wire  _T_5593; // @[Bitwise.scala 50:65:@5622.4]
  wire  _T_5594; // @[Bitwise.scala 50:65:@5623.4]
  wire  _T_5595; // @[Bitwise.scala 50:65:@5624.4]
  wire  _T_5596; // @[Bitwise.scala 50:65:@5625.4]
  wire  _T_5597; // @[Bitwise.scala 50:65:@5626.4]
  wire  _T_5598; // @[Bitwise.scala 50:65:@5627.4]
  wire [1:0] _T_5599; // @[Bitwise.scala 48:55:@5628.4]
  wire [1:0] _T_5600; // @[Bitwise.scala 48:55:@5629.4]
  wire [2:0] _T_5601; // @[Bitwise.scala 48:55:@5630.4]
  wire [1:0] _T_5602; // @[Bitwise.scala 48:55:@5631.4]
  wire [1:0] _T_5603; // @[Bitwise.scala 48:55:@5632.4]
  wire [2:0] _T_5604; // @[Bitwise.scala 48:55:@5633.4]
  wire [3:0] _T_5605; // @[Bitwise.scala 48:55:@5634.4]
  wire [1:0] _T_5606; // @[Bitwise.scala 48:55:@5635.4]
  wire [1:0] _T_5607; // @[Bitwise.scala 48:55:@5636.4]
  wire [2:0] _T_5608; // @[Bitwise.scala 48:55:@5637.4]
  wire [1:0] _T_5609; // @[Bitwise.scala 48:55:@5638.4]
  wire [1:0] _T_5610; // @[Bitwise.scala 48:55:@5639.4]
  wire [1:0] _GEN_669; // @[Bitwise.scala 48:55:@5640.4]
  wire [2:0] _T_5611; // @[Bitwise.scala 48:55:@5640.4]
  wire [2:0] _GEN_670; // @[Bitwise.scala 48:55:@5641.4]
  wire [3:0] _T_5612; // @[Bitwise.scala 48:55:@5641.4]
  wire [3:0] _GEN_671; // @[Bitwise.scala 48:55:@5642.4]
  wire [4:0] _T_5613; // @[Bitwise.scala 48:55:@5642.4]
  wire [4:0] _GEN_672; // @[Bitwise.scala 48:55:@5643.4]
  wire [5:0] _T_5614; // @[Bitwise.scala 48:55:@5643.4]
  wire [1:0] _T_5615; // @[Bitwise.scala 48:55:@5644.4]
  wire [1:0] _T_5616; // @[Bitwise.scala 48:55:@5645.4]
  wire [2:0] _T_5617; // @[Bitwise.scala 48:55:@5646.4]
  wire [1:0] _T_5618; // @[Bitwise.scala 48:55:@5647.4]
  wire [1:0] _T_5619; // @[Bitwise.scala 48:55:@5648.4]
  wire [1:0] _GEN_673; // @[Bitwise.scala 48:55:@5649.4]
  wire [2:0] _T_5620; // @[Bitwise.scala 48:55:@5649.4]
  wire [2:0] _GEN_674; // @[Bitwise.scala 48:55:@5650.4]
  wire [3:0] _T_5621; // @[Bitwise.scala 48:55:@5650.4]
  wire [3:0] _GEN_675; // @[Bitwise.scala 48:55:@5651.4]
  wire [4:0] _T_5622; // @[Bitwise.scala 48:55:@5651.4]
  wire [1:0] _T_5623; // @[Bitwise.scala 48:55:@5652.4]
  wire [1:0] _T_5624; // @[Bitwise.scala 48:55:@5653.4]
  wire [2:0] _T_5625; // @[Bitwise.scala 48:55:@5654.4]
  wire [1:0] _T_5626; // @[Bitwise.scala 48:55:@5655.4]
  wire [1:0] _T_5627; // @[Bitwise.scala 48:55:@5656.4]
  wire [1:0] _GEN_676; // @[Bitwise.scala 48:55:@5657.4]
  wire [2:0] _T_5628; // @[Bitwise.scala 48:55:@5657.4]
  wire [2:0] _GEN_677; // @[Bitwise.scala 48:55:@5658.4]
  wire [3:0] _T_5629; // @[Bitwise.scala 48:55:@5658.4]
  wire [3:0] _GEN_678; // @[Bitwise.scala 48:55:@5659.4]
  wire [4:0] _T_5630; // @[Bitwise.scala 48:55:@5659.4]
  wire [5:0] _T_5631; // @[Bitwise.scala 48:55:@5660.4]
  wire [6:0] _T_5632; // @[Bitwise.scala 48:55:@5661.4]
  wire [35:0] _T_5696; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5726.4]
  wire  _T_5697; // @[Bitwise.scala 50:65:@5727.4]
  wire  _T_5698; // @[Bitwise.scala 50:65:@5728.4]
  wire  _T_5699; // @[Bitwise.scala 50:65:@5729.4]
  wire  _T_5700; // @[Bitwise.scala 50:65:@5730.4]
  wire  _T_5701; // @[Bitwise.scala 50:65:@5731.4]
  wire  _T_5702; // @[Bitwise.scala 50:65:@5732.4]
  wire  _T_5703; // @[Bitwise.scala 50:65:@5733.4]
  wire  _T_5704; // @[Bitwise.scala 50:65:@5734.4]
  wire  _T_5705; // @[Bitwise.scala 50:65:@5735.4]
  wire  _T_5706; // @[Bitwise.scala 50:65:@5736.4]
  wire  _T_5707; // @[Bitwise.scala 50:65:@5737.4]
  wire  _T_5708; // @[Bitwise.scala 50:65:@5738.4]
  wire  _T_5709; // @[Bitwise.scala 50:65:@5739.4]
  wire  _T_5710; // @[Bitwise.scala 50:65:@5740.4]
  wire  _T_5711; // @[Bitwise.scala 50:65:@5741.4]
  wire  _T_5712; // @[Bitwise.scala 50:65:@5742.4]
  wire  _T_5713; // @[Bitwise.scala 50:65:@5743.4]
  wire  _T_5714; // @[Bitwise.scala 50:65:@5744.4]
  wire  _T_5715; // @[Bitwise.scala 50:65:@5745.4]
  wire  _T_5716; // @[Bitwise.scala 50:65:@5746.4]
  wire  _T_5717; // @[Bitwise.scala 50:65:@5747.4]
  wire  _T_5718; // @[Bitwise.scala 50:65:@5748.4]
  wire  _T_5719; // @[Bitwise.scala 50:65:@5749.4]
  wire  _T_5720; // @[Bitwise.scala 50:65:@5750.4]
  wire  _T_5721; // @[Bitwise.scala 50:65:@5751.4]
  wire  _T_5722; // @[Bitwise.scala 50:65:@5752.4]
  wire  _T_5723; // @[Bitwise.scala 50:65:@5753.4]
  wire  _T_5724; // @[Bitwise.scala 50:65:@5754.4]
  wire  _T_5725; // @[Bitwise.scala 50:65:@5755.4]
  wire  _T_5726; // @[Bitwise.scala 50:65:@5756.4]
  wire  _T_5727; // @[Bitwise.scala 50:65:@5757.4]
  wire  _T_5728; // @[Bitwise.scala 50:65:@5758.4]
  wire  _T_5729; // @[Bitwise.scala 50:65:@5759.4]
  wire  _T_5730; // @[Bitwise.scala 50:65:@5760.4]
  wire  _T_5731; // @[Bitwise.scala 50:65:@5761.4]
  wire  _T_5732; // @[Bitwise.scala 50:65:@5762.4]
  wire [1:0] _T_5733; // @[Bitwise.scala 48:55:@5763.4]
  wire [1:0] _T_5734; // @[Bitwise.scala 48:55:@5764.4]
  wire [2:0] _T_5735; // @[Bitwise.scala 48:55:@5765.4]
  wire [1:0] _T_5736; // @[Bitwise.scala 48:55:@5766.4]
  wire [1:0] _T_5737; // @[Bitwise.scala 48:55:@5767.4]
  wire [1:0] _GEN_679; // @[Bitwise.scala 48:55:@5768.4]
  wire [2:0] _T_5738; // @[Bitwise.scala 48:55:@5768.4]
  wire [2:0] _GEN_680; // @[Bitwise.scala 48:55:@5769.4]
  wire [3:0] _T_5739; // @[Bitwise.scala 48:55:@5769.4]
  wire [3:0] _GEN_681; // @[Bitwise.scala 48:55:@5770.4]
  wire [4:0] _T_5740; // @[Bitwise.scala 48:55:@5770.4]
  wire [1:0] _T_5741; // @[Bitwise.scala 48:55:@5771.4]
  wire [1:0] _T_5742; // @[Bitwise.scala 48:55:@5772.4]
  wire [2:0] _T_5743; // @[Bitwise.scala 48:55:@5773.4]
  wire [1:0] _T_5744; // @[Bitwise.scala 48:55:@5774.4]
  wire [1:0] _T_5745; // @[Bitwise.scala 48:55:@5775.4]
  wire [1:0] _GEN_682; // @[Bitwise.scala 48:55:@5776.4]
  wire [2:0] _T_5746; // @[Bitwise.scala 48:55:@5776.4]
  wire [2:0] _GEN_683; // @[Bitwise.scala 48:55:@5777.4]
  wire [3:0] _T_5747; // @[Bitwise.scala 48:55:@5777.4]
  wire [3:0] _GEN_684; // @[Bitwise.scala 48:55:@5778.4]
  wire [4:0] _T_5748; // @[Bitwise.scala 48:55:@5778.4]
  wire [5:0] _T_5749; // @[Bitwise.scala 48:55:@5779.4]
  wire [1:0] _T_5750; // @[Bitwise.scala 48:55:@5780.4]
  wire [1:0] _T_5751; // @[Bitwise.scala 48:55:@5781.4]
  wire [2:0] _T_5752; // @[Bitwise.scala 48:55:@5782.4]
  wire [1:0] _T_5753; // @[Bitwise.scala 48:55:@5783.4]
  wire [1:0] _T_5754; // @[Bitwise.scala 48:55:@5784.4]
  wire [1:0] _GEN_685; // @[Bitwise.scala 48:55:@5785.4]
  wire [2:0] _T_5755; // @[Bitwise.scala 48:55:@5785.4]
  wire [2:0] _GEN_686; // @[Bitwise.scala 48:55:@5786.4]
  wire [3:0] _T_5756; // @[Bitwise.scala 48:55:@5786.4]
  wire [3:0] _GEN_687; // @[Bitwise.scala 48:55:@5787.4]
  wire [4:0] _T_5757; // @[Bitwise.scala 48:55:@5787.4]
  wire [1:0] _T_5758; // @[Bitwise.scala 48:55:@5788.4]
  wire [1:0] _T_5759; // @[Bitwise.scala 48:55:@5789.4]
  wire [2:0] _T_5760; // @[Bitwise.scala 48:55:@5790.4]
  wire [1:0] _T_5761; // @[Bitwise.scala 48:55:@5791.4]
  wire [1:0] _T_5762; // @[Bitwise.scala 48:55:@5792.4]
  wire [1:0] _GEN_688; // @[Bitwise.scala 48:55:@5793.4]
  wire [2:0] _T_5763; // @[Bitwise.scala 48:55:@5793.4]
  wire [2:0] _GEN_689; // @[Bitwise.scala 48:55:@5794.4]
  wire [3:0] _T_5764; // @[Bitwise.scala 48:55:@5794.4]
  wire [3:0] _GEN_690; // @[Bitwise.scala 48:55:@5795.4]
  wire [4:0] _T_5765; // @[Bitwise.scala 48:55:@5795.4]
  wire [5:0] _T_5766; // @[Bitwise.scala 48:55:@5796.4]
  wire [6:0] _T_5767; // @[Bitwise.scala 48:55:@5797.4]
  wire [36:0] _T_5831; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5862.4]
  wire  _T_5832; // @[Bitwise.scala 50:65:@5863.4]
  wire  _T_5833; // @[Bitwise.scala 50:65:@5864.4]
  wire  _T_5834; // @[Bitwise.scala 50:65:@5865.4]
  wire  _T_5835; // @[Bitwise.scala 50:65:@5866.4]
  wire  _T_5836; // @[Bitwise.scala 50:65:@5867.4]
  wire  _T_5837; // @[Bitwise.scala 50:65:@5868.4]
  wire  _T_5838; // @[Bitwise.scala 50:65:@5869.4]
  wire  _T_5839; // @[Bitwise.scala 50:65:@5870.4]
  wire  _T_5840; // @[Bitwise.scala 50:65:@5871.4]
  wire  _T_5841; // @[Bitwise.scala 50:65:@5872.4]
  wire  _T_5842; // @[Bitwise.scala 50:65:@5873.4]
  wire  _T_5843; // @[Bitwise.scala 50:65:@5874.4]
  wire  _T_5844; // @[Bitwise.scala 50:65:@5875.4]
  wire  _T_5845; // @[Bitwise.scala 50:65:@5876.4]
  wire  _T_5846; // @[Bitwise.scala 50:65:@5877.4]
  wire  _T_5847; // @[Bitwise.scala 50:65:@5878.4]
  wire  _T_5848; // @[Bitwise.scala 50:65:@5879.4]
  wire  _T_5849; // @[Bitwise.scala 50:65:@5880.4]
  wire  _T_5850; // @[Bitwise.scala 50:65:@5881.4]
  wire  _T_5851; // @[Bitwise.scala 50:65:@5882.4]
  wire  _T_5852; // @[Bitwise.scala 50:65:@5883.4]
  wire  _T_5853; // @[Bitwise.scala 50:65:@5884.4]
  wire  _T_5854; // @[Bitwise.scala 50:65:@5885.4]
  wire  _T_5855; // @[Bitwise.scala 50:65:@5886.4]
  wire  _T_5856; // @[Bitwise.scala 50:65:@5887.4]
  wire  _T_5857; // @[Bitwise.scala 50:65:@5888.4]
  wire  _T_5858; // @[Bitwise.scala 50:65:@5889.4]
  wire  _T_5859; // @[Bitwise.scala 50:65:@5890.4]
  wire  _T_5860; // @[Bitwise.scala 50:65:@5891.4]
  wire  _T_5861; // @[Bitwise.scala 50:65:@5892.4]
  wire  _T_5862; // @[Bitwise.scala 50:65:@5893.4]
  wire  _T_5863; // @[Bitwise.scala 50:65:@5894.4]
  wire  _T_5864; // @[Bitwise.scala 50:65:@5895.4]
  wire  _T_5865; // @[Bitwise.scala 50:65:@5896.4]
  wire  _T_5866; // @[Bitwise.scala 50:65:@5897.4]
  wire  _T_5867; // @[Bitwise.scala 50:65:@5898.4]
  wire  _T_5868; // @[Bitwise.scala 50:65:@5899.4]
  wire [1:0] _T_5869; // @[Bitwise.scala 48:55:@5900.4]
  wire [1:0] _T_5870; // @[Bitwise.scala 48:55:@5901.4]
  wire [2:0] _T_5871; // @[Bitwise.scala 48:55:@5902.4]
  wire [1:0] _T_5872; // @[Bitwise.scala 48:55:@5903.4]
  wire [1:0] _T_5873; // @[Bitwise.scala 48:55:@5904.4]
  wire [1:0] _GEN_691; // @[Bitwise.scala 48:55:@5905.4]
  wire [2:0] _T_5874; // @[Bitwise.scala 48:55:@5905.4]
  wire [2:0] _GEN_692; // @[Bitwise.scala 48:55:@5906.4]
  wire [3:0] _T_5875; // @[Bitwise.scala 48:55:@5906.4]
  wire [3:0] _GEN_693; // @[Bitwise.scala 48:55:@5907.4]
  wire [4:0] _T_5876; // @[Bitwise.scala 48:55:@5907.4]
  wire [1:0] _T_5877; // @[Bitwise.scala 48:55:@5908.4]
  wire [1:0] _T_5878; // @[Bitwise.scala 48:55:@5909.4]
  wire [2:0] _T_5879; // @[Bitwise.scala 48:55:@5910.4]
  wire [1:0] _T_5880; // @[Bitwise.scala 48:55:@5911.4]
  wire [1:0] _T_5881; // @[Bitwise.scala 48:55:@5912.4]
  wire [1:0] _GEN_694; // @[Bitwise.scala 48:55:@5913.4]
  wire [2:0] _T_5882; // @[Bitwise.scala 48:55:@5913.4]
  wire [2:0] _GEN_695; // @[Bitwise.scala 48:55:@5914.4]
  wire [3:0] _T_5883; // @[Bitwise.scala 48:55:@5914.4]
  wire [3:0] _GEN_696; // @[Bitwise.scala 48:55:@5915.4]
  wire [4:0] _T_5884; // @[Bitwise.scala 48:55:@5915.4]
  wire [5:0] _T_5885; // @[Bitwise.scala 48:55:@5916.4]
  wire [1:0] _T_5886; // @[Bitwise.scala 48:55:@5917.4]
  wire [1:0] _T_5887; // @[Bitwise.scala 48:55:@5918.4]
  wire [2:0] _T_5888; // @[Bitwise.scala 48:55:@5919.4]
  wire [1:0] _T_5889; // @[Bitwise.scala 48:55:@5920.4]
  wire [1:0] _T_5890; // @[Bitwise.scala 48:55:@5921.4]
  wire [1:0] _GEN_697; // @[Bitwise.scala 48:55:@5922.4]
  wire [2:0] _T_5891; // @[Bitwise.scala 48:55:@5922.4]
  wire [2:0] _GEN_698; // @[Bitwise.scala 48:55:@5923.4]
  wire [3:0] _T_5892; // @[Bitwise.scala 48:55:@5923.4]
  wire [3:0] _GEN_699; // @[Bitwise.scala 48:55:@5924.4]
  wire [4:0] _T_5893; // @[Bitwise.scala 48:55:@5924.4]
  wire [1:0] _T_5894; // @[Bitwise.scala 48:55:@5925.4]
  wire [1:0] _T_5895; // @[Bitwise.scala 48:55:@5926.4]
  wire [1:0] _GEN_700; // @[Bitwise.scala 48:55:@5927.4]
  wire [2:0] _T_5896; // @[Bitwise.scala 48:55:@5927.4]
  wire [2:0] _GEN_701; // @[Bitwise.scala 48:55:@5928.4]
  wire [3:0] _T_5897; // @[Bitwise.scala 48:55:@5928.4]
  wire [1:0] _T_5898; // @[Bitwise.scala 48:55:@5929.4]
  wire [1:0] _T_5899; // @[Bitwise.scala 48:55:@5930.4]
  wire [1:0] _GEN_702; // @[Bitwise.scala 48:55:@5931.4]
  wire [2:0] _T_5900; // @[Bitwise.scala 48:55:@5931.4]
  wire [2:0] _GEN_703; // @[Bitwise.scala 48:55:@5932.4]
  wire [3:0] _T_5901; // @[Bitwise.scala 48:55:@5932.4]
  wire [4:0] _T_5902; // @[Bitwise.scala 48:55:@5933.4]
  wire [5:0] _T_5903; // @[Bitwise.scala 48:55:@5934.4]
  wire [6:0] _T_5904; // @[Bitwise.scala 48:55:@5935.4]
  wire [37:0] _T_5968; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6000.4]
  wire  _T_5969; // @[Bitwise.scala 50:65:@6001.4]
  wire  _T_5970; // @[Bitwise.scala 50:65:@6002.4]
  wire  _T_5971; // @[Bitwise.scala 50:65:@6003.4]
  wire  _T_5972; // @[Bitwise.scala 50:65:@6004.4]
  wire  _T_5973; // @[Bitwise.scala 50:65:@6005.4]
  wire  _T_5974; // @[Bitwise.scala 50:65:@6006.4]
  wire  _T_5975; // @[Bitwise.scala 50:65:@6007.4]
  wire  _T_5976; // @[Bitwise.scala 50:65:@6008.4]
  wire  _T_5977; // @[Bitwise.scala 50:65:@6009.4]
  wire  _T_5978; // @[Bitwise.scala 50:65:@6010.4]
  wire  _T_5979; // @[Bitwise.scala 50:65:@6011.4]
  wire  _T_5980; // @[Bitwise.scala 50:65:@6012.4]
  wire  _T_5981; // @[Bitwise.scala 50:65:@6013.4]
  wire  _T_5982; // @[Bitwise.scala 50:65:@6014.4]
  wire  _T_5983; // @[Bitwise.scala 50:65:@6015.4]
  wire  _T_5984; // @[Bitwise.scala 50:65:@6016.4]
  wire  _T_5985; // @[Bitwise.scala 50:65:@6017.4]
  wire  _T_5986; // @[Bitwise.scala 50:65:@6018.4]
  wire  _T_5987; // @[Bitwise.scala 50:65:@6019.4]
  wire  _T_5988; // @[Bitwise.scala 50:65:@6020.4]
  wire  _T_5989; // @[Bitwise.scala 50:65:@6021.4]
  wire  _T_5990; // @[Bitwise.scala 50:65:@6022.4]
  wire  _T_5991; // @[Bitwise.scala 50:65:@6023.4]
  wire  _T_5992; // @[Bitwise.scala 50:65:@6024.4]
  wire  _T_5993; // @[Bitwise.scala 50:65:@6025.4]
  wire  _T_5994; // @[Bitwise.scala 50:65:@6026.4]
  wire  _T_5995; // @[Bitwise.scala 50:65:@6027.4]
  wire  _T_5996; // @[Bitwise.scala 50:65:@6028.4]
  wire  _T_5997; // @[Bitwise.scala 50:65:@6029.4]
  wire  _T_5998; // @[Bitwise.scala 50:65:@6030.4]
  wire  _T_5999; // @[Bitwise.scala 50:65:@6031.4]
  wire  _T_6000; // @[Bitwise.scala 50:65:@6032.4]
  wire  _T_6001; // @[Bitwise.scala 50:65:@6033.4]
  wire  _T_6002; // @[Bitwise.scala 50:65:@6034.4]
  wire  _T_6003; // @[Bitwise.scala 50:65:@6035.4]
  wire  _T_6004; // @[Bitwise.scala 50:65:@6036.4]
  wire  _T_6005; // @[Bitwise.scala 50:65:@6037.4]
  wire  _T_6006; // @[Bitwise.scala 50:65:@6038.4]
  wire [1:0] _T_6007; // @[Bitwise.scala 48:55:@6039.4]
  wire [1:0] _T_6008; // @[Bitwise.scala 48:55:@6040.4]
  wire [2:0] _T_6009; // @[Bitwise.scala 48:55:@6041.4]
  wire [1:0] _T_6010; // @[Bitwise.scala 48:55:@6042.4]
  wire [1:0] _T_6011; // @[Bitwise.scala 48:55:@6043.4]
  wire [1:0] _GEN_704; // @[Bitwise.scala 48:55:@6044.4]
  wire [2:0] _T_6012; // @[Bitwise.scala 48:55:@6044.4]
  wire [2:0] _GEN_705; // @[Bitwise.scala 48:55:@6045.4]
  wire [3:0] _T_6013; // @[Bitwise.scala 48:55:@6045.4]
  wire [3:0] _GEN_706; // @[Bitwise.scala 48:55:@6046.4]
  wire [4:0] _T_6014; // @[Bitwise.scala 48:55:@6046.4]
  wire [1:0] _T_6015; // @[Bitwise.scala 48:55:@6047.4]
  wire [1:0] _T_6016; // @[Bitwise.scala 48:55:@6048.4]
  wire [1:0] _GEN_707; // @[Bitwise.scala 48:55:@6049.4]
  wire [2:0] _T_6017; // @[Bitwise.scala 48:55:@6049.4]
  wire [2:0] _GEN_708; // @[Bitwise.scala 48:55:@6050.4]
  wire [3:0] _T_6018; // @[Bitwise.scala 48:55:@6050.4]
  wire [1:0] _T_6019; // @[Bitwise.scala 48:55:@6051.4]
  wire [1:0] _T_6020; // @[Bitwise.scala 48:55:@6052.4]
  wire [1:0] _GEN_709; // @[Bitwise.scala 48:55:@6053.4]
  wire [2:0] _T_6021; // @[Bitwise.scala 48:55:@6053.4]
  wire [2:0] _GEN_710; // @[Bitwise.scala 48:55:@6054.4]
  wire [3:0] _T_6022; // @[Bitwise.scala 48:55:@6054.4]
  wire [4:0] _T_6023; // @[Bitwise.scala 48:55:@6055.4]
  wire [5:0] _T_6024; // @[Bitwise.scala 48:55:@6056.4]
  wire [1:0] _T_6025; // @[Bitwise.scala 48:55:@6057.4]
  wire [1:0] _T_6026; // @[Bitwise.scala 48:55:@6058.4]
  wire [2:0] _T_6027; // @[Bitwise.scala 48:55:@6059.4]
  wire [1:0] _T_6028; // @[Bitwise.scala 48:55:@6060.4]
  wire [1:0] _T_6029; // @[Bitwise.scala 48:55:@6061.4]
  wire [1:0] _GEN_711; // @[Bitwise.scala 48:55:@6062.4]
  wire [2:0] _T_6030; // @[Bitwise.scala 48:55:@6062.4]
  wire [2:0] _GEN_712; // @[Bitwise.scala 48:55:@6063.4]
  wire [3:0] _T_6031; // @[Bitwise.scala 48:55:@6063.4]
  wire [3:0] _GEN_713; // @[Bitwise.scala 48:55:@6064.4]
  wire [4:0] _T_6032; // @[Bitwise.scala 48:55:@6064.4]
  wire [1:0] _T_6033; // @[Bitwise.scala 48:55:@6065.4]
  wire [1:0] _T_6034; // @[Bitwise.scala 48:55:@6066.4]
  wire [1:0] _GEN_714; // @[Bitwise.scala 48:55:@6067.4]
  wire [2:0] _T_6035; // @[Bitwise.scala 48:55:@6067.4]
  wire [2:0] _GEN_715; // @[Bitwise.scala 48:55:@6068.4]
  wire [3:0] _T_6036; // @[Bitwise.scala 48:55:@6068.4]
  wire [1:0] _T_6037; // @[Bitwise.scala 48:55:@6069.4]
  wire [1:0] _T_6038; // @[Bitwise.scala 48:55:@6070.4]
  wire [1:0] _GEN_716; // @[Bitwise.scala 48:55:@6071.4]
  wire [2:0] _T_6039; // @[Bitwise.scala 48:55:@6071.4]
  wire [2:0] _GEN_717; // @[Bitwise.scala 48:55:@6072.4]
  wire [3:0] _T_6040; // @[Bitwise.scala 48:55:@6072.4]
  wire [4:0] _T_6041; // @[Bitwise.scala 48:55:@6073.4]
  wire [5:0] _T_6042; // @[Bitwise.scala 48:55:@6074.4]
  wire [6:0] _T_6043; // @[Bitwise.scala 48:55:@6075.4]
  wire [38:0] _T_6107; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6140.4]
  wire  _T_6108; // @[Bitwise.scala 50:65:@6141.4]
  wire  _T_6109; // @[Bitwise.scala 50:65:@6142.4]
  wire  _T_6110; // @[Bitwise.scala 50:65:@6143.4]
  wire  _T_6111; // @[Bitwise.scala 50:65:@6144.4]
  wire  _T_6112; // @[Bitwise.scala 50:65:@6145.4]
  wire  _T_6113; // @[Bitwise.scala 50:65:@6146.4]
  wire  _T_6114; // @[Bitwise.scala 50:65:@6147.4]
  wire  _T_6115; // @[Bitwise.scala 50:65:@6148.4]
  wire  _T_6116; // @[Bitwise.scala 50:65:@6149.4]
  wire  _T_6117; // @[Bitwise.scala 50:65:@6150.4]
  wire  _T_6118; // @[Bitwise.scala 50:65:@6151.4]
  wire  _T_6119; // @[Bitwise.scala 50:65:@6152.4]
  wire  _T_6120; // @[Bitwise.scala 50:65:@6153.4]
  wire  _T_6121; // @[Bitwise.scala 50:65:@6154.4]
  wire  _T_6122; // @[Bitwise.scala 50:65:@6155.4]
  wire  _T_6123; // @[Bitwise.scala 50:65:@6156.4]
  wire  _T_6124; // @[Bitwise.scala 50:65:@6157.4]
  wire  _T_6125; // @[Bitwise.scala 50:65:@6158.4]
  wire  _T_6126; // @[Bitwise.scala 50:65:@6159.4]
  wire  _T_6127; // @[Bitwise.scala 50:65:@6160.4]
  wire  _T_6128; // @[Bitwise.scala 50:65:@6161.4]
  wire  _T_6129; // @[Bitwise.scala 50:65:@6162.4]
  wire  _T_6130; // @[Bitwise.scala 50:65:@6163.4]
  wire  _T_6131; // @[Bitwise.scala 50:65:@6164.4]
  wire  _T_6132; // @[Bitwise.scala 50:65:@6165.4]
  wire  _T_6133; // @[Bitwise.scala 50:65:@6166.4]
  wire  _T_6134; // @[Bitwise.scala 50:65:@6167.4]
  wire  _T_6135; // @[Bitwise.scala 50:65:@6168.4]
  wire  _T_6136; // @[Bitwise.scala 50:65:@6169.4]
  wire  _T_6137; // @[Bitwise.scala 50:65:@6170.4]
  wire  _T_6138; // @[Bitwise.scala 50:65:@6171.4]
  wire  _T_6139; // @[Bitwise.scala 50:65:@6172.4]
  wire  _T_6140; // @[Bitwise.scala 50:65:@6173.4]
  wire  _T_6141; // @[Bitwise.scala 50:65:@6174.4]
  wire  _T_6142; // @[Bitwise.scala 50:65:@6175.4]
  wire  _T_6143; // @[Bitwise.scala 50:65:@6176.4]
  wire  _T_6144; // @[Bitwise.scala 50:65:@6177.4]
  wire  _T_6145; // @[Bitwise.scala 50:65:@6178.4]
  wire  _T_6146; // @[Bitwise.scala 50:65:@6179.4]
  wire [1:0] _T_6147; // @[Bitwise.scala 48:55:@6180.4]
  wire [1:0] _T_6148; // @[Bitwise.scala 48:55:@6181.4]
  wire [2:0] _T_6149; // @[Bitwise.scala 48:55:@6182.4]
  wire [1:0] _T_6150; // @[Bitwise.scala 48:55:@6183.4]
  wire [1:0] _T_6151; // @[Bitwise.scala 48:55:@6184.4]
  wire [1:0] _GEN_718; // @[Bitwise.scala 48:55:@6185.4]
  wire [2:0] _T_6152; // @[Bitwise.scala 48:55:@6185.4]
  wire [2:0] _GEN_719; // @[Bitwise.scala 48:55:@6186.4]
  wire [3:0] _T_6153; // @[Bitwise.scala 48:55:@6186.4]
  wire [3:0] _GEN_720; // @[Bitwise.scala 48:55:@6187.4]
  wire [4:0] _T_6154; // @[Bitwise.scala 48:55:@6187.4]
  wire [1:0] _T_6155; // @[Bitwise.scala 48:55:@6188.4]
  wire [1:0] _T_6156; // @[Bitwise.scala 48:55:@6189.4]
  wire [1:0] _GEN_721; // @[Bitwise.scala 48:55:@6190.4]
  wire [2:0] _T_6157; // @[Bitwise.scala 48:55:@6190.4]
  wire [2:0] _GEN_722; // @[Bitwise.scala 48:55:@6191.4]
  wire [3:0] _T_6158; // @[Bitwise.scala 48:55:@6191.4]
  wire [1:0] _T_6159; // @[Bitwise.scala 48:55:@6192.4]
  wire [1:0] _T_6160; // @[Bitwise.scala 48:55:@6193.4]
  wire [1:0] _GEN_723; // @[Bitwise.scala 48:55:@6194.4]
  wire [2:0] _T_6161; // @[Bitwise.scala 48:55:@6194.4]
  wire [2:0] _GEN_724; // @[Bitwise.scala 48:55:@6195.4]
  wire [3:0] _T_6162; // @[Bitwise.scala 48:55:@6195.4]
  wire [4:0] _T_6163; // @[Bitwise.scala 48:55:@6196.4]
  wire [5:0] _T_6164; // @[Bitwise.scala 48:55:@6197.4]
  wire [1:0] _T_6165; // @[Bitwise.scala 48:55:@6198.4]
  wire [1:0] _T_6166; // @[Bitwise.scala 48:55:@6199.4]
  wire [1:0] _GEN_725; // @[Bitwise.scala 48:55:@6200.4]
  wire [2:0] _T_6167; // @[Bitwise.scala 48:55:@6200.4]
  wire [2:0] _GEN_726; // @[Bitwise.scala 48:55:@6201.4]
  wire [3:0] _T_6168; // @[Bitwise.scala 48:55:@6201.4]
  wire [1:0] _T_6169; // @[Bitwise.scala 48:55:@6202.4]
  wire [1:0] _T_6170; // @[Bitwise.scala 48:55:@6203.4]
  wire [1:0] _GEN_727; // @[Bitwise.scala 48:55:@6204.4]
  wire [2:0] _T_6171; // @[Bitwise.scala 48:55:@6204.4]
  wire [2:0] _GEN_728; // @[Bitwise.scala 48:55:@6205.4]
  wire [3:0] _T_6172; // @[Bitwise.scala 48:55:@6205.4]
  wire [4:0] _T_6173; // @[Bitwise.scala 48:55:@6206.4]
  wire [1:0] _T_6174; // @[Bitwise.scala 48:55:@6207.4]
  wire [1:0] _T_6175; // @[Bitwise.scala 48:55:@6208.4]
  wire [1:0] _GEN_729; // @[Bitwise.scala 48:55:@6209.4]
  wire [2:0] _T_6176; // @[Bitwise.scala 48:55:@6209.4]
  wire [2:0] _GEN_730; // @[Bitwise.scala 48:55:@6210.4]
  wire [3:0] _T_6177; // @[Bitwise.scala 48:55:@6210.4]
  wire [1:0] _T_6178; // @[Bitwise.scala 48:55:@6211.4]
  wire [1:0] _T_6179; // @[Bitwise.scala 48:55:@6212.4]
  wire [1:0] _GEN_731; // @[Bitwise.scala 48:55:@6213.4]
  wire [2:0] _T_6180; // @[Bitwise.scala 48:55:@6213.4]
  wire [2:0] _GEN_732; // @[Bitwise.scala 48:55:@6214.4]
  wire [3:0] _T_6181; // @[Bitwise.scala 48:55:@6214.4]
  wire [4:0] _T_6182; // @[Bitwise.scala 48:55:@6215.4]
  wire [5:0] _T_6183; // @[Bitwise.scala 48:55:@6216.4]
  wire [6:0] _T_6184; // @[Bitwise.scala 48:55:@6217.4]
  wire [39:0] _T_6248; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6282.4]
  wire  _T_6249; // @[Bitwise.scala 50:65:@6283.4]
  wire  _T_6250; // @[Bitwise.scala 50:65:@6284.4]
  wire  _T_6251; // @[Bitwise.scala 50:65:@6285.4]
  wire  _T_6252; // @[Bitwise.scala 50:65:@6286.4]
  wire  _T_6253; // @[Bitwise.scala 50:65:@6287.4]
  wire  _T_6254; // @[Bitwise.scala 50:65:@6288.4]
  wire  _T_6255; // @[Bitwise.scala 50:65:@6289.4]
  wire  _T_6256; // @[Bitwise.scala 50:65:@6290.4]
  wire  _T_6257; // @[Bitwise.scala 50:65:@6291.4]
  wire  _T_6258; // @[Bitwise.scala 50:65:@6292.4]
  wire  _T_6259; // @[Bitwise.scala 50:65:@6293.4]
  wire  _T_6260; // @[Bitwise.scala 50:65:@6294.4]
  wire  _T_6261; // @[Bitwise.scala 50:65:@6295.4]
  wire  _T_6262; // @[Bitwise.scala 50:65:@6296.4]
  wire  _T_6263; // @[Bitwise.scala 50:65:@6297.4]
  wire  _T_6264; // @[Bitwise.scala 50:65:@6298.4]
  wire  _T_6265; // @[Bitwise.scala 50:65:@6299.4]
  wire  _T_6266; // @[Bitwise.scala 50:65:@6300.4]
  wire  _T_6267; // @[Bitwise.scala 50:65:@6301.4]
  wire  _T_6268; // @[Bitwise.scala 50:65:@6302.4]
  wire  _T_6269; // @[Bitwise.scala 50:65:@6303.4]
  wire  _T_6270; // @[Bitwise.scala 50:65:@6304.4]
  wire  _T_6271; // @[Bitwise.scala 50:65:@6305.4]
  wire  _T_6272; // @[Bitwise.scala 50:65:@6306.4]
  wire  _T_6273; // @[Bitwise.scala 50:65:@6307.4]
  wire  _T_6274; // @[Bitwise.scala 50:65:@6308.4]
  wire  _T_6275; // @[Bitwise.scala 50:65:@6309.4]
  wire  _T_6276; // @[Bitwise.scala 50:65:@6310.4]
  wire  _T_6277; // @[Bitwise.scala 50:65:@6311.4]
  wire  _T_6278; // @[Bitwise.scala 50:65:@6312.4]
  wire  _T_6279; // @[Bitwise.scala 50:65:@6313.4]
  wire  _T_6280; // @[Bitwise.scala 50:65:@6314.4]
  wire  _T_6281; // @[Bitwise.scala 50:65:@6315.4]
  wire  _T_6282; // @[Bitwise.scala 50:65:@6316.4]
  wire  _T_6283; // @[Bitwise.scala 50:65:@6317.4]
  wire  _T_6284; // @[Bitwise.scala 50:65:@6318.4]
  wire  _T_6285; // @[Bitwise.scala 50:65:@6319.4]
  wire  _T_6286; // @[Bitwise.scala 50:65:@6320.4]
  wire  _T_6287; // @[Bitwise.scala 50:65:@6321.4]
  wire  _T_6288; // @[Bitwise.scala 50:65:@6322.4]
  wire [1:0] _T_6289; // @[Bitwise.scala 48:55:@6323.4]
  wire [1:0] _T_6290; // @[Bitwise.scala 48:55:@6324.4]
  wire [1:0] _GEN_733; // @[Bitwise.scala 48:55:@6325.4]
  wire [2:0] _T_6291; // @[Bitwise.scala 48:55:@6325.4]
  wire [2:0] _GEN_734; // @[Bitwise.scala 48:55:@6326.4]
  wire [3:0] _T_6292; // @[Bitwise.scala 48:55:@6326.4]
  wire [1:0] _T_6293; // @[Bitwise.scala 48:55:@6327.4]
  wire [1:0] _T_6294; // @[Bitwise.scala 48:55:@6328.4]
  wire [1:0] _GEN_735; // @[Bitwise.scala 48:55:@6329.4]
  wire [2:0] _T_6295; // @[Bitwise.scala 48:55:@6329.4]
  wire [2:0] _GEN_736; // @[Bitwise.scala 48:55:@6330.4]
  wire [3:0] _T_6296; // @[Bitwise.scala 48:55:@6330.4]
  wire [4:0] _T_6297; // @[Bitwise.scala 48:55:@6331.4]
  wire [1:0] _T_6298; // @[Bitwise.scala 48:55:@6332.4]
  wire [1:0] _T_6299; // @[Bitwise.scala 48:55:@6333.4]
  wire [1:0] _GEN_737; // @[Bitwise.scala 48:55:@6334.4]
  wire [2:0] _T_6300; // @[Bitwise.scala 48:55:@6334.4]
  wire [2:0] _GEN_738; // @[Bitwise.scala 48:55:@6335.4]
  wire [3:0] _T_6301; // @[Bitwise.scala 48:55:@6335.4]
  wire [1:0] _T_6302; // @[Bitwise.scala 48:55:@6336.4]
  wire [1:0] _T_6303; // @[Bitwise.scala 48:55:@6337.4]
  wire [1:0] _GEN_739; // @[Bitwise.scala 48:55:@6338.4]
  wire [2:0] _T_6304; // @[Bitwise.scala 48:55:@6338.4]
  wire [2:0] _GEN_740; // @[Bitwise.scala 48:55:@6339.4]
  wire [3:0] _T_6305; // @[Bitwise.scala 48:55:@6339.4]
  wire [4:0] _T_6306; // @[Bitwise.scala 48:55:@6340.4]
  wire [5:0] _T_6307; // @[Bitwise.scala 48:55:@6341.4]
  wire [1:0] _T_6308; // @[Bitwise.scala 48:55:@6342.4]
  wire [1:0] _T_6309; // @[Bitwise.scala 48:55:@6343.4]
  wire [1:0] _GEN_741; // @[Bitwise.scala 48:55:@6344.4]
  wire [2:0] _T_6310; // @[Bitwise.scala 48:55:@6344.4]
  wire [2:0] _GEN_742; // @[Bitwise.scala 48:55:@6345.4]
  wire [3:0] _T_6311; // @[Bitwise.scala 48:55:@6345.4]
  wire [1:0] _T_6312; // @[Bitwise.scala 48:55:@6346.4]
  wire [1:0] _T_6313; // @[Bitwise.scala 48:55:@6347.4]
  wire [1:0] _GEN_743; // @[Bitwise.scala 48:55:@6348.4]
  wire [2:0] _T_6314; // @[Bitwise.scala 48:55:@6348.4]
  wire [2:0] _GEN_744; // @[Bitwise.scala 48:55:@6349.4]
  wire [3:0] _T_6315; // @[Bitwise.scala 48:55:@6349.4]
  wire [4:0] _T_6316; // @[Bitwise.scala 48:55:@6350.4]
  wire [1:0] _T_6317; // @[Bitwise.scala 48:55:@6351.4]
  wire [1:0] _T_6318; // @[Bitwise.scala 48:55:@6352.4]
  wire [1:0] _GEN_745; // @[Bitwise.scala 48:55:@6353.4]
  wire [2:0] _T_6319; // @[Bitwise.scala 48:55:@6353.4]
  wire [2:0] _GEN_746; // @[Bitwise.scala 48:55:@6354.4]
  wire [3:0] _T_6320; // @[Bitwise.scala 48:55:@6354.4]
  wire [1:0] _T_6321; // @[Bitwise.scala 48:55:@6355.4]
  wire [1:0] _T_6322; // @[Bitwise.scala 48:55:@6356.4]
  wire [1:0] _GEN_747; // @[Bitwise.scala 48:55:@6357.4]
  wire [2:0] _T_6323; // @[Bitwise.scala 48:55:@6357.4]
  wire [2:0] _GEN_748; // @[Bitwise.scala 48:55:@6358.4]
  wire [3:0] _T_6324; // @[Bitwise.scala 48:55:@6358.4]
  wire [4:0] _T_6325; // @[Bitwise.scala 48:55:@6359.4]
  wire [5:0] _T_6326; // @[Bitwise.scala 48:55:@6360.4]
  wire [6:0] _T_6327; // @[Bitwise.scala 48:55:@6361.4]
  wire [40:0] _T_6391; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6426.4]
  wire  _T_6392; // @[Bitwise.scala 50:65:@6427.4]
  wire  _T_6393; // @[Bitwise.scala 50:65:@6428.4]
  wire  _T_6394; // @[Bitwise.scala 50:65:@6429.4]
  wire  _T_6395; // @[Bitwise.scala 50:65:@6430.4]
  wire  _T_6396; // @[Bitwise.scala 50:65:@6431.4]
  wire  _T_6397; // @[Bitwise.scala 50:65:@6432.4]
  wire  _T_6398; // @[Bitwise.scala 50:65:@6433.4]
  wire  _T_6399; // @[Bitwise.scala 50:65:@6434.4]
  wire  _T_6400; // @[Bitwise.scala 50:65:@6435.4]
  wire  _T_6401; // @[Bitwise.scala 50:65:@6436.4]
  wire  _T_6402; // @[Bitwise.scala 50:65:@6437.4]
  wire  _T_6403; // @[Bitwise.scala 50:65:@6438.4]
  wire  _T_6404; // @[Bitwise.scala 50:65:@6439.4]
  wire  _T_6405; // @[Bitwise.scala 50:65:@6440.4]
  wire  _T_6406; // @[Bitwise.scala 50:65:@6441.4]
  wire  _T_6407; // @[Bitwise.scala 50:65:@6442.4]
  wire  _T_6408; // @[Bitwise.scala 50:65:@6443.4]
  wire  _T_6409; // @[Bitwise.scala 50:65:@6444.4]
  wire  _T_6410; // @[Bitwise.scala 50:65:@6445.4]
  wire  _T_6411; // @[Bitwise.scala 50:65:@6446.4]
  wire  _T_6412; // @[Bitwise.scala 50:65:@6447.4]
  wire  _T_6413; // @[Bitwise.scala 50:65:@6448.4]
  wire  _T_6414; // @[Bitwise.scala 50:65:@6449.4]
  wire  _T_6415; // @[Bitwise.scala 50:65:@6450.4]
  wire  _T_6416; // @[Bitwise.scala 50:65:@6451.4]
  wire  _T_6417; // @[Bitwise.scala 50:65:@6452.4]
  wire  _T_6418; // @[Bitwise.scala 50:65:@6453.4]
  wire  _T_6419; // @[Bitwise.scala 50:65:@6454.4]
  wire  _T_6420; // @[Bitwise.scala 50:65:@6455.4]
  wire  _T_6421; // @[Bitwise.scala 50:65:@6456.4]
  wire  _T_6422; // @[Bitwise.scala 50:65:@6457.4]
  wire  _T_6423; // @[Bitwise.scala 50:65:@6458.4]
  wire  _T_6424; // @[Bitwise.scala 50:65:@6459.4]
  wire  _T_6425; // @[Bitwise.scala 50:65:@6460.4]
  wire  _T_6426; // @[Bitwise.scala 50:65:@6461.4]
  wire  _T_6427; // @[Bitwise.scala 50:65:@6462.4]
  wire  _T_6428; // @[Bitwise.scala 50:65:@6463.4]
  wire  _T_6429; // @[Bitwise.scala 50:65:@6464.4]
  wire  _T_6430; // @[Bitwise.scala 50:65:@6465.4]
  wire  _T_6431; // @[Bitwise.scala 50:65:@6466.4]
  wire  _T_6432; // @[Bitwise.scala 50:65:@6467.4]
  wire [1:0] _T_6433; // @[Bitwise.scala 48:55:@6468.4]
  wire [1:0] _T_6434; // @[Bitwise.scala 48:55:@6469.4]
  wire [1:0] _GEN_749; // @[Bitwise.scala 48:55:@6470.4]
  wire [2:0] _T_6435; // @[Bitwise.scala 48:55:@6470.4]
  wire [2:0] _GEN_750; // @[Bitwise.scala 48:55:@6471.4]
  wire [3:0] _T_6436; // @[Bitwise.scala 48:55:@6471.4]
  wire [1:0] _T_6437; // @[Bitwise.scala 48:55:@6472.4]
  wire [1:0] _T_6438; // @[Bitwise.scala 48:55:@6473.4]
  wire [1:0] _GEN_751; // @[Bitwise.scala 48:55:@6474.4]
  wire [2:0] _T_6439; // @[Bitwise.scala 48:55:@6474.4]
  wire [2:0] _GEN_752; // @[Bitwise.scala 48:55:@6475.4]
  wire [3:0] _T_6440; // @[Bitwise.scala 48:55:@6475.4]
  wire [4:0] _T_6441; // @[Bitwise.scala 48:55:@6476.4]
  wire [1:0] _T_6442; // @[Bitwise.scala 48:55:@6477.4]
  wire [1:0] _T_6443; // @[Bitwise.scala 48:55:@6478.4]
  wire [1:0] _GEN_753; // @[Bitwise.scala 48:55:@6479.4]
  wire [2:0] _T_6444; // @[Bitwise.scala 48:55:@6479.4]
  wire [2:0] _GEN_754; // @[Bitwise.scala 48:55:@6480.4]
  wire [3:0] _T_6445; // @[Bitwise.scala 48:55:@6480.4]
  wire [1:0] _T_6446; // @[Bitwise.scala 48:55:@6481.4]
  wire [1:0] _T_6447; // @[Bitwise.scala 48:55:@6482.4]
  wire [1:0] _GEN_755; // @[Bitwise.scala 48:55:@6483.4]
  wire [2:0] _T_6448; // @[Bitwise.scala 48:55:@6483.4]
  wire [2:0] _GEN_756; // @[Bitwise.scala 48:55:@6484.4]
  wire [3:0] _T_6449; // @[Bitwise.scala 48:55:@6484.4]
  wire [4:0] _T_6450; // @[Bitwise.scala 48:55:@6485.4]
  wire [5:0] _T_6451; // @[Bitwise.scala 48:55:@6486.4]
  wire [1:0] _T_6452; // @[Bitwise.scala 48:55:@6487.4]
  wire [1:0] _T_6453; // @[Bitwise.scala 48:55:@6488.4]
  wire [1:0] _GEN_757; // @[Bitwise.scala 48:55:@6489.4]
  wire [2:0] _T_6454; // @[Bitwise.scala 48:55:@6489.4]
  wire [2:0] _GEN_758; // @[Bitwise.scala 48:55:@6490.4]
  wire [3:0] _T_6455; // @[Bitwise.scala 48:55:@6490.4]
  wire [1:0] _T_6456; // @[Bitwise.scala 48:55:@6491.4]
  wire [1:0] _T_6457; // @[Bitwise.scala 48:55:@6492.4]
  wire [1:0] _GEN_759; // @[Bitwise.scala 48:55:@6493.4]
  wire [2:0] _T_6458; // @[Bitwise.scala 48:55:@6493.4]
  wire [2:0] _GEN_760; // @[Bitwise.scala 48:55:@6494.4]
  wire [3:0] _T_6459; // @[Bitwise.scala 48:55:@6494.4]
  wire [4:0] _T_6460; // @[Bitwise.scala 48:55:@6495.4]
  wire [1:0] _T_6461; // @[Bitwise.scala 48:55:@6496.4]
  wire [1:0] _T_6462; // @[Bitwise.scala 48:55:@6497.4]
  wire [1:0] _GEN_761; // @[Bitwise.scala 48:55:@6498.4]
  wire [2:0] _T_6463; // @[Bitwise.scala 48:55:@6498.4]
  wire [2:0] _GEN_762; // @[Bitwise.scala 48:55:@6499.4]
  wire [3:0] _T_6464; // @[Bitwise.scala 48:55:@6499.4]
  wire [1:0] _T_6465; // @[Bitwise.scala 48:55:@6500.4]
  wire [1:0] _GEN_763; // @[Bitwise.scala 48:55:@6501.4]
  wire [2:0] _T_6466; // @[Bitwise.scala 48:55:@6501.4]
  wire [1:0] _T_6467; // @[Bitwise.scala 48:55:@6502.4]
  wire [1:0] _GEN_764; // @[Bitwise.scala 48:55:@6503.4]
  wire [2:0] _T_6468; // @[Bitwise.scala 48:55:@6503.4]
  wire [3:0] _T_6469; // @[Bitwise.scala 48:55:@6504.4]
  wire [4:0] _T_6470; // @[Bitwise.scala 48:55:@6505.4]
  wire [5:0] _T_6471; // @[Bitwise.scala 48:55:@6506.4]
  wire [6:0] _T_6472; // @[Bitwise.scala 48:55:@6507.4]
  wire [41:0] _T_6536; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6572.4]
  wire  _T_6537; // @[Bitwise.scala 50:65:@6573.4]
  wire  _T_6538; // @[Bitwise.scala 50:65:@6574.4]
  wire  _T_6539; // @[Bitwise.scala 50:65:@6575.4]
  wire  _T_6540; // @[Bitwise.scala 50:65:@6576.4]
  wire  _T_6541; // @[Bitwise.scala 50:65:@6577.4]
  wire  _T_6542; // @[Bitwise.scala 50:65:@6578.4]
  wire  _T_6543; // @[Bitwise.scala 50:65:@6579.4]
  wire  _T_6544; // @[Bitwise.scala 50:65:@6580.4]
  wire  _T_6545; // @[Bitwise.scala 50:65:@6581.4]
  wire  _T_6546; // @[Bitwise.scala 50:65:@6582.4]
  wire  _T_6547; // @[Bitwise.scala 50:65:@6583.4]
  wire  _T_6548; // @[Bitwise.scala 50:65:@6584.4]
  wire  _T_6549; // @[Bitwise.scala 50:65:@6585.4]
  wire  _T_6550; // @[Bitwise.scala 50:65:@6586.4]
  wire  _T_6551; // @[Bitwise.scala 50:65:@6587.4]
  wire  _T_6552; // @[Bitwise.scala 50:65:@6588.4]
  wire  _T_6553; // @[Bitwise.scala 50:65:@6589.4]
  wire  _T_6554; // @[Bitwise.scala 50:65:@6590.4]
  wire  _T_6555; // @[Bitwise.scala 50:65:@6591.4]
  wire  _T_6556; // @[Bitwise.scala 50:65:@6592.4]
  wire  _T_6557; // @[Bitwise.scala 50:65:@6593.4]
  wire  _T_6558; // @[Bitwise.scala 50:65:@6594.4]
  wire  _T_6559; // @[Bitwise.scala 50:65:@6595.4]
  wire  _T_6560; // @[Bitwise.scala 50:65:@6596.4]
  wire  _T_6561; // @[Bitwise.scala 50:65:@6597.4]
  wire  _T_6562; // @[Bitwise.scala 50:65:@6598.4]
  wire  _T_6563; // @[Bitwise.scala 50:65:@6599.4]
  wire  _T_6564; // @[Bitwise.scala 50:65:@6600.4]
  wire  _T_6565; // @[Bitwise.scala 50:65:@6601.4]
  wire  _T_6566; // @[Bitwise.scala 50:65:@6602.4]
  wire  _T_6567; // @[Bitwise.scala 50:65:@6603.4]
  wire  _T_6568; // @[Bitwise.scala 50:65:@6604.4]
  wire  _T_6569; // @[Bitwise.scala 50:65:@6605.4]
  wire  _T_6570; // @[Bitwise.scala 50:65:@6606.4]
  wire  _T_6571; // @[Bitwise.scala 50:65:@6607.4]
  wire  _T_6572; // @[Bitwise.scala 50:65:@6608.4]
  wire  _T_6573; // @[Bitwise.scala 50:65:@6609.4]
  wire  _T_6574; // @[Bitwise.scala 50:65:@6610.4]
  wire  _T_6575; // @[Bitwise.scala 50:65:@6611.4]
  wire  _T_6576; // @[Bitwise.scala 50:65:@6612.4]
  wire  _T_6577; // @[Bitwise.scala 50:65:@6613.4]
  wire  _T_6578; // @[Bitwise.scala 50:65:@6614.4]
  wire [1:0] _T_6579; // @[Bitwise.scala 48:55:@6615.4]
  wire [1:0] _T_6580; // @[Bitwise.scala 48:55:@6616.4]
  wire [1:0] _GEN_765; // @[Bitwise.scala 48:55:@6617.4]
  wire [2:0] _T_6581; // @[Bitwise.scala 48:55:@6617.4]
  wire [2:0] _GEN_766; // @[Bitwise.scala 48:55:@6618.4]
  wire [3:0] _T_6582; // @[Bitwise.scala 48:55:@6618.4]
  wire [1:0] _T_6583; // @[Bitwise.scala 48:55:@6619.4]
  wire [1:0] _T_6584; // @[Bitwise.scala 48:55:@6620.4]
  wire [1:0] _GEN_767; // @[Bitwise.scala 48:55:@6621.4]
  wire [2:0] _T_6585; // @[Bitwise.scala 48:55:@6621.4]
  wire [2:0] _GEN_768; // @[Bitwise.scala 48:55:@6622.4]
  wire [3:0] _T_6586; // @[Bitwise.scala 48:55:@6622.4]
  wire [4:0] _T_6587; // @[Bitwise.scala 48:55:@6623.4]
  wire [1:0] _T_6588; // @[Bitwise.scala 48:55:@6624.4]
  wire [1:0] _T_6589; // @[Bitwise.scala 48:55:@6625.4]
  wire [1:0] _GEN_769; // @[Bitwise.scala 48:55:@6626.4]
  wire [2:0] _T_6590; // @[Bitwise.scala 48:55:@6626.4]
  wire [2:0] _GEN_770; // @[Bitwise.scala 48:55:@6627.4]
  wire [3:0] _T_6591; // @[Bitwise.scala 48:55:@6627.4]
  wire [1:0] _T_6592; // @[Bitwise.scala 48:55:@6628.4]
  wire [1:0] _GEN_771; // @[Bitwise.scala 48:55:@6629.4]
  wire [2:0] _T_6593; // @[Bitwise.scala 48:55:@6629.4]
  wire [1:0] _T_6594; // @[Bitwise.scala 48:55:@6630.4]
  wire [1:0] _GEN_772; // @[Bitwise.scala 48:55:@6631.4]
  wire [2:0] _T_6595; // @[Bitwise.scala 48:55:@6631.4]
  wire [3:0] _T_6596; // @[Bitwise.scala 48:55:@6632.4]
  wire [4:0] _T_6597; // @[Bitwise.scala 48:55:@6633.4]
  wire [5:0] _T_6598; // @[Bitwise.scala 48:55:@6634.4]
  wire [1:0] _T_6599; // @[Bitwise.scala 48:55:@6635.4]
  wire [1:0] _T_6600; // @[Bitwise.scala 48:55:@6636.4]
  wire [1:0] _GEN_773; // @[Bitwise.scala 48:55:@6637.4]
  wire [2:0] _T_6601; // @[Bitwise.scala 48:55:@6637.4]
  wire [2:0] _GEN_774; // @[Bitwise.scala 48:55:@6638.4]
  wire [3:0] _T_6602; // @[Bitwise.scala 48:55:@6638.4]
  wire [1:0] _T_6603; // @[Bitwise.scala 48:55:@6639.4]
  wire [1:0] _T_6604; // @[Bitwise.scala 48:55:@6640.4]
  wire [1:0] _GEN_775; // @[Bitwise.scala 48:55:@6641.4]
  wire [2:0] _T_6605; // @[Bitwise.scala 48:55:@6641.4]
  wire [2:0] _GEN_776; // @[Bitwise.scala 48:55:@6642.4]
  wire [3:0] _T_6606; // @[Bitwise.scala 48:55:@6642.4]
  wire [4:0] _T_6607; // @[Bitwise.scala 48:55:@6643.4]
  wire [1:0] _T_6608; // @[Bitwise.scala 48:55:@6644.4]
  wire [1:0] _T_6609; // @[Bitwise.scala 48:55:@6645.4]
  wire [1:0] _GEN_777; // @[Bitwise.scala 48:55:@6646.4]
  wire [2:0] _T_6610; // @[Bitwise.scala 48:55:@6646.4]
  wire [2:0] _GEN_778; // @[Bitwise.scala 48:55:@6647.4]
  wire [3:0] _T_6611; // @[Bitwise.scala 48:55:@6647.4]
  wire [1:0] _T_6612; // @[Bitwise.scala 48:55:@6648.4]
  wire [1:0] _GEN_779; // @[Bitwise.scala 48:55:@6649.4]
  wire [2:0] _T_6613; // @[Bitwise.scala 48:55:@6649.4]
  wire [1:0] _T_6614; // @[Bitwise.scala 48:55:@6650.4]
  wire [1:0] _GEN_780; // @[Bitwise.scala 48:55:@6651.4]
  wire [2:0] _T_6615; // @[Bitwise.scala 48:55:@6651.4]
  wire [3:0] _T_6616; // @[Bitwise.scala 48:55:@6652.4]
  wire [4:0] _T_6617; // @[Bitwise.scala 48:55:@6653.4]
  wire [5:0] _T_6618; // @[Bitwise.scala 48:55:@6654.4]
  wire [6:0] _T_6619; // @[Bitwise.scala 48:55:@6655.4]
  wire [42:0] _T_6683; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6720.4]
  wire  _T_6684; // @[Bitwise.scala 50:65:@6721.4]
  wire  _T_6685; // @[Bitwise.scala 50:65:@6722.4]
  wire  _T_6686; // @[Bitwise.scala 50:65:@6723.4]
  wire  _T_6687; // @[Bitwise.scala 50:65:@6724.4]
  wire  _T_6688; // @[Bitwise.scala 50:65:@6725.4]
  wire  _T_6689; // @[Bitwise.scala 50:65:@6726.4]
  wire  _T_6690; // @[Bitwise.scala 50:65:@6727.4]
  wire  _T_6691; // @[Bitwise.scala 50:65:@6728.4]
  wire  _T_6692; // @[Bitwise.scala 50:65:@6729.4]
  wire  _T_6693; // @[Bitwise.scala 50:65:@6730.4]
  wire  _T_6694; // @[Bitwise.scala 50:65:@6731.4]
  wire  _T_6695; // @[Bitwise.scala 50:65:@6732.4]
  wire  _T_6696; // @[Bitwise.scala 50:65:@6733.4]
  wire  _T_6697; // @[Bitwise.scala 50:65:@6734.4]
  wire  _T_6698; // @[Bitwise.scala 50:65:@6735.4]
  wire  _T_6699; // @[Bitwise.scala 50:65:@6736.4]
  wire  _T_6700; // @[Bitwise.scala 50:65:@6737.4]
  wire  _T_6701; // @[Bitwise.scala 50:65:@6738.4]
  wire  _T_6702; // @[Bitwise.scala 50:65:@6739.4]
  wire  _T_6703; // @[Bitwise.scala 50:65:@6740.4]
  wire  _T_6704; // @[Bitwise.scala 50:65:@6741.4]
  wire  _T_6705; // @[Bitwise.scala 50:65:@6742.4]
  wire  _T_6706; // @[Bitwise.scala 50:65:@6743.4]
  wire  _T_6707; // @[Bitwise.scala 50:65:@6744.4]
  wire  _T_6708; // @[Bitwise.scala 50:65:@6745.4]
  wire  _T_6709; // @[Bitwise.scala 50:65:@6746.4]
  wire  _T_6710; // @[Bitwise.scala 50:65:@6747.4]
  wire  _T_6711; // @[Bitwise.scala 50:65:@6748.4]
  wire  _T_6712; // @[Bitwise.scala 50:65:@6749.4]
  wire  _T_6713; // @[Bitwise.scala 50:65:@6750.4]
  wire  _T_6714; // @[Bitwise.scala 50:65:@6751.4]
  wire  _T_6715; // @[Bitwise.scala 50:65:@6752.4]
  wire  _T_6716; // @[Bitwise.scala 50:65:@6753.4]
  wire  _T_6717; // @[Bitwise.scala 50:65:@6754.4]
  wire  _T_6718; // @[Bitwise.scala 50:65:@6755.4]
  wire  _T_6719; // @[Bitwise.scala 50:65:@6756.4]
  wire  _T_6720; // @[Bitwise.scala 50:65:@6757.4]
  wire  _T_6721; // @[Bitwise.scala 50:65:@6758.4]
  wire  _T_6722; // @[Bitwise.scala 50:65:@6759.4]
  wire  _T_6723; // @[Bitwise.scala 50:65:@6760.4]
  wire  _T_6724; // @[Bitwise.scala 50:65:@6761.4]
  wire  _T_6725; // @[Bitwise.scala 50:65:@6762.4]
  wire  _T_6726; // @[Bitwise.scala 50:65:@6763.4]
  wire [1:0] _T_6727; // @[Bitwise.scala 48:55:@6764.4]
  wire [1:0] _T_6728; // @[Bitwise.scala 48:55:@6765.4]
  wire [1:0] _GEN_781; // @[Bitwise.scala 48:55:@6766.4]
  wire [2:0] _T_6729; // @[Bitwise.scala 48:55:@6766.4]
  wire [2:0] _GEN_782; // @[Bitwise.scala 48:55:@6767.4]
  wire [3:0] _T_6730; // @[Bitwise.scala 48:55:@6767.4]
  wire [1:0] _T_6731; // @[Bitwise.scala 48:55:@6768.4]
  wire [1:0] _T_6732; // @[Bitwise.scala 48:55:@6769.4]
  wire [1:0] _GEN_783; // @[Bitwise.scala 48:55:@6770.4]
  wire [2:0] _T_6733; // @[Bitwise.scala 48:55:@6770.4]
  wire [2:0] _GEN_784; // @[Bitwise.scala 48:55:@6771.4]
  wire [3:0] _T_6734; // @[Bitwise.scala 48:55:@6771.4]
  wire [4:0] _T_6735; // @[Bitwise.scala 48:55:@6772.4]
  wire [1:0] _T_6736; // @[Bitwise.scala 48:55:@6773.4]
  wire [1:0] _T_6737; // @[Bitwise.scala 48:55:@6774.4]
  wire [1:0] _GEN_785; // @[Bitwise.scala 48:55:@6775.4]
  wire [2:0] _T_6738; // @[Bitwise.scala 48:55:@6775.4]
  wire [2:0] _GEN_786; // @[Bitwise.scala 48:55:@6776.4]
  wire [3:0] _T_6739; // @[Bitwise.scala 48:55:@6776.4]
  wire [1:0] _T_6740; // @[Bitwise.scala 48:55:@6777.4]
  wire [1:0] _GEN_787; // @[Bitwise.scala 48:55:@6778.4]
  wire [2:0] _T_6741; // @[Bitwise.scala 48:55:@6778.4]
  wire [1:0] _T_6742; // @[Bitwise.scala 48:55:@6779.4]
  wire [1:0] _GEN_788; // @[Bitwise.scala 48:55:@6780.4]
  wire [2:0] _T_6743; // @[Bitwise.scala 48:55:@6780.4]
  wire [3:0] _T_6744; // @[Bitwise.scala 48:55:@6781.4]
  wire [4:0] _T_6745; // @[Bitwise.scala 48:55:@6782.4]
  wire [5:0] _T_6746; // @[Bitwise.scala 48:55:@6783.4]
  wire [1:0] _T_6747; // @[Bitwise.scala 48:55:@6784.4]
  wire [1:0] _T_6748; // @[Bitwise.scala 48:55:@6785.4]
  wire [1:0] _GEN_789; // @[Bitwise.scala 48:55:@6786.4]
  wire [2:0] _T_6749; // @[Bitwise.scala 48:55:@6786.4]
  wire [2:0] _GEN_790; // @[Bitwise.scala 48:55:@6787.4]
  wire [3:0] _T_6750; // @[Bitwise.scala 48:55:@6787.4]
  wire [1:0] _T_6751; // @[Bitwise.scala 48:55:@6788.4]
  wire [1:0] _GEN_791; // @[Bitwise.scala 48:55:@6789.4]
  wire [2:0] _T_6752; // @[Bitwise.scala 48:55:@6789.4]
  wire [1:0] _T_6753; // @[Bitwise.scala 48:55:@6790.4]
  wire [1:0] _GEN_792; // @[Bitwise.scala 48:55:@6791.4]
  wire [2:0] _T_6754; // @[Bitwise.scala 48:55:@6791.4]
  wire [3:0] _T_6755; // @[Bitwise.scala 48:55:@6792.4]
  wire [4:0] _T_6756; // @[Bitwise.scala 48:55:@6793.4]
  wire [1:0] _T_6757; // @[Bitwise.scala 48:55:@6794.4]
  wire [1:0] _T_6758; // @[Bitwise.scala 48:55:@6795.4]
  wire [1:0] _GEN_793; // @[Bitwise.scala 48:55:@6796.4]
  wire [2:0] _T_6759; // @[Bitwise.scala 48:55:@6796.4]
  wire [2:0] _GEN_794; // @[Bitwise.scala 48:55:@6797.4]
  wire [3:0] _T_6760; // @[Bitwise.scala 48:55:@6797.4]
  wire [1:0] _T_6761; // @[Bitwise.scala 48:55:@6798.4]
  wire [1:0] _GEN_795; // @[Bitwise.scala 48:55:@6799.4]
  wire [2:0] _T_6762; // @[Bitwise.scala 48:55:@6799.4]
  wire [1:0] _T_6763; // @[Bitwise.scala 48:55:@6800.4]
  wire [1:0] _GEN_796; // @[Bitwise.scala 48:55:@6801.4]
  wire [2:0] _T_6764; // @[Bitwise.scala 48:55:@6801.4]
  wire [3:0] _T_6765; // @[Bitwise.scala 48:55:@6802.4]
  wire [4:0] _T_6766; // @[Bitwise.scala 48:55:@6803.4]
  wire [5:0] _T_6767; // @[Bitwise.scala 48:55:@6804.4]
  wire [6:0] _T_6768; // @[Bitwise.scala 48:55:@6805.4]
  wire [43:0] _T_6832; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6870.4]
  wire  _T_6833; // @[Bitwise.scala 50:65:@6871.4]
  wire  _T_6834; // @[Bitwise.scala 50:65:@6872.4]
  wire  _T_6835; // @[Bitwise.scala 50:65:@6873.4]
  wire  _T_6836; // @[Bitwise.scala 50:65:@6874.4]
  wire  _T_6837; // @[Bitwise.scala 50:65:@6875.4]
  wire  _T_6838; // @[Bitwise.scala 50:65:@6876.4]
  wire  _T_6839; // @[Bitwise.scala 50:65:@6877.4]
  wire  _T_6840; // @[Bitwise.scala 50:65:@6878.4]
  wire  _T_6841; // @[Bitwise.scala 50:65:@6879.4]
  wire  _T_6842; // @[Bitwise.scala 50:65:@6880.4]
  wire  _T_6843; // @[Bitwise.scala 50:65:@6881.4]
  wire  _T_6844; // @[Bitwise.scala 50:65:@6882.4]
  wire  _T_6845; // @[Bitwise.scala 50:65:@6883.4]
  wire  _T_6846; // @[Bitwise.scala 50:65:@6884.4]
  wire  _T_6847; // @[Bitwise.scala 50:65:@6885.4]
  wire  _T_6848; // @[Bitwise.scala 50:65:@6886.4]
  wire  _T_6849; // @[Bitwise.scala 50:65:@6887.4]
  wire  _T_6850; // @[Bitwise.scala 50:65:@6888.4]
  wire  _T_6851; // @[Bitwise.scala 50:65:@6889.4]
  wire  _T_6852; // @[Bitwise.scala 50:65:@6890.4]
  wire  _T_6853; // @[Bitwise.scala 50:65:@6891.4]
  wire  _T_6854; // @[Bitwise.scala 50:65:@6892.4]
  wire  _T_6855; // @[Bitwise.scala 50:65:@6893.4]
  wire  _T_6856; // @[Bitwise.scala 50:65:@6894.4]
  wire  _T_6857; // @[Bitwise.scala 50:65:@6895.4]
  wire  _T_6858; // @[Bitwise.scala 50:65:@6896.4]
  wire  _T_6859; // @[Bitwise.scala 50:65:@6897.4]
  wire  _T_6860; // @[Bitwise.scala 50:65:@6898.4]
  wire  _T_6861; // @[Bitwise.scala 50:65:@6899.4]
  wire  _T_6862; // @[Bitwise.scala 50:65:@6900.4]
  wire  _T_6863; // @[Bitwise.scala 50:65:@6901.4]
  wire  _T_6864; // @[Bitwise.scala 50:65:@6902.4]
  wire  _T_6865; // @[Bitwise.scala 50:65:@6903.4]
  wire  _T_6866; // @[Bitwise.scala 50:65:@6904.4]
  wire  _T_6867; // @[Bitwise.scala 50:65:@6905.4]
  wire  _T_6868; // @[Bitwise.scala 50:65:@6906.4]
  wire  _T_6869; // @[Bitwise.scala 50:65:@6907.4]
  wire  _T_6870; // @[Bitwise.scala 50:65:@6908.4]
  wire  _T_6871; // @[Bitwise.scala 50:65:@6909.4]
  wire  _T_6872; // @[Bitwise.scala 50:65:@6910.4]
  wire  _T_6873; // @[Bitwise.scala 50:65:@6911.4]
  wire  _T_6874; // @[Bitwise.scala 50:65:@6912.4]
  wire  _T_6875; // @[Bitwise.scala 50:65:@6913.4]
  wire  _T_6876; // @[Bitwise.scala 50:65:@6914.4]
  wire [1:0] _T_6877; // @[Bitwise.scala 48:55:@6915.4]
  wire [1:0] _T_6878; // @[Bitwise.scala 48:55:@6916.4]
  wire [1:0] _GEN_797; // @[Bitwise.scala 48:55:@6917.4]
  wire [2:0] _T_6879; // @[Bitwise.scala 48:55:@6917.4]
  wire [2:0] _GEN_798; // @[Bitwise.scala 48:55:@6918.4]
  wire [3:0] _T_6880; // @[Bitwise.scala 48:55:@6918.4]
  wire [1:0] _T_6881; // @[Bitwise.scala 48:55:@6919.4]
  wire [1:0] _GEN_799; // @[Bitwise.scala 48:55:@6920.4]
  wire [2:0] _T_6882; // @[Bitwise.scala 48:55:@6920.4]
  wire [1:0] _T_6883; // @[Bitwise.scala 48:55:@6921.4]
  wire [1:0] _GEN_800; // @[Bitwise.scala 48:55:@6922.4]
  wire [2:0] _T_6884; // @[Bitwise.scala 48:55:@6922.4]
  wire [3:0] _T_6885; // @[Bitwise.scala 48:55:@6923.4]
  wire [4:0] _T_6886; // @[Bitwise.scala 48:55:@6924.4]
  wire [1:0] _T_6887; // @[Bitwise.scala 48:55:@6925.4]
  wire [1:0] _T_6888; // @[Bitwise.scala 48:55:@6926.4]
  wire [1:0] _GEN_801; // @[Bitwise.scala 48:55:@6927.4]
  wire [2:0] _T_6889; // @[Bitwise.scala 48:55:@6927.4]
  wire [2:0] _GEN_802; // @[Bitwise.scala 48:55:@6928.4]
  wire [3:0] _T_6890; // @[Bitwise.scala 48:55:@6928.4]
  wire [1:0] _T_6891; // @[Bitwise.scala 48:55:@6929.4]
  wire [1:0] _GEN_803; // @[Bitwise.scala 48:55:@6930.4]
  wire [2:0] _T_6892; // @[Bitwise.scala 48:55:@6930.4]
  wire [1:0] _T_6893; // @[Bitwise.scala 48:55:@6931.4]
  wire [1:0] _GEN_804; // @[Bitwise.scala 48:55:@6932.4]
  wire [2:0] _T_6894; // @[Bitwise.scala 48:55:@6932.4]
  wire [3:0] _T_6895; // @[Bitwise.scala 48:55:@6933.4]
  wire [4:0] _T_6896; // @[Bitwise.scala 48:55:@6934.4]
  wire [5:0] _T_6897; // @[Bitwise.scala 48:55:@6935.4]
  wire [1:0] _T_6898; // @[Bitwise.scala 48:55:@6936.4]
  wire [1:0] _T_6899; // @[Bitwise.scala 48:55:@6937.4]
  wire [1:0] _GEN_805; // @[Bitwise.scala 48:55:@6938.4]
  wire [2:0] _T_6900; // @[Bitwise.scala 48:55:@6938.4]
  wire [2:0] _GEN_806; // @[Bitwise.scala 48:55:@6939.4]
  wire [3:0] _T_6901; // @[Bitwise.scala 48:55:@6939.4]
  wire [1:0] _T_6902; // @[Bitwise.scala 48:55:@6940.4]
  wire [1:0] _GEN_807; // @[Bitwise.scala 48:55:@6941.4]
  wire [2:0] _T_6903; // @[Bitwise.scala 48:55:@6941.4]
  wire [1:0] _T_6904; // @[Bitwise.scala 48:55:@6942.4]
  wire [1:0] _GEN_808; // @[Bitwise.scala 48:55:@6943.4]
  wire [2:0] _T_6905; // @[Bitwise.scala 48:55:@6943.4]
  wire [3:0] _T_6906; // @[Bitwise.scala 48:55:@6944.4]
  wire [4:0] _T_6907; // @[Bitwise.scala 48:55:@6945.4]
  wire [1:0] _T_6908; // @[Bitwise.scala 48:55:@6946.4]
  wire [1:0] _T_6909; // @[Bitwise.scala 48:55:@6947.4]
  wire [1:0] _GEN_809; // @[Bitwise.scala 48:55:@6948.4]
  wire [2:0] _T_6910; // @[Bitwise.scala 48:55:@6948.4]
  wire [2:0] _GEN_810; // @[Bitwise.scala 48:55:@6949.4]
  wire [3:0] _T_6911; // @[Bitwise.scala 48:55:@6949.4]
  wire [1:0] _T_6912; // @[Bitwise.scala 48:55:@6950.4]
  wire [1:0] _GEN_811; // @[Bitwise.scala 48:55:@6951.4]
  wire [2:0] _T_6913; // @[Bitwise.scala 48:55:@6951.4]
  wire [1:0] _T_6914; // @[Bitwise.scala 48:55:@6952.4]
  wire [1:0] _GEN_812; // @[Bitwise.scala 48:55:@6953.4]
  wire [2:0] _T_6915; // @[Bitwise.scala 48:55:@6953.4]
  wire [3:0] _T_6916; // @[Bitwise.scala 48:55:@6954.4]
  wire [4:0] _T_6917; // @[Bitwise.scala 48:55:@6955.4]
  wire [5:0] _T_6918; // @[Bitwise.scala 48:55:@6956.4]
  wire [6:0] _T_6919; // @[Bitwise.scala 48:55:@6957.4]
  wire [44:0] _T_6983; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7022.4]
  wire  _T_6984; // @[Bitwise.scala 50:65:@7023.4]
  wire  _T_6985; // @[Bitwise.scala 50:65:@7024.4]
  wire  _T_6986; // @[Bitwise.scala 50:65:@7025.4]
  wire  _T_6987; // @[Bitwise.scala 50:65:@7026.4]
  wire  _T_6988; // @[Bitwise.scala 50:65:@7027.4]
  wire  _T_6989; // @[Bitwise.scala 50:65:@7028.4]
  wire  _T_6990; // @[Bitwise.scala 50:65:@7029.4]
  wire  _T_6991; // @[Bitwise.scala 50:65:@7030.4]
  wire  _T_6992; // @[Bitwise.scala 50:65:@7031.4]
  wire  _T_6993; // @[Bitwise.scala 50:65:@7032.4]
  wire  _T_6994; // @[Bitwise.scala 50:65:@7033.4]
  wire  _T_6995; // @[Bitwise.scala 50:65:@7034.4]
  wire  _T_6996; // @[Bitwise.scala 50:65:@7035.4]
  wire  _T_6997; // @[Bitwise.scala 50:65:@7036.4]
  wire  _T_6998; // @[Bitwise.scala 50:65:@7037.4]
  wire  _T_6999; // @[Bitwise.scala 50:65:@7038.4]
  wire  _T_7000; // @[Bitwise.scala 50:65:@7039.4]
  wire  _T_7001; // @[Bitwise.scala 50:65:@7040.4]
  wire  _T_7002; // @[Bitwise.scala 50:65:@7041.4]
  wire  _T_7003; // @[Bitwise.scala 50:65:@7042.4]
  wire  _T_7004; // @[Bitwise.scala 50:65:@7043.4]
  wire  _T_7005; // @[Bitwise.scala 50:65:@7044.4]
  wire  _T_7006; // @[Bitwise.scala 50:65:@7045.4]
  wire  _T_7007; // @[Bitwise.scala 50:65:@7046.4]
  wire  _T_7008; // @[Bitwise.scala 50:65:@7047.4]
  wire  _T_7009; // @[Bitwise.scala 50:65:@7048.4]
  wire  _T_7010; // @[Bitwise.scala 50:65:@7049.4]
  wire  _T_7011; // @[Bitwise.scala 50:65:@7050.4]
  wire  _T_7012; // @[Bitwise.scala 50:65:@7051.4]
  wire  _T_7013; // @[Bitwise.scala 50:65:@7052.4]
  wire  _T_7014; // @[Bitwise.scala 50:65:@7053.4]
  wire  _T_7015; // @[Bitwise.scala 50:65:@7054.4]
  wire  _T_7016; // @[Bitwise.scala 50:65:@7055.4]
  wire  _T_7017; // @[Bitwise.scala 50:65:@7056.4]
  wire  _T_7018; // @[Bitwise.scala 50:65:@7057.4]
  wire  _T_7019; // @[Bitwise.scala 50:65:@7058.4]
  wire  _T_7020; // @[Bitwise.scala 50:65:@7059.4]
  wire  _T_7021; // @[Bitwise.scala 50:65:@7060.4]
  wire  _T_7022; // @[Bitwise.scala 50:65:@7061.4]
  wire  _T_7023; // @[Bitwise.scala 50:65:@7062.4]
  wire  _T_7024; // @[Bitwise.scala 50:65:@7063.4]
  wire  _T_7025; // @[Bitwise.scala 50:65:@7064.4]
  wire  _T_7026; // @[Bitwise.scala 50:65:@7065.4]
  wire  _T_7027; // @[Bitwise.scala 50:65:@7066.4]
  wire  _T_7028; // @[Bitwise.scala 50:65:@7067.4]
  wire [1:0] _T_7029; // @[Bitwise.scala 48:55:@7068.4]
  wire [1:0] _T_7030; // @[Bitwise.scala 48:55:@7069.4]
  wire [1:0] _GEN_813; // @[Bitwise.scala 48:55:@7070.4]
  wire [2:0] _T_7031; // @[Bitwise.scala 48:55:@7070.4]
  wire [2:0] _GEN_814; // @[Bitwise.scala 48:55:@7071.4]
  wire [3:0] _T_7032; // @[Bitwise.scala 48:55:@7071.4]
  wire [1:0] _T_7033; // @[Bitwise.scala 48:55:@7072.4]
  wire [1:0] _GEN_815; // @[Bitwise.scala 48:55:@7073.4]
  wire [2:0] _T_7034; // @[Bitwise.scala 48:55:@7073.4]
  wire [1:0] _T_7035; // @[Bitwise.scala 48:55:@7074.4]
  wire [1:0] _GEN_816; // @[Bitwise.scala 48:55:@7075.4]
  wire [2:0] _T_7036; // @[Bitwise.scala 48:55:@7075.4]
  wire [3:0] _T_7037; // @[Bitwise.scala 48:55:@7076.4]
  wire [4:0] _T_7038; // @[Bitwise.scala 48:55:@7077.4]
  wire [1:0] _T_7039; // @[Bitwise.scala 48:55:@7078.4]
  wire [1:0] _T_7040; // @[Bitwise.scala 48:55:@7079.4]
  wire [1:0] _GEN_817; // @[Bitwise.scala 48:55:@7080.4]
  wire [2:0] _T_7041; // @[Bitwise.scala 48:55:@7080.4]
  wire [2:0] _GEN_818; // @[Bitwise.scala 48:55:@7081.4]
  wire [3:0] _T_7042; // @[Bitwise.scala 48:55:@7081.4]
  wire [1:0] _T_7043; // @[Bitwise.scala 48:55:@7082.4]
  wire [1:0] _GEN_819; // @[Bitwise.scala 48:55:@7083.4]
  wire [2:0] _T_7044; // @[Bitwise.scala 48:55:@7083.4]
  wire [1:0] _T_7045; // @[Bitwise.scala 48:55:@7084.4]
  wire [1:0] _GEN_820; // @[Bitwise.scala 48:55:@7085.4]
  wire [2:0] _T_7046; // @[Bitwise.scala 48:55:@7085.4]
  wire [3:0] _T_7047; // @[Bitwise.scala 48:55:@7086.4]
  wire [4:0] _T_7048; // @[Bitwise.scala 48:55:@7087.4]
  wire [5:0] _T_7049; // @[Bitwise.scala 48:55:@7088.4]
  wire [1:0] _T_7050; // @[Bitwise.scala 48:55:@7089.4]
  wire [1:0] _T_7051; // @[Bitwise.scala 48:55:@7090.4]
  wire [1:0] _GEN_821; // @[Bitwise.scala 48:55:@7091.4]
  wire [2:0] _T_7052; // @[Bitwise.scala 48:55:@7091.4]
  wire [2:0] _GEN_822; // @[Bitwise.scala 48:55:@7092.4]
  wire [3:0] _T_7053; // @[Bitwise.scala 48:55:@7092.4]
  wire [1:0] _T_7054; // @[Bitwise.scala 48:55:@7093.4]
  wire [1:0] _GEN_823; // @[Bitwise.scala 48:55:@7094.4]
  wire [2:0] _T_7055; // @[Bitwise.scala 48:55:@7094.4]
  wire [1:0] _T_7056; // @[Bitwise.scala 48:55:@7095.4]
  wire [1:0] _GEN_824; // @[Bitwise.scala 48:55:@7096.4]
  wire [2:0] _T_7057; // @[Bitwise.scala 48:55:@7096.4]
  wire [3:0] _T_7058; // @[Bitwise.scala 48:55:@7097.4]
  wire [4:0] _T_7059; // @[Bitwise.scala 48:55:@7098.4]
  wire [1:0] _T_7060; // @[Bitwise.scala 48:55:@7099.4]
  wire [1:0] _GEN_825; // @[Bitwise.scala 48:55:@7100.4]
  wire [2:0] _T_7061; // @[Bitwise.scala 48:55:@7100.4]
  wire [1:0] _T_7062; // @[Bitwise.scala 48:55:@7101.4]
  wire [1:0] _GEN_826; // @[Bitwise.scala 48:55:@7102.4]
  wire [2:0] _T_7063; // @[Bitwise.scala 48:55:@7102.4]
  wire [3:0] _T_7064; // @[Bitwise.scala 48:55:@7103.4]
  wire [1:0] _T_7065; // @[Bitwise.scala 48:55:@7104.4]
  wire [1:0] _GEN_827; // @[Bitwise.scala 48:55:@7105.4]
  wire [2:0] _T_7066; // @[Bitwise.scala 48:55:@7105.4]
  wire [1:0] _T_7067; // @[Bitwise.scala 48:55:@7106.4]
  wire [1:0] _GEN_828; // @[Bitwise.scala 48:55:@7107.4]
  wire [2:0] _T_7068; // @[Bitwise.scala 48:55:@7107.4]
  wire [3:0] _T_7069; // @[Bitwise.scala 48:55:@7108.4]
  wire [4:0] _T_7070; // @[Bitwise.scala 48:55:@7109.4]
  wire [5:0] _T_7071; // @[Bitwise.scala 48:55:@7110.4]
  wire [6:0] _T_7072; // @[Bitwise.scala 48:55:@7111.4]
  wire [45:0] _T_7136; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7176.4]
  wire  _T_7137; // @[Bitwise.scala 50:65:@7177.4]
  wire  _T_7138; // @[Bitwise.scala 50:65:@7178.4]
  wire  _T_7139; // @[Bitwise.scala 50:65:@7179.4]
  wire  _T_7140; // @[Bitwise.scala 50:65:@7180.4]
  wire  _T_7141; // @[Bitwise.scala 50:65:@7181.4]
  wire  _T_7142; // @[Bitwise.scala 50:65:@7182.4]
  wire  _T_7143; // @[Bitwise.scala 50:65:@7183.4]
  wire  _T_7144; // @[Bitwise.scala 50:65:@7184.4]
  wire  _T_7145; // @[Bitwise.scala 50:65:@7185.4]
  wire  _T_7146; // @[Bitwise.scala 50:65:@7186.4]
  wire  _T_7147; // @[Bitwise.scala 50:65:@7187.4]
  wire  _T_7148; // @[Bitwise.scala 50:65:@7188.4]
  wire  _T_7149; // @[Bitwise.scala 50:65:@7189.4]
  wire  _T_7150; // @[Bitwise.scala 50:65:@7190.4]
  wire  _T_7151; // @[Bitwise.scala 50:65:@7191.4]
  wire  _T_7152; // @[Bitwise.scala 50:65:@7192.4]
  wire  _T_7153; // @[Bitwise.scala 50:65:@7193.4]
  wire  _T_7154; // @[Bitwise.scala 50:65:@7194.4]
  wire  _T_7155; // @[Bitwise.scala 50:65:@7195.4]
  wire  _T_7156; // @[Bitwise.scala 50:65:@7196.4]
  wire  _T_7157; // @[Bitwise.scala 50:65:@7197.4]
  wire  _T_7158; // @[Bitwise.scala 50:65:@7198.4]
  wire  _T_7159; // @[Bitwise.scala 50:65:@7199.4]
  wire  _T_7160; // @[Bitwise.scala 50:65:@7200.4]
  wire  _T_7161; // @[Bitwise.scala 50:65:@7201.4]
  wire  _T_7162; // @[Bitwise.scala 50:65:@7202.4]
  wire  _T_7163; // @[Bitwise.scala 50:65:@7203.4]
  wire  _T_7164; // @[Bitwise.scala 50:65:@7204.4]
  wire  _T_7165; // @[Bitwise.scala 50:65:@7205.4]
  wire  _T_7166; // @[Bitwise.scala 50:65:@7206.4]
  wire  _T_7167; // @[Bitwise.scala 50:65:@7207.4]
  wire  _T_7168; // @[Bitwise.scala 50:65:@7208.4]
  wire  _T_7169; // @[Bitwise.scala 50:65:@7209.4]
  wire  _T_7170; // @[Bitwise.scala 50:65:@7210.4]
  wire  _T_7171; // @[Bitwise.scala 50:65:@7211.4]
  wire  _T_7172; // @[Bitwise.scala 50:65:@7212.4]
  wire  _T_7173; // @[Bitwise.scala 50:65:@7213.4]
  wire  _T_7174; // @[Bitwise.scala 50:65:@7214.4]
  wire  _T_7175; // @[Bitwise.scala 50:65:@7215.4]
  wire  _T_7176; // @[Bitwise.scala 50:65:@7216.4]
  wire  _T_7177; // @[Bitwise.scala 50:65:@7217.4]
  wire  _T_7178; // @[Bitwise.scala 50:65:@7218.4]
  wire  _T_7179; // @[Bitwise.scala 50:65:@7219.4]
  wire  _T_7180; // @[Bitwise.scala 50:65:@7220.4]
  wire  _T_7181; // @[Bitwise.scala 50:65:@7221.4]
  wire  _T_7182; // @[Bitwise.scala 50:65:@7222.4]
  wire [1:0] _T_7183; // @[Bitwise.scala 48:55:@7223.4]
  wire [1:0] _T_7184; // @[Bitwise.scala 48:55:@7224.4]
  wire [1:0] _GEN_829; // @[Bitwise.scala 48:55:@7225.4]
  wire [2:0] _T_7185; // @[Bitwise.scala 48:55:@7225.4]
  wire [2:0] _GEN_830; // @[Bitwise.scala 48:55:@7226.4]
  wire [3:0] _T_7186; // @[Bitwise.scala 48:55:@7226.4]
  wire [1:0] _T_7187; // @[Bitwise.scala 48:55:@7227.4]
  wire [1:0] _GEN_831; // @[Bitwise.scala 48:55:@7228.4]
  wire [2:0] _T_7188; // @[Bitwise.scala 48:55:@7228.4]
  wire [1:0] _T_7189; // @[Bitwise.scala 48:55:@7229.4]
  wire [1:0] _GEN_832; // @[Bitwise.scala 48:55:@7230.4]
  wire [2:0] _T_7190; // @[Bitwise.scala 48:55:@7230.4]
  wire [3:0] _T_7191; // @[Bitwise.scala 48:55:@7231.4]
  wire [4:0] _T_7192; // @[Bitwise.scala 48:55:@7232.4]
  wire [1:0] _T_7193; // @[Bitwise.scala 48:55:@7233.4]
  wire [1:0] _GEN_833; // @[Bitwise.scala 48:55:@7234.4]
  wire [2:0] _T_7194; // @[Bitwise.scala 48:55:@7234.4]
  wire [1:0] _T_7195; // @[Bitwise.scala 48:55:@7235.4]
  wire [1:0] _GEN_834; // @[Bitwise.scala 48:55:@7236.4]
  wire [2:0] _T_7196; // @[Bitwise.scala 48:55:@7236.4]
  wire [3:0] _T_7197; // @[Bitwise.scala 48:55:@7237.4]
  wire [1:0] _T_7198; // @[Bitwise.scala 48:55:@7238.4]
  wire [1:0] _GEN_835; // @[Bitwise.scala 48:55:@7239.4]
  wire [2:0] _T_7199; // @[Bitwise.scala 48:55:@7239.4]
  wire [1:0] _T_7200; // @[Bitwise.scala 48:55:@7240.4]
  wire [1:0] _GEN_836; // @[Bitwise.scala 48:55:@7241.4]
  wire [2:0] _T_7201; // @[Bitwise.scala 48:55:@7241.4]
  wire [3:0] _T_7202; // @[Bitwise.scala 48:55:@7242.4]
  wire [4:0] _T_7203; // @[Bitwise.scala 48:55:@7243.4]
  wire [5:0] _T_7204; // @[Bitwise.scala 48:55:@7244.4]
  wire [1:0] _T_7205; // @[Bitwise.scala 48:55:@7245.4]
  wire [1:0] _T_7206; // @[Bitwise.scala 48:55:@7246.4]
  wire [1:0] _GEN_837; // @[Bitwise.scala 48:55:@7247.4]
  wire [2:0] _T_7207; // @[Bitwise.scala 48:55:@7247.4]
  wire [2:0] _GEN_838; // @[Bitwise.scala 48:55:@7248.4]
  wire [3:0] _T_7208; // @[Bitwise.scala 48:55:@7248.4]
  wire [1:0] _T_7209; // @[Bitwise.scala 48:55:@7249.4]
  wire [1:0] _GEN_839; // @[Bitwise.scala 48:55:@7250.4]
  wire [2:0] _T_7210; // @[Bitwise.scala 48:55:@7250.4]
  wire [1:0] _T_7211; // @[Bitwise.scala 48:55:@7251.4]
  wire [1:0] _GEN_840; // @[Bitwise.scala 48:55:@7252.4]
  wire [2:0] _T_7212; // @[Bitwise.scala 48:55:@7252.4]
  wire [3:0] _T_7213; // @[Bitwise.scala 48:55:@7253.4]
  wire [4:0] _T_7214; // @[Bitwise.scala 48:55:@7254.4]
  wire [1:0] _T_7215; // @[Bitwise.scala 48:55:@7255.4]
  wire [1:0] _GEN_841; // @[Bitwise.scala 48:55:@7256.4]
  wire [2:0] _T_7216; // @[Bitwise.scala 48:55:@7256.4]
  wire [1:0] _T_7217; // @[Bitwise.scala 48:55:@7257.4]
  wire [1:0] _GEN_842; // @[Bitwise.scala 48:55:@7258.4]
  wire [2:0] _T_7218; // @[Bitwise.scala 48:55:@7258.4]
  wire [3:0] _T_7219; // @[Bitwise.scala 48:55:@7259.4]
  wire [1:0] _T_7220; // @[Bitwise.scala 48:55:@7260.4]
  wire [1:0] _GEN_843; // @[Bitwise.scala 48:55:@7261.4]
  wire [2:0] _T_7221; // @[Bitwise.scala 48:55:@7261.4]
  wire [1:0] _T_7222; // @[Bitwise.scala 48:55:@7262.4]
  wire [1:0] _GEN_844; // @[Bitwise.scala 48:55:@7263.4]
  wire [2:0] _T_7223; // @[Bitwise.scala 48:55:@7263.4]
  wire [3:0] _T_7224; // @[Bitwise.scala 48:55:@7264.4]
  wire [4:0] _T_7225; // @[Bitwise.scala 48:55:@7265.4]
  wire [5:0] _T_7226; // @[Bitwise.scala 48:55:@7266.4]
  wire [6:0] _T_7227; // @[Bitwise.scala 48:55:@7267.4]
  wire [46:0] _T_7291; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7332.4]
  wire  _T_7292; // @[Bitwise.scala 50:65:@7333.4]
  wire  _T_7293; // @[Bitwise.scala 50:65:@7334.4]
  wire  _T_7294; // @[Bitwise.scala 50:65:@7335.4]
  wire  _T_7295; // @[Bitwise.scala 50:65:@7336.4]
  wire  _T_7296; // @[Bitwise.scala 50:65:@7337.4]
  wire  _T_7297; // @[Bitwise.scala 50:65:@7338.4]
  wire  _T_7298; // @[Bitwise.scala 50:65:@7339.4]
  wire  _T_7299; // @[Bitwise.scala 50:65:@7340.4]
  wire  _T_7300; // @[Bitwise.scala 50:65:@7341.4]
  wire  _T_7301; // @[Bitwise.scala 50:65:@7342.4]
  wire  _T_7302; // @[Bitwise.scala 50:65:@7343.4]
  wire  _T_7303; // @[Bitwise.scala 50:65:@7344.4]
  wire  _T_7304; // @[Bitwise.scala 50:65:@7345.4]
  wire  _T_7305; // @[Bitwise.scala 50:65:@7346.4]
  wire  _T_7306; // @[Bitwise.scala 50:65:@7347.4]
  wire  _T_7307; // @[Bitwise.scala 50:65:@7348.4]
  wire  _T_7308; // @[Bitwise.scala 50:65:@7349.4]
  wire  _T_7309; // @[Bitwise.scala 50:65:@7350.4]
  wire  _T_7310; // @[Bitwise.scala 50:65:@7351.4]
  wire  _T_7311; // @[Bitwise.scala 50:65:@7352.4]
  wire  _T_7312; // @[Bitwise.scala 50:65:@7353.4]
  wire  _T_7313; // @[Bitwise.scala 50:65:@7354.4]
  wire  _T_7314; // @[Bitwise.scala 50:65:@7355.4]
  wire  _T_7315; // @[Bitwise.scala 50:65:@7356.4]
  wire  _T_7316; // @[Bitwise.scala 50:65:@7357.4]
  wire  _T_7317; // @[Bitwise.scala 50:65:@7358.4]
  wire  _T_7318; // @[Bitwise.scala 50:65:@7359.4]
  wire  _T_7319; // @[Bitwise.scala 50:65:@7360.4]
  wire  _T_7320; // @[Bitwise.scala 50:65:@7361.4]
  wire  _T_7321; // @[Bitwise.scala 50:65:@7362.4]
  wire  _T_7322; // @[Bitwise.scala 50:65:@7363.4]
  wire  _T_7323; // @[Bitwise.scala 50:65:@7364.4]
  wire  _T_7324; // @[Bitwise.scala 50:65:@7365.4]
  wire  _T_7325; // @[Bitwise.scala 50:65:@7366.4]
  wire  _T_7326; // @[Bitwise.scala 50:65:@7367.4]
  wire  _T_7327; // @[Bitwise.scala 50:65:@7368.4]
  wire  _T_7328; // @[Bitwise.scala 50:65:@7369.4]
  wire  _T_7329; // @[Bitwise.scala 50:65:@7370.4]
  wire  _T_7330; // @[Bitwise.scala 50:65:@7371.4]
  wire  _T_7331; // @[Bitwise.scala 50:65:@7372.4]
  wire  _T_7332; // @[Bitwise.scala 50:65:@7373.4]
  wire  _T_7333; // @[Bitwise.scala 50:65:@7374.4]
  wire  _T_7334; // @[Bitwise.scala 50:65:@7375.4]
  wire  _T_7335; // @[Bitwise.scala 50:65:@7376.4]
  wire  _T_7336; // @[Bitwise.scala 50:65:@7377.4]
  wire  _T_7337; // @[Bitwise.scala 50:65:@7378.4]
  wire  _T_7338; // @[Bitwise.scala 50:65:@7379.4]
  wire [1:0] _T_7339; // @[Bitwise.scala 48:55:@7380.4]
  wire [1:0] _T_7340; // @[Bitwise.scala 48:55:@7381.4]
  wire [1:0] _GEN_845; // @[Bitwise.scala 48:55:@7382.4]
  wire [2:0] _T_7341; // @[Bitwise.scala 48:55:@7382.4]
  wire [2:0] _GEN_846; // @[Bitwise.scala 48:55:@7383.4]
  wire [3:0] _T_7342; // @[Bitwise.scala 48:55:@7383.4]
  wire [1:0] _T_7343; // @[Bitwise.scala 48:55:@7384.4]
  wire [1:0] _GEN_847; // @[Bitwise.scala 48:55:@7385.4]
  wire [2:0] _T_7344; // @[Bitwise.scala 48:55:@7385.4]
  wire [1:0] _T_7345; // @[Bitwise.scala 48:55:@7386.4]
  wire [1:0] _GEN_848; // @[Bitwise.scala 48:55:@7387.4]
  wire [2:0] _T_7346; // @[Bitwise.scala 48:55:@7387.4]
  wire [3:0] _T_7347; // @[Bitwise.scala 48:55:@7388.4]
  wire [4:0] _T_7348; // @[Bitwise.scala 48:55:@7389.4]
  wire [1:0] _T_7349; // @[Bitwise.scala 48:55:@7390.4]
  wire [1:0] _GEN_849; // @[Bitwise.scala 48:55:@7391.4]
  wire [2:0] _T_7350; // @[Bitwise.scala 48:55:@7391.4]
  wire [1:0] _T_7351; // @[Bitwise.scala 48:55:@7392.4]
  wire [1:0] _GEN_850; // @[Bitwise.scala 48:55:@7393.4]
  wire [2:0] _T_7352; // @[Bitwise.scala 48:55:@7393.4]
  wire [3:0] _T_7353; // @[Bitwise.scala 48:55:@7394.4]
  wire [1:0] _T_7354; // @[Bitwise.scala 48:55:@7395.4]
  wire [1:0] _GEN_851; // @[Bitwise.scala 48:55:@7396.4]
  wire [2:0] _T_7355; // @[Bitwise.scala 48:55:@7396.4]
  wire [1:0] _T_7356; // @[Bitwise.scala 48:55:@7397.4]
  wire [1:0] _GEN_852; // @[Bitwise.scala 48:55:@7398.4]
  wire [2:0] _T_7357; // @[Bitwise.scala 48:55:@7398.4]
  wire [3:0] _T_7358; // @[Bitwise.scala 48:55:@7399.4]
  wire [4:0] _T_7359; // @[Bitwise.scala 48:55:@7400.4]
  wire [5:0] _T_7360; // @[Bitwise.scala 48:55:@7401.4]
  wire [1:0] _T_7361; // @[Bitwise.scala 48:55:@7402.4]
  wire [1:0] _GEN_853; // @[Bitwise.scala 48:55:@7403.4]
  wire [2:0] _T_7362; // @[Bitwise.scala 48:55:@7403.4]
  wire [1:0] _T_7363; // @[Bitwise.scala 48:55:@7404.4]
  wire [1:0] _GEN_854; // @[Bitwise.scala 48:55:@7405.4]
  wire [2:0] _T_7364; // @[Bitwise.scala 48:55:@7405.4]
  wire [3:0] _T_7365; // @[Bitwise.scala 48:55:@7406.4]
  wire [1:0] _T_7366; // @[Bitwise.scala 48:55:@7407.4]
  wire [1:0] _GEN_855; // @[Bitwise.scala 48:55:@7408.4]
  wire [2:0] _T_7367; // @[Bitwise.scala 48:55:@7408.4]
  wire [1:0] _T_7368; // @[Bitwise.scala 48:55:@7409.4]
  wire [1:0] _GEN_856; // @[Bitwise.scala 48:55:@7410.4]
  wire [2:0] _T_7369; // @[Bitwise.scala 48:55:@7410.4]
  wire [3:0] _T_7370; // @[Bitwise.scala 48:55:@7411.4]
  wire [4:0] _T_7371; // @[Bitwise.scala 48:55:@7412.4]
  wire [1:0] _T_7372; // @[Bitwise.scala 48:55:@7413.4]
  wire [1:0] _GEN_857; // @[Bitwise.scala 48:55:@7414.4]
  wire [2:0] _T_7373; // @[Bitwise.scala 48:55:@7414.4]
  wire [1:0] _T_7374; // @[Bitwise.scala 48:55:@7415.4]
  wire [1:0] _GEN_858; // @[Bitwise.scala 48:55:@7416.4]
  wire [2:0] _T_7375; // @[Bitwise.scala 48:55:@7416.4]
  wire [3:0] _T_7376; // @[Bitwise.scala 48:55:@7417.4]
  wire [1:0] _T_7377; // @[Bitwise.scala 48:55:@7418.4]
  wire [1:0] _GEN_859; // @[Bitwise.scala 48:55:@7419.4]
  wire [2:0] _T_7378; // @[Bitwise.scala 48:55:@7419.4]
  wire [1:0] _T_7379; // @[Bitwise.scala 48:55:@7420.4]
  wire [1:0] _GEN_860; // @[Bitwise.scala 48:55:@7421.4]
  wire [2:0] _T_7380; // @[Bitwise.scala 48:55:@7421.4]
  wire [3:0] _T_7381; // @[Bitwise.scala 48:55:@7422.4]
  wire [4:0] _T_7382; // @[Bitwise.scala 48:55:@7423.4]
  wire [5:0] _T_7383; // @[Bitwise.scala 48:55:@7424.4]
  wire [6:0] _T_7384; // @[Bitwise.scala 48:55:@7425.4]
  wire [47:0] _T_7448; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7490.4]
  wire  _T_7449; // @[Bitwise.scala 50:65:@7491.4]
  wire  _T_7450; // @[Bitwise.scala 50:65:@7492.4]
  wire  _T_7451; // @[Bitwise.scala 50:65:@7493.4]
  wire  _T_7452; // @[Bitwise.scala 50:65:@7494.4]
  wire  _T_7453; // @[Bitwise.scala 50:65:@7495.4]
  wire  _T_7454; // @[Bitwise.scala 50:65:@7496.4]
  wire  _T_7455; // @[Bitwise.scala 50:65:@7497.4]
  wire  _T_7456; // @[Bitwise.scala 50:65:@7498.4]
  wire  _T_7457; // @[Bitwise.scala 50:65:@7499.4]
  wire  _T_7458; // @[Bitwise.scala 50:65:@7500.4]
  wire  _T_7459; // @[Bitwise.scala 50:65:@7501.4]
  wire  _T_7460; // @[Bitwise.scala 50:65:@7502.4]
  wire  _T_7461; // @[Bitwise.scala 50:65:@7503.4]
  wire  _T_7462; // @[Bitwise.scala 50:65:@7504.4]
  wire  _T_7463; // @[Bitwise.scala 50:65:@7505.4]
  wire  _T_7464; // @[Bitwise.scala 50:65:@7506.4]
  wire  _T_7465; // @[Bitwise.scala 50:65:@7507.4]
  wire  _T_7466; // @[Bitwise.scala 50:65:@7508.4]
  wire  _T_7467; // @[Bitwise.scala 50:65:@7509.4]
  wire  _T_7468; // @[Bitwise.scala 50:65:@7510.4]
  wire  _T_7469; // @[Bitwise.scala 50:65:@7511.4]
  wire  _T_7470; // @[Bitwise.scala 50:65:@7512.4]
  wire  _T_7471; // @[Bitwise.scala 50:65:@7513.4]
  wire  _T_7472; // @[Bitwise.scala 50:65:@7514.4]
  wire  _T_7473; // @[Bitwise.scala 50:65:@7515.4]
  wire  _T_7474; // @[Bitwise.scala 50:65:@7516.4]
  wire  _T_7475; // @[Bitwise.scala 50:65:@7517.4]
  wire  _T_7476; // @[Bitwise.scala 50:65:@7518.4]
  wire  _T_7477; // @[Bitwise.scala 50:65:@7519.4]
  wire  _T_7478; // @[Bitwise.scala 50:65:@7520.4]
  wire  _T_7479; // @[Bitwise.scala 50:65:@7521.4]
  wire  _T_7480; // @[Bitwise.scala 50:65:@7522.4]
  wire  _T_7481; // @[Bitwise.scala 50:65:@7523.4]
  wire  _T_7482; // @[Bitwise.scala 50:65:@7524.4]
  wire  _T_7483; // @[Bitwise.scala 50:65:@7525.4]
  wire  _T_7484; // @[Bitwise.scala 50:65:@7526.4]
  wire  _T_7485; // @[Bitwise.scala 50:65:@7527.4]
  wire  _T_7486; // @[Bitwise.scala 50:65:@7528.4]
  wire  _T_7487; // @[Bitwise.scala 50:65:@7529.4]
  wire  _T_7488; // @[Bitwise.scala 50:65:@7530.4]
  wire  _T_7489; // @[Bitwise.scala 50:65:@7531.4]
  wire  _T_7490; // @[Bitwise.scala 50:65:@7532.4]
  wire  _T_7491; // @[Bitwise.scala 50:65:@7533.4]
  wire  _T_7492; // @[Bitwise.scala 50:65:@7534.4]
  wire  _T_7493; // @[Bitwise.scala 50:65:@7535.4]
  wire  _T_7494; // @[Bitwise.scala 50:65:@7536.4]
  wire  _T_7495; // @[Bitwise.scala 50:65:@7537.4]
  wire  _T_7496; // @[Bitwise.scala 50:65:@7538.4]
  wire [1:0] _T_7497; // @[Bitwise.scala 48:55:@7539.4]
  wire [1:0] _GEN_861; // @[Bitwise.scala 48:55:@7540.4]
  wire [2:0] _T_7498; // @[Bitwise.scala 48:55:@7540.4]
  wire [1:0] _T_7499; // @[Bitwise.scala 48:55:@7541.4]
  wire [1:0] _GEN_862; // @[Bitwise.scala 48:55:@7542.4]
  wire [2:0] _T_7500; // @[Bitwise.scala 48:55:@7542.4]
  wire [3:0] _T_7501; // @[Bitwise.scala 48:55:@7543.4]
  wire [1:0] _T_7502; // @[Bitwise.scala 48:55:@7544.4]
  wire [1:0] _GEN_863; // @[Bitwise.scala 48:55:@7545.4]
  wire [2:0] _T_7503; // @[Bitwise.scala 48:55:@7545.4]
  wire [1:0] _T_7504; // @[Bitwise.scala 48:55:@7546.4]
  wire [1:0] _GEN_864; // @[Bitwise.scala 48:55:@7547.4]
  wire [2:0] _T_7505; // @[Bitwise.scala 48:55:@7547.4]
  wire [3:0] _T_7506; // @[Bitwise.scala 48:55:@7548.4]
  wire [4:0] _T_7507; // @[Bitwise.scala 48:55:@7549.4]
  wire [1:0] _T_7508; // @[Bitwise.scala 48:55:@7550.4]
  wire [1:0] _GEN_865; // @[Bitwise.scala 48:55:@7551.4]
  wire [2:0] _T_7509; // @[Bitwise.scala 48:55:@7551.4]
  wire [1:0] _T_7510; // @[Bitwise.scala 48:55:@7552.4]
  wire [1:0] _GEN_866; // @[Bitwise.scala 48:55:@7553.4]
  wire [2:0] _T_7511; // @[Bitwise.scala 48:55:@7553.4]
  wire [3:0] _T_7512; // @[Bitwise.scala 48:55:@7554.4]
  wire [1:0] _T_7513; // @[Bitwise.scala 48:55:@7555.4]
  wire [1:0] _GEN_867; // @[Bitwise.scala 48:55:@7556.4]
  wire [2:0] _T_7514; // @[Bitwise.scala 48:55:@7556.4]
  wire [1:0] _T_7515; // @[Bitwise.scala 48:55:@7557.4]
  wire [1:0] _GEN_868; // @[Bitwise.scala 48:55:@7558.4]
  wire [2:0] _T_7516; // @[Bitwise.scala 48:55:@7558.4]
  wire [3:0] _T_7517; // @[Bitwise.scala 48:55:@7559.4]
  wire [4:0] _T_7518; // @[Bitwise.scala 48:55:@7560.4]
  wire [5:0] _T_7519; // @[Bitwise.scala 48:55:@7561.4]
  wire [1:0] _T_7520; // @[Bitwise.scala 48:55:@7562.4]
  wire [1:0] _GEN_869; // @[Bitwise.scala 48:55:@7563.4]
  wire [2:0] _T_7521; // @[Bitwise.scala 48:55:@7563.4]
  wire [1:0] _T_7522; // @[Bitwise.scala 48:55:@7564.4]
  wire [1:0] _GEN_870; // @[Bitwise.scala 48:55:@7565.4]
  wire [2:0] _T_7523; // @[Bitwise.scala 48:55:@7565.4]
  wire [3:0] _T_7524; // @[Bitwise.scala 48:55:@7566.4]
  wire [1:0] _T_7525; // @[Bitwise.scala 48:55:@7567.4]
  wire [1:0] _GEN_871; // @[Bitwise.scala 48:55:@7568.4]
  wire [2:0] _T_7526; // @[Bitwise.scala 48:55:@7568.4]
  wire [1:0] _T_7527; // @[Bitwise.scala 48:55:@7569.4]
  wire [1:0] _GEN_872; // @[Bitwise.scala 48:55:@7570.4]
  wire [2:0] _T_7528; // @[Bitwise.scala 48:55:@7570.4]
  wire [3:0] _T_7529; // @[Bitwise.scala 48:55:@7571.4]
  wire [4:0] _T_7530; // @[Bitwise.scala 48:55:@7572.4]
  wire [1:0] _T_7531; // @[Bitwise.scala 48:55:@7573.4]
  wire [1:0] _GEN_873; // @[Bitwise.scala 48:55:@7574.4]
  wire [2:0] _T_7532; // @[Bitwise.scala 48:55:@7574.4]
  wire [1:0] _T_7533; // @[Bitwise.scala 48:55:@7575.4]
  wire [1:0] _GEN_874; // @[Bitwise.scala 48:55:@7576.4]
  wire [2:0] _T_7534; // @[Bitwise.scala 48:55:@7576.4]
  wire [3:0] _T_7535; // @[Bitwise.scala 48:55:@7577.4]
  wire [1:0] _T_7536; // @[Bitwise.scala 48:55:@7578.4]
  wire [1:0] _GEN_875; // @[Bitwise.scala 48:55:@7579.4]
  wire [2:0] _T_7537; // @[Bitwise.scala 48:55:@7579.4]
  wire [1:0] _T_7538; // @[Bitwise.scala 48:55:@7580.4]
  wire [1:0] _GEN_876; // @[Bitwise.scala 48:55:@7581.4]
  wire [2:0] _T_7539; // @[Bitwise.scala 48:55:@7581.4]
  wire [3:0] _T_7540; // @[Bitwise.scala 48:55:@7582.4]
  wire [4:0] _T_7541; // @[Bitwise.scala 48:55:@7583.4]
  wire [5:0] _T_7542; // @[Bitwise.scala 48:55:@7584.4]
  wire [6:0] _T_7543; // @[Bitwise.scala 48:55:@7585.4]
  wire [48:0] _T_7607; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7650.4]
  wire  _T_7608; // @[Bitwise.scala 50:65:@7651.4]
  wire  _T_7609; // @[Bitwise.scala 50:65:@7652.4]
  wire  _T_7610; // @[Bitwise.scala 50:65:@7653.4]
  wire  _T_7611; // @[Bitwise.scala 50:65:@7654.4]
  wire  _T_7612; // @[Bitwise.scala 50:65:@7655.4]
  wire  _T_7613; // @[Bitwise.scala 50:65:@7656.4]
  wire  _T_7614; // @[Bitwise.scala 50:65:@7657.4]
  wire  _T_7615; // @[Bitwise.scala 50:65:@7658.4]
  wire  _T_7616; // @[Bitwise.scala 50:65:@7659.4]
  wire  _T_7617; // @[Bitwise.scala 50:65:@7660.4]
  wire  _T_7618; // @[Bitwise.scala 50:65:@7661.4]
  wire  _T_7619; // @[Bitwise.scala 50:65:@7662.4]
  wire  _T_7620; // @[Bitwise.scala 50:65:@7663.4]
  wire  _T_7621; // @[Bitwise.scala 50:65:@7664.4]
  wire  _T_7622; // @[Bitwise.scala 50:65:@7665.4]
  wire  _T_7623; // @[Bitwise.scala 50:65:@7666.4]
  wire  _T_7624; // @[Bitwise.scala 50:65:@7667.4]
  wire  _T_7625; // @[Bitwise.scala 50:65:@7668.4]
  wire  _T_7626; // @[Bitwise.scala 50:65:@7669.4]
  wire  _T_7627; // @[Bitwise.scala 50:65:@7670.4]
  wire  _T_7628; // @[Bitwise.scala 50:65:@7671.4]
  wire  _T_7629; // @[Bitwise.scala 50:65:@7672.4]
  wire  _T_7630; // @[Bitwise.scala 50:65:@7673.4]
  wire  _T_7631; // @[Bitwise.scala 50:65:@7674.4]
  wire  _T_7632; // @[Bitwise.scala 50:65:@7675.4]
  wire  _T_7633; // @[Bitwise.scala 50:65:@7676.4]
  wire  _T_7634; // @[Bitwise.scala 50:65:@7677.4]
  wire  _T_7635; // @[Bitwise.scala 50:65:@7678.4]
  wire  _T_7636; // @[Bitwise.scala 50:65:@7679.4]
  wire  _T_7637; // @[Bitwise.scala 50:65:@7680.4]
  wire  _T_7638; // @[Bitwise.scala 50:65:@7681.4]
  wire  _T_7639; // @[Bitwise.scala 50:65:@7682.4]
  wire  _T_7640; // @[Bitwise.scala 50:65:@7683.4]
  wire  _T_7641; // @[Bitwise.scala 50:65:@7684.4]
  wire  _T_7642; // @[Bitwise.scala 50:65:@7685.4]
  wire  _T_7643; // @[Bitwise.scala 50:65:@7686.4]
  wire  _T_7644; // @[Bitwise.scala 50:65:@7687.4]
  wire  _T_7645; // @[Bitwise.scala 50:65:@7688.4]
  wire  _T_7646; // @[Bitwise.scala 50:65:@7689.4]
  wire  _T_7647; // @[Bitwise.scala 50:65:@7690.4]
  wire  _T_7648; // @[Bitwise.scala 50:65:@7691.4]
  wire  _T_7649; // @[Bitwise.scala 50:65:@7692.4]
  wire  _T_7650; // @[Bitwise.scala 50:65:@7693.4]
  wire  _T_7651; // @[Bitwise.scala 50:65:@7694.4]
  wire  _T_7652; // @[Bitwise.scala 50:65:@7695.4]
  wire  _T_7653; // @[Bitwise.scala 50:65:@7696.4]
  wire  _T_7654; // @[Bitwise.scala 50:65:@7697.4]
  wire  _T_7655; // @[Bitwise.scala 50:65:@7698.4]
  wire  _T_7656; // @[Bitwise.scala 50:65:@7699.4]
  wire [1:0] _T_7657; // @[Bitwise.scala 48:55:@7700.4]
  wire [1:0] _GEN_877; // @[Bitwise.scala 48:55:@7701.4]
  wire [2:0] _T_7658; // @[Bitwise.scala 48:55:@7701.4]
  wire [1:0] _T_7659; // @[Bitwise.scala 48:55:@7702.4]
  wire [1:0] _GEN_878; // @[Bitwise.scala 48:55:@7703.4]
  wire [2:0] _T_7660; // @[Bitwise.scala 48:55:@7703.4]
  wire [3:0] _T_7661; // @[Bitwise.scala 48:55:@7704.4]
  wire [1:0] _T_7662; // @[Bitwise.scala 48:55:@7705.4]
  wire [1:0] _GEN_879; // @[Bitwise.scala 48:55:@7706.4]
  wire [2:0] _T_7663; // @[Bitwise.scala 48:55:@7706.4]
  wire [1:0] _T_7664; // @[Bitwise.scala 48:55:@7707.4]
  wire [1:0] _GEN_880; // @[Bitwise.scala 48:55:@7708.4]
  wire [2:0] _T_7665; // @[Bitwise.scala 48:55:@7708.4]
  wire [3:0] _T_7666; // @[Bitwise.scala 48:55:@7709.4]
  wire [4:0] _T_7667; // @[Bitwise.scala 48:55:@7710.4]
  wire [1:0] _T_7668; // @[Bitwise.scala 48:55:@7711.4]
  wire [1:0] _GEN_881; // @[Bitwise.scala 48:55:@7712.4]
  wire [2:0] _T_7669; // @[Bitwise.scala 48:55:@7712.4]
  wire [1:0] _T_7670; // @[Bitwise.scala 48:55:@7713.4]
  wire [1:0] _GEN_882; // @[Bitwise.scala 48:55:@7714.4]
  wire [2:0] _T_7671; // @[Bitwise.scala 48:55:@7714.4]
  wire [3:0] _T_7672; // @[Bitwise.scala 48:55:@7715.4]
  wire [1:0] _T_7673; // @[Bitwise.scala 48:55:@7716.4]
  wire [1:0] _GEN_883; // @[Bitwise.scala 48:55:@7717.4]
  wire [2:0] _T_7674; // @[Bitwise.scala 48:55:@7717.4]
  wire [1:0] _T_7675; // @[Bitwise.scala 48:55:@7718.4]
  wire [1:0] _GEN_884; // @[Bitwise.scala 48:55:@7719.4]
  wire [2:0] _T_7676; // @[Bitwise.scala 48:55:@7719.4]
  wire [3:0] _T_7677; // @[Bitwise.scala 48:55:@7720.4]
  wire [4:0] _T_7678; // @[Bitwise.scala 48:55:@7721.4]
  wire [5:0] _T_7679; // @[Bitwise.scala 48:55:@7722.4]
  wire [1:0] _T_7680; // @[Bitwise.scala 48:55:@7723.4]
  wire [1:0] _GEN_885; // @[Bitwise.scala 48:55:@7724.4]
  wire [2:0] _T_7681; // @[Bitwise.scala 48:55:@7724.4]
  wire [1:0] _T_7682; // @[Bitwise.scala 48:55:@7725.4]
  wire [1:0] _GEN_886; // @[Bitwise.scala 48:55:@7726.4]
  wire [2:0] _T_7683; // @[Bitwise.scala 48:55:@7726.4]
  wire [3:0] _T_7684; // @[Bitwise.scala 48:55:@7727.4]
  wire [1:0] _T_7685; // @[Bitwise.scala 48:55:@7728.4]
  wire [1:0] _GEN_887; // @[Bitwise.scala 48:55:@7729.4]
  wire [2:0] _T_7686; // @[Bitwise.scala 48:55:@7729.4]
  wire [1:0] _T_7687; // @[Bitwise.scala 48:55:@7730.4]
  wire [1:0] _GEN_888; // @[Bitwise.scala 48:55:@7731.4]
  wire [2:0] _T_7688; // @[Bitwise.scala 48:55:@7731.4]
  wire [3:0] _T_7689; // @[Bitwise.scala 48:55:@7732.4]
  wire [4:0] _T_7690; // @[Bitwise.scala 48:55:@7733.4]
  wire [1:0] _T_7691; // @[Bitwise.scala 48:55:@7734.4]
  wire [1:0] _GEN_889; // @[Bitwise.scala 48:55:@7735.4]
  wire [2:0] _T_7692; // @[Bitwise.scala 48:55:@7735.4]
  wire [1:0] _T_7693; // @[Bitwise.scala 48:55:@7736.4]
  wire [1:0] _GEN_890; // @[Bitwise.scala 48:55:@7737.4]
  wire [2:0] _T_7694; // @[Bitwise.scala 48:55:@7737.4]
  wire [3:0] _T_7695; // @[Bitwise.scala 48:55:@7738.4]
  wire [1:0] _T_7696; // @[Bitwise.scala 48:55:@7739.4]
  wire [1:0] _GEN_891; // @[Bitwise.scala 48:55:@7740.4]
  wire [2:0] _T_7697; // @[Bitwise.scala 48:55:@7740.4]
  wire [1:0] _T_7698; // @[Bitwise.scala 48:55:@7741.4]
  wire [1:0] _T_7699; // @[Bitwise.scala 48:55:@7742.4]
  wire [2:0] _T_7700; // @[Bitwise.scala 48:55:@7743.4]
  wire [3:0] _T_7701; // @[Bitwise.scala 48:55:@7744.4]
  wire [4:0] _T_7702; // @[Bitwise.scala 48:55:@7745.4]
  wire [5:0] _T_7703; // @[Bitwise.scala 48:55:@7746.4]
  wire [6:0] _T_7704; // @[Bitwise.scala 48:55:@7747.4]
  wire [49:0] _T_7768; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7812.4]
  wire  _T_7769; // @[Bitwise.scala 50:65:@7813.4]
  wire  _T_7770; // @[Bitwise.scala 50:65:@7814.4]
  wire  _T_7771; // @[Bitwise.scala 50:65:@7815.4]
  wire  _T_7772; // @[Bitwise.scala 50:65:@7816.4]
  wire  _T_7773; // @[Bitwise.scala 50:65:@7817.4]
  wire  _T_7774; // @[Bitwise.scala 50:65:@7818.4]
  wire  _T_7775; // @[Bitwise.scala 50:65:@7819.4]
  wire  _T_7776; // @[Bitwise.scala 50:65:@7820.4]
  wire  _T_7777; // @[Bitwise.scala 50:65:@7821.4]
  wire  _T_7778; // @[Bitwise.scala 50:65:@7822.4]
  wire  _T_7779; // @[Bitwise.scala 50:65:@7823.4]
  wire  _T_7780; // @[Bitwise.scala 50:65:@7824.4]
  wire  _T_7781; // @[Bitwise.scala 50:65:@7825.4]
  wire  _T_7782; // @[Bitwise.scala 50:65:@7826.4]
  wire  _T_7783; // @[Bitwise.scala 50:65:@7827.4]
  wire  _T_7784; // @[Bitwise.scala 50:65:@7828.4]
  wire  _T_7785; // @[Bitwise.scala 50:65:@7829.4]
  wire  _T_7786; // @[Bitwise.scala 50:65:@7830.4]
  wire  _T_7787; // @[Bitwise.scala 50:65:@7831.4]
  wire  _T_7788; // @[Bitwise.scala 50:65:@7832.4]
  wire  _T_7789; // @[Bitwise.scala 50:65:@7833.4]
  wire  _T_7790; // @[Bitwise.scala 50:65:@7834.4]
  wire  _T_7791; // @[Bitwise.scala 50:65:@7835.4]
  wire  _T_7792; // @[Bitwise.scala 50:65:@7836.4]
  wire  _T_7793; // @[Bitwise.scala 50:65:@7837.4]
  wire  _T_7794; // @[Bitwise.scala 50:65:@7838.4]
  wire  _T_7795; // @[Bitwise.scala 50:65:@7839.4]
  wire  _T_7796; // @[Bitwise.scala 50:65:@7840.4]
  wire  _T_7797; // @[Bitwise.scala 50:65:@7841.4]
  wire  _T_7798; // @[Bitwise.scala 50:65:@7842.4]
  wire  _T_7799; // @[Bitwise.scala 50:65:@7843.4]
  wire  _T_7800; // @[Bitwise.scala 50:65:@7844.4]
  wire  _T_7801; // @[Bitwise.scala 50:65:@7845.4]
  wire  _T_7802; // @[Bitwise.scala 50:65:@7846.4]
  wire  _T_7803; // @[Bitwise.scala 50:65:@7847.4]
  wire  _T_7804; // @[Bitwise.scala 50:65:@7848.4]
  wire  _T_7805; // @[Bitwise.scala 50:65:@7849.4]
  wire  _T_7806; // @[Bitwise.scala 50:65:@7850.4]
  wire  _T_7807; // @[Bitwise.scala 50:65:@7851.4]
  wire  _T_7808; // @[Bitwise.scala 50:65:@7852.4]
  wire  _T_7809; // @[Bitwise.scala 50:65:@7853.4]
  wire  _T_7810; // @[Bitwise.scala 50:65:@7854.4]
  wire  _T_7811; // @[Bitwise.scala 50:65:@7855.4]
  wire  _T_7812; // @[Bitwise.scala 50:65:@7856.4]
  wire  _T_7813; // @[Bitwise.scala 50:65:@7857.4]
  wire  _T_7814; // @[Bitwise.scala 50:65:@7858.4]
  wire  _T_7815; // @[Bitwise.scala 50:65:@7859.4]
  wire  _T_7816; // @[Bitwise.scala 50:65:@7860.4]
  wire  _T_7817; // @[Bitwise.scala 50:65:@7861.4]
  wire  _T_7818; // @[Bitwise.scala 50:65:@7862.4]
  wire [1:0] _T_7819; // @[Bitwise.scala 48:55:@7863.4]
  wire [1:0] _GEN_892; // @[Bitwise.scala 48:55:@7864.4]
  wire [2:0] _T_7820; // @[Bitwise.scala 48:55:@7864.4]
  wire [1:0] _T_7821; // @[Bitwise.scala 48:55:@7865.4]
  wire [1:0] _GEN_893; // @[Bitwise.scala 48:55:@7866.4]
  wire [2:0] _T_7822; // @[Bitwise.scala 48:55:@7866.4]
  wire [3:0] _T_7823; // @[Bitwise.scala 48:55:@7867.4]
  wire [1:0] _T_7824; // @[Bitwise.scala 48:55:@7868.4]
  wire [1:0] _GEN_894; // @[Bitwise.scala 48:55:@7869.4]
  wire [2:0] _T_7825; // @[Bitwise.scala 48:55:@7869.4]
  wire [1:0] _T_7826; // @[Bitwise.scala 48:55:@7870.4]
  wire [1:0] _GEN_895; // @[Bitwise.scala 48:55:@7871.4]
  wire [2:0] _T_7827; // @[Bitwise.scala 48:55:@7871.4]
  wire [3:0] _T_7828; // @[Bitwise.scala 48:55:@7872.4]
  wire [4:0] _T_7829; // @[Bitwise.scala 48:55:@7873.4]
  wire [1:0] _T_7830; // @[Bitwise.scala 48:55:@7874.4]
  wire [1:0] _GEN_896; // @[Bitwise.scala 48:55:@7875.4]
  wire [2:0] _T_7831; // @[Bitwise.scala 48:55:@7875.4]
  wire [1:0] _T_7832; // @[Bitwise.scala 48:55:@7876.4]
  wire [1:0] _GEN_897; // @[Bitwise.scala 48:55:@7877.4]
  wire [2:0] _T_7833; // @[Bitwise.scala 48:55:@7877.4]
  wire [3:0] _T_7834; // @[Bitwise.scala 48:55:@7878.4]
  wire [1:0] _T_7835; // @[Bitwise.scala 48:55:@7879.4]
  wire [1:0] _GEN_898; // @[Bitwise.scala 48:55:@7880.4]
  wire [2:0] _T_7836; // @[Bitwise.scala 48:55:@7880.4]
  wire [1:0] _T_7837; // @[Bitwise.scala 48:55:@7881.4]
  wire [1:0] _T_7838; // @[Bitwise.scala 48:55:@7882.4]
  wire [2:0] _T_7839; // @[Bitwise.scala 48:55:@7883.4]
  wire [3:0] _T_7840; // @[Bitwise.scala 48:55:@7884.4]
  wire [4:0] _T_7841; // @[Bitwise.scala 48:55:@7885.4]
  wire [5:0] _T_7842; // @[Bitwise.scala 48:55:@7886.4]
  wire [1:0] _T_7843; // @[Bitwise.scala 48:55:@7887.4]
  wire [1:0] _GEN_899; // @[Bitwise.scala 48:55:@7888.4]
  wire [2:0] _T_7844; // @[Bitwise.scala 48:55:@7888.4]
  wire [1:0] _T_7845; // @[Bitwise.scala 48:55:@7889.4]
  wire [1:0] _GEN_900; // @[Bitwise.scala 48:55:@7890.4]
  wire [2:0] _T_7846; // @[Bitwise.scala 48:55:@7890.4]
  wire [3:0] _T_7847; // @[Bitwise.scala 48:55:@7891.4]
  wire [1:0] _T_7848; // @[Bitwise.scala 48:55:@7892.4]
  wire [1:0] _GEN_901; // @[Bitwise.scala 48:55:@7893.4]
  wire [2:0] _T_7849; // @[Bitwise.scala 48:55:@7893.4]
  wire [1:0] _T_7850; // @[Bitwise.scala 48:55:@7894.4]
  wire [1:0] _GEN_902; // @[Bitwise.scala 48:55:@7895.4]
  wire [2:0] _T_7851; // @[Bitwise.scala 48:55:@7895.4]
  wire [3:0] _T_7852; // @[Bitwise.scala 48:55:@7896.4]
  wire [4:0] _T_7853; // @[Bitwise.scala 48:55:@7897.4]
  wire [1:0] _T_7854; // @[Bitwise.scala 48:55:@7898.4]
  wire [1:0] _GEN_903; // @[Bitwise.scala 48:55:@7899.4]
  wire [2:0] _T_7855; // @[Bitwise.scala 48:55:@7899.4]
  wire [1:0] _T_7856; // @[Bitwise.scala 48:55:@7900.4]
  wire [1:0] _GEN_904; // @[Bitwise.scala 48:55:@7901.4]
  wire [2:0] _T_7857; // @[Bitwise.scala 48:55:@7901.4]
  wire [3:0] _T_7858; // @[Bitwise.scala 48:55:@7902.4]
  wire [1:0] _T_7859; // @[Bitwise.scala 48:55:@7903.4]
  wire [1:0] _GEN_905; // @[Bitwise.scala 48:55:@7904.4]
  wire [2:0] _T_7860; // @[Bitwise.scala 48:55:@7904.4]
  wire [1:0] _T_7861; // @[Bitwise.scala 48:55:@7905.4]
  wire [1:0] _T_7862; // @[Bitwise.scala 48:55:@7906.4]
  wire [2:0] _T_7863; // @[Bitwise.scala 48:55:@7907.4]
  wire [3:0] _T_7864; // @[Bitwise.scala 48:55:@7908.4]
  wire [4:0] _T_7865; // @[Bitwise.scala 48:55:@7909.4]
  wire [5:0] _T_7866; // @[Bitwise.scala 48:55:@7910.4]
  wire [6:0] _T_7867; // @[Bitwise.scala 48:55:@7911.4]
  wire [50:0] _T_7931; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7976.4]
  wire  _T_7932; // @[Bitwise.scala 50:65:@7977.4]
  wire  _T_7933; // @[Bitwise.scala 50:65:@7978.4]
  wire  _T_7934; // @[Bitwise.scala 50:65:@7979.4]
  wire  _T_7935; // @[Bitwise.scala 50:65:@7980.4]
  wire  _T_7936; // @[Bitwise.scala 50:65:@7981.4]
  wire  _T_7937; // @[Bitwise.scala 50:65:@7982.4]
  wire  _T_7938; // @[Bitwise.scala 50:65:@7983.4]
  wire  _T_7939; // @[Bitwise.scala 50:65:@7984.4]
  wire  _T_7940; // @[Bitwise.scala 50:65:@7985.4]
  wire  _T_7941; // @[Bitwise.scala 50:65:@7986.4]
  wire  _T_7942; // @[Bitwise.scala 50:65:@7987.4]
  wire  _T_7943; // @[Bitwise.scala 50:65:@7988.4]
  wire  _T_7944; // @[Bitwise.scala 50:65:@7989.4]
  wire  _T_7945; // @[Bitwise.scala 50:65:@7990.4]
  wire  _T_7946; // @[Bitwise.scala 50:65:@7991.4]
  wire  _T_7947; // @[Bitwise.scala 50:65:@7992.4]
  wire  _T_7948; // @[Bitwise.scala 50:65:@7993.4]
  wire  _T_7949; // @[Bitwise.scala 50:65:@7994.4]
  wire  _T_7950; // @[Bitwise.scala 50:65:@7995.4]
  wire  _T_7951; // @[Bitwise.scala 50:65:@7996.4]
  wire  _T_7952; // @[Bitwise.scala 50:65:@7997.4]
  wire  _T_7953; // @[Bitwise.scala 50:65:@7998.4]
  wire  _T_7954; // @[Bitwise.scala 50:65:@7999.4]
  wire  _T_7955; // @[Bitwise.scala 50:65:@8000.4]
  wire  _T_7956; // @[Bitwise.scala 50:65:@8001.4]
  wire  _T_7957; // @[Bitwise.scala 50:65:@8002.4]
  wire  _T_7958; // @[Bitwise.scala 50:65:@8003.4]
  wire  _T_7959; // @[Bitwise.scala 50:65:@8004.4]
  wire  _T_7960; // @[Bitwise.scala 50:65:@8005.4]
  wire  _T_7961; // @[Bitwise.scala 50:65:@8006.4]
  wire  _T_7962; // @[Bitwise.scala 50:65:@8007.4]
  wire  _T_7963; // @[Bitwise.scala 50:65:@8008.4]
  wire  _T_7964; // @[Bitwise.scala 50:65:@8009.4]
  wire  _T_7965; // @[Bitwise.scala 50:65:@8010.4]
  wire  _T_7966; // @[Bitwise.scala 50:65:@8011.4]
  wire  _T_7967; // @[Bitwise.scala 50:65:@8012.4]
  wire  _T_7968; // @[Bitwise.scala 50:65:@8013.4]
  wire  _T_7969; // @[Bitwise.scala 50:65:@8014.4]
  wire  _T_7970; // @[Bitwise.scala 50:65:@8015.4]
  wire  _T_7971; // @[Bitwise.scala 50:65:@8016.4]
  wire  _T_7972; // @[Bitwise.scala 50:65:@8017.4]
  wire  _T_7973; // @[Bitwise.scala 50:65:@8018.4]
  wire  _T_7974; // @[Bitwise.scala 50:65:@8019.4]
  wire  _T_7975; // @[Bitwise.scala 50:65:@8020.4]
  wire  _T_7976; // @[Bitwise.scala 50:65:@8021.4]
  wire  _T_7977; // @[Bitwise.scala 50:65:@8022.4]
  wire  _T_7978; // @[Bitwise.scala 50:65:@8023.4]
  wire  _T_7979; // @[Bitwise.scala 50:65:@8024.4]
  wire  _T_7980; // @[Bitwise.scala 50:65:@8025.4]
  wire  _T_7981; // @[Bitwise.scala 50:65:@8026.4]
  wire  _T_7982; // @[Bitwise.scala 50:65:@8027.4]
  wire [1:0] _T_7983; // @[Bitwise.scala 48:55:@8028.4]
  wire [1:0] _GEN_906; // @[Bitwise.scala 48:55:@8029.4]
  wire [2:0] _T_7984; // @[Bitwise.scala 48:55:@8029.4]
  wire [1:0] _T_7985; // @[Bitwise.scala 48:55:@8030.4]
  wire [1:0] _GEN_907; // @[Bitwise.scala 48:55:@8031.4]
  wire [2:0] _T_7986; // @[Bitwise.scala 48:55:@8031.4]
  wire [3:0] _T_7987; // @[Bitwise.scala 48:55:@8032.4]
  wire [1:0] _T_7988; // @[Bitwise.scala 48:55:@8033.4]
  wire [1:0] _GEN_908; // @[Bitwise.scala 48:55:@8034.4]
  wire [2:0] _T_7989; // @[Bitwise.scala 48:55:@8034.4]
  wire [1:0] _T_7990; // @[Bitwise.scala 48:55:@8035.4]
  wire [1:0] _GEN_909; // @[Bitwise.scala 48:55:@8036.4]
  wire [2:0] _T_7991; // @[Bitwise.scala 48:55:@8036.4]
  wire [3:0] _T_7992; // @[Bitwise.scala 48:55:@8037.4]
  wire [4:0] _T_7993; // @[Bitwise.scala 48:55:@8038.4]
  wire [1:0] _T_7994; // @[Bitwise.scala 48:55:@8039.4]
  wire [1:0] _GEN_910; // @[Bitwise.scala 48:55:@8040.4]
  wire [2:0] _T_7995; // @[Bitwise.scala 48:55:@8040.4]
  wire [1:0] _T_7996; // @[Bitwise.scala 48:55:@8041.4]
  wire [1:0] _GEN_911; // @[Bitwise.scala 48:55:@8042.4]
  wire [2:0] _T_7997; // @[Bitwise.scala 48:55:@8042.4]
  wire [3:0] _T_7998; // @[Bitwise.scala 48:55:@8043.4]
  wire [1:0] _T_7999; // @[Bitwise.scala 48:55:@8044.4]
  wire [1:0] _GEN_912; // @[Bitwise.scala 48:55:@8045.4]
  wire [2:0] _T_8000; // @[Bitwise.scala 48:55:@8045.4]
  wire [1:0] _T_8001; // @[Bitwise.scala 48:55:@8046.4]
  wire [1:0] _T_8002; // @[Bitwise.scala 48:55:@8047.4]
  wire [2:0] _T_8003; // @[Bitwise.scala 48:55:@8048.4]
  wire [3:0] _T_8004; // @[Bitwise.scala 48:55:@8049.4]
  wire [4:0] _T_8005; // @[Bitwise.scala 48:55:@8050.4]
  wire [5:0] _T_8006; // @[Bitwise.scala 48:55:@8051.4]
  wire [1:0] _T_8007; // @[Bitwise.scala 48:55:@8052.4]
  wire [1:0] _GEN_913; // @[Bitwise.scala 48:55:@8053.4]
  wire [2:0] _T_8008; // @[Bitwise.scala 48:55:@8053.4]
  wire [1:0] _T_8009; // @[Bitwise.scala 48:55:@8054.4]
  wire [1:0] _GEN_914; // @[Bitwise.scala 48:55:@8055.4]
  wire [2:0] _T_8010; // @[Bitwise.scala 48:55:@8055.4]
  wire [3:0] _T_8011; // @[Bitwise.scala 48:55:@8056.4]
  wire [1:0] _T_8012; // @[Bitwise.scala 48:55:@8057.4]
  wire [1:0] _GEN_915; // @[Bitwise.scala 48:55:@8058.4]
  wire [2:0] _T_8013; // @[Bitwise.scala 48:55:@8058.4]
  wire [1:0] _T_8014; // @[Bitwise.scala 48:55:@8059.4]
  wire [1:0] _T_8015; // @[Bitwise.scala 48:55:@8060.4]
  wire [2:0] _T_8016; // @[Bitwise.scala 48:55:@8061.4]
  wire [3:0] _T_8017; // @[Bitwise.scala 48:55:@8062.4]
  wire [4:0] _T_8018; // @[Bitwise.scala 48:55:@8063.4]
  wire [1:0] _T_8019; // @[Bitwise.scala 48:55:@8064.4]
  wire [1:0] _GEN_916; // @[Bitwise.scala 48:55:@8065.4]
  wire [2:0] _T_8020; // @[Bitwise.scala 48:55:@8065.4]
  wire [1:0] _T_8021; // @[Bitwise.scala 48:55:@8066.4]
  wire [1:0] _GEN_917; // @[Bitwise.scala 48:55:@8067.4]
  wire [2:0] _T_8022; // @[Bitwise.scala 48:55:@8067.4]
  wire [3:0] _T_8023; // @[Bitwise.scala 48:55:@8068.4]
  wire [1:0] _T_8024; // @[Bitwise.scala 48:55:@8069.4]
  wire [1:0] _GEN_918; // @[Bitwise.scala 48:55:@8070.4]
  wire [2:0] _T_8025; // @[Bitwise.scala 48:55:@8070.4]
  wire [1:0] _T_8026; // @[Bitwise.scala 48:55:@8071.4]
  wire [1:0] _T_8027; // @[Bitwise.scala 48:55:@8072.4]
  wire [2:0] _T_8028; // @[Bitwise.scala 48:55:@8073.4]
  wire [3:0] _T_8029; // @[Bitwise.scala 48:55:@8074.4]
  wire [4:0] _T_8030; // @[Bitwise.scala 48:55:@8075.4]
  wire [5:0] _T_8031; // @[Bitwise.scala 48:55:@8076.4]
  wire [6:0] _T_8032; // @[Bitwise.scala 48:55:@8077.4]
  wire [51:0] _T_8096; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@8142.4]
  wire  _T_8097; // @[Bitwise.scala 50:65:@8143.4]
  wire  _T_8098; // @[Bitwise.scala 50:65:@8144.4]
  wire  _T_8099; // @[Bitwise.scala 50:65:@8145.4]
  wire  _T_8100; // @[Bitwise.scala 50:65:@8146.4]
  wire  _T_8101; // @[Bitwise.scala 50:65:@8147.4]
  wire  _T_8102; // @[Bitwise.scala 50:65:@8148.4]
  wire  _T_8103; // @[Bitwise.scala 50:65:@8149.4]
  wire  _T_8104; // @[Bitwise.scala 50:65:@8150.4]
  wire  _T_8105; // @[Bitwise.scala 50:65:@8151.4]
  wire  _T_8106; // @[Bitwise.scala 50:65:@8152.4]
  wire  _T_8107; // @[Bitwise.scala 50:65:@8153.4]
  wire  _T_8108; // @[Bitwise.scala 50:65:@8154.4]
  wire  _T_8109; // @[Bitwise.scala 50:65:@8155.4]
  wire  _T_8110; // @[Bitwise.scala 50:65:@8156.4]
  wire  _T_8111; // @[Bitwise.scala 50:65:@8157.4]
  wire  _T_8112; // @[Bitwise.scala 50:65:@8158.4]
  wire  _T_8113; // @[Bitwise.scala 50:65:@8159.4]
  wire  _T_8114; // @[Bitwise.scala 50:65:@8160.4]
  wire  _T_8115; // @[Bitwise.scala 50:65:@8161.4]
  wire  _T_8116; // @[Bitwise.scala 50:65:@8162.4]
  wire  _T_8117; // @[Bitwise.scala 50:65:@8163.4]
  wire  _T_8118; // @[Bitwise.scala 50:65:@8164.4]
  wire  _T_8119; // @[Bitwise.scala 50:65:@8165.4]
  wire  _T_8120; // @[Bitwise.scala 50:65:@8166.4]
  wire  _T_8121; // @[Bitwise.scala 50:65:@8167.4]
  wire  _T_8122; // @[Bitwise.scala 50:65:@8168.4]
  wire  _T_8123; // @[Bitwise.scala 50:65:@8169.4]
  wire  _T_8124; // @[Bitwise.scala 50:65:@8170.4]
  wire  _T_8125; // @[Bitwise.scala 50:65:@8171.4]
  wire  _T_8126; // @[Bitwise.scala 50:65:@8172.4]
  wire  _T_8127; // @[Bitwise.scala 50:65:@8173.4]
  wire  _T_8128; // @[Bitwise.scala 50:65:@8174.4]
  wire  _T_8129; // @[Bitwise.scala 50:65:@8175.4]
  wire  _T_8130; // @[Bitwise.scala 50:65:@8176.4]
  wire  _T_8131; // @[Bitwise.scala 50:65:@8177.4]
  wire  _T_8132; // @[Bitwise.scala 50:65:@8178.4]
  wire  _T_8133; // @[Bitwise.scala 50:65:@8179.4]
  wire  _T_8134; // @[Bitwise.scala 50:65:@8180.4]
  wire  _T_8135; // @[Bitwise.scala 50:65:@8181.4]
  wire  _T_8136; // @[Bitwise.scala 50:65:@8182.4]
  wire  _T_8137; // @[Bitwise.scala 50:65:@8183.4]
  wire  _T_8138; // @[Bitwise.scala 50:65:@8184.4]
  wire  _T_8139; // @[Bitwise.scala 50:65:@8185.4]
  wire  _T_8140; // @[Bitwise.scala 50:65:@8186.4]
  wire  _T_8141; // @[Bitwise.scala 50:65:@8187.4]
  wire  _T_8142; // @[Bitwise.scala 50:65:@8188.4]
  wire  _T_8143; // @[Bitwise.scala 50:65:@8189.4]
  wire  _T_8144; // @[Bitwise.scala 50:65:@8190.4]
  wire  _T_8145; // @[Bitwise.scala 50:65:@8191.4]
  wire  _T_8146; // @[Bitwise.scala 50:65:@8192.4]
  wire  _T_8147; // @[Bitwise.scala 50:65:@8193.4]
  wire  _T_8148; // @[Bitwise.scala 50:65:@8194.4]
  wire [1:0] _T_8149; // @[Bitwise.scala 48:55:@8195.4]
  wire [1:0] _GEN_919; // @[Bitwise.scala 48:55:@8196.4]
  wire [2:0] _T_8150; // @[Bitwise.scala 48:55:@8196.4]
  wire [1:0] _T_8151; // @[Bitwise.scala 48:55:@8197.4]
  wire [1:0] _GEN_920; // @[Bitwise.scala 48:55:@8198.4]
  wire [2:0] _T_8152; // @[Bitwise.scala 48:55:@8198.4]
  wire [3:0] _T_8153; // @[Bitwise.scala 48:55:@8199.4]
  wire [1:0] _T_8154; // @[Bitwise.scala 48:55:@8200.4]
  wire [1:0] _GEN_921; // @[Bitwise.scala 48:55:@8201.4]
  wire [2:0] _T_8155; // @[Bitwise.scala 48:55:@8201.4]
  wire [1:0] _T_8156; // @[Bitwise.scala 48:55:@8202.4]
  wire [1:0] _T_8157; // @[Bitwise.scala 48:55:@8203.4]
  wire [2:0] _T_8158; // @[Bitwise.scala 48:55:@8204.4]
  wire [3:0] _T_8159; // @[Bitwise.scala 48:55:@8205.4]
  wire [4:0] _T_8160; // @[Bitwise.scala 48:55:@8206.4]
  wire [1:0] _T_8161; // @[Bitwise.scala 48:55:@8207.4]
  wire [1:0] _GEN_922; // @[Bitwise.scala 48:55:@8208.4]
  wire [2:0] _T_8162; // @[Bitwise.scala 48:55:@8208.4]
  wire [1:0] _T_8163; // @[Bitwise.scala 48:55:@8209.4]
  wire [1:0] _GEN_923; // @[Bitwise.scala 48:55:@8210.4]
  wire [2:0] _T_8164; // @[Bitwise.scala 48:55:@8210.4]
  wire [3:0] _T_8165; // @[Bitwise.scala 48:55:@8211.4]
  wire [1:0] _T_8166; // @[Bitwise.scala 48:55:@8212.4]
  wire [1:0] _GEN_924; // @[Bitwise.scala 48:55:@8213.4]
  wire [2:0] _T_8167; // @[Bitwise.scala 48:55:@8213.4]
  wire [1:0] _T_8168; // @[Bitwise.scala 48:55:@8214.4]
  wire [1:0] _T_8169; // @[Bitwise.scala 48:55:@8215.4]
  wire [2:0] _T_8170; // @[Bitwise.scala 48:55:@8216.4]
  wire [3:0] _T_8171; // @[Bitwise.scala 48:55:@8217.4]
  wire [4:0] _T_8172; // @[Bitwise.scala 48:55:@8218.4]
  wire [5:0] _T_8173; // @[Bitwise.scala 48:55:@8219.4]
  wire [1:0] _T_8174; // @[Bitwise.scala 48:55:@8220.4]
  wire [1:0] _GEN_925; // @[Bitwise.scala 48:55:@8221.4]
  wire [2:0] _T_8175; // @[Bitwise.scala 48:55:@8221.4]
  wire [1:0] _T_8176; // @[Bitwise.scala 48:55:@8222.4]
  wire [1:0] _GEN_926; // @[Bitwise.scala 48:55:@8223.4]
  wire [2:0] _T_8177; // @[Bitwise.scala 48:55:@8223.4]
  wire [3:0] _T_8178; // @[Bitwise.scala 48:55:@8224.4]
  wire [1:0] _T_8179; // @[Bitwise.scala 48:55:@8225.4]
  wire [1:0] _GEN_927; // @[Bitwise.scala 48:55:@8226.4]
  wire [2:0] _T_8180; // @[Bitwise.scala 48:55:@8226.4]
  wire [1:0] _T_8181; // @[Bitwise.scala 48:55:@8227.4]
  wire [1:0] _T_8182; // @[Bitwise.scala 48:55:@8228.4]
  wire [2:0] _T_8183; // @[Bitwise.scala 48:55:@8229.4]
  wire [3:0] _T_8184; // @[Bitwise.scala 48:55:@8230.4]
  wire [4:0] _T_8185; // @[Bitwise.scala 48:55:@8231.4]
  wire [1:0] _T_8186; // @[Bitwise.scala 48:55:@8232.4]
  wire [1:0] _GEN_928; // @[Bitwise.scala 48:55:@8233.4]
  wire [2:0] _T_8187; // @[Bitwise.scala 48:55:@8233.4]
  wire [1:0] _T_8188; // @[Bitwise.scala 48:55:@8234.4]
  wire [1:0] _GEN_929; // @[Bitwise.scala 48:55:@8235.4]
  wire [2:0] _T_8189; // @[Bitwise.scala 48:55:@8235.4]
  wire [3:0] _T_8190; // @[Bitwise.scala 48:55:@8236.4]
  wire [1:0] _T_8191; // @[Bitwise.scala 48:55:@8237.4]
  wire [1:0] _GEN_930; // @[Bitwise.scala 48:55:@8238.4]
  wire [2:0] _T_8192; // @[Bitwise.scala 48:55:@8238.4]
  wire [1:0] _T_8193; // @[Bitwise.scala 48:55:@8239.4]
  wire [1:0] _T_8194; // @[Bitwise.scala 48:55:@8240.4]
  wire [2:0] _T_8195; // @[Bitwise.scala 48:55:@8241.4]
  wire [3:0] _T_8196; // @[Bitwise.scala 48:55:@8242.4]
  wire [4:0] _T_8197; // @[Bitwise.scala 48:55:@8243.4]
  wire [5:0] _T_8198; // @[Bitwise.scala 48:55:@8244.4]
  wire [6:0] _T_8199; // @[Bitwise.scala 48:55:@8245.4]
  wire [52:0] _T_8263; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@8310.4]
  wire  _T_8264; // @[Bitwise.scala 50:65:@8311.4]
  wire  _T_8265; // @[Bitwise.scala 50:65:@8312.4]
  wire  _T_8266; // @[Bitwise.scala 50:65:@8313.4]
  wire  _T_8267; // @[Bitwise.scala 50:65:@8314.4]
  wire  _T_8268; // @[Bitwise.scala 50:65:@8315.4]
  wire  _T_8269; // @[Bitwise.scala 50:65:@8316.4]
  wire  _T_8270; // @[Bitwise.scala 50:65:@8317.4]
  wire  _T_8271; // @[Bitwise.scala 50:65:@8318.4]
  wire  _T_8272; // @[Bitwise.scala 50:65:@8319.4]
  wire  _T_8273; // @[Bitwise.scala 50:65:@8320.4]
  wire  _T_8274; // @[Bitwise.scala 50:65:@8321.4]
  wire  _T_8275; // @[Bitwise.scala 50:65:@8322.4]
  wire  _T_8276; // @[Bitwise.scala 50:65:@8323.4]
  wire  _T_8277; // @[Bitwise.scala 50:65:@8324.4]
  wire  _T_8278; // @[Bitwise.scala 50:65:@8325.4]
  wire  _T_8279; // @[Bitwise.scala 50:65:@8326.4]
  wire  _T_8280; // @[Bitwise.scala 50:65:@8327.4]
  wire  _T_8281; // @[Bitwise.scala 50:65:@8328.4]
  wire  _T_8282; // @[Bitwise.scala 50:65:@8329.4]
  wire  _T_8283; // @[Bitwise.scala 50:65:@8330.4]
  wire  _T_8284; // @[Bitwise.scala 50:65:@8331.4]
  wire  _T_8285; // @[Bitwise.scala 50:65:@8332.4]
  wire  _T_8286; // @[Bitwise.scala 50:65:@8333.4]
  wire  _T_8287; // @[Bitwise.scala 50:65:@8334.4]
  wire  _T_8288; // @[Bitwise.scala 50:65:@8335.4]
  wire  _T_8289; // @[Bitwise.scala 50:65:@8336.4]
  wire  _T_8290; // @[Bitwise.scala 50:65:@8337.4]
  wire  _T_8291; // @[Bitwise.scala 50:65:@8338.4]
  wire  _T_8292; // @[Bitwise.scala 50:65:@8339.4]
  wire  _T_8293; // @[Bitwise.scala 50:65:@8340.4]
  wire  _T_8294; // @[Bitwise.scala 50:65:@8341.4]
  wire  _T_8295; // @[Bitwise.scala 50:65:@8342.4]
  wire  _T_8296; // @[Bitwise.scala 50:65:@8343.4]
  wire  _T_8297; // @[Bitwise.scala 50:65:@8344.4]
  wire  _T_8298; // @[Bitwise.scala 50:65:@8345.4]
  wire  _T_8299; // @[Bitwise.scala 50:65:@8346.4]
  wire  _T_8300; // @[Bitwise.scala 50:65:@8347.4]
  wire  _T_8301; // @[Bitwise.scala 50:65:@8348.4]
  wire  _T_8302; // @[Bitwise.scala 50:65:@8349.4]
  wire  _T_8303; // @[Bitwise.scala 50:65:@8350.4]
  wire  _T_8304; // @[Bitwise.scala 50:65:@8351.4]
  wire  _T_8305; // @[Bitwise.scala 50:65:@8352.4]
  wire  _T_8306; // @[Bitwise.scala 50:65:@8353.4]
  wire  _T_8307; // @[Bitwise.scala 50:65:@8354.4]
  wire  _T_8308; // @[Bitwise.scala 50:65:@8355.4]
  wire  _T_8309; // @[Bitwise.scala 50:65:@8356.4]
  wire  _T_8310; // @[Bitwise.scala 50:65:@8357.4]
  wire  _T_8311; // @[Bitwise.scala 50:65:@8358.4]
  wire  _T_8312; // @[Bitwise.scala 50:65:@8359.4]
  wire  _T_8313; // @[Bitwise.scala 50:65:@8360.4]
  wire  _T_8314; // @[Bitwise.scala 50:65:@8361.4]
  wire  _T_8315; // @[Bitwise.scala 50:65:@8362.4]
  wire  _T_8316; // @[Bitwise.scala 50:65:@8363.4]
  wire [1:0] _T_8317; // @[Bitwise.scala 48:55:@8364.4]
  wire [1:0] _GEN_931; // @[Bitwise.scala 48:55:@8365.4]
  wire [2:0] _T_8318; // @[Bitwise.scala 48:55:@8365.4]
  wire [1:0] _T_8319; // @[Bitwise.scala 48:55:@8366.4]
  wire [1:0] _GEN_932; // @[Bitwise.scala 48:55:@8367.4]
  wire [2:0] _T_8320; // @[Bitwise.scala 48:55:@8367.4]
  wire [3:0] _T_8321; // @[Bitwise.scala 48:55:@8368.4]
  wire [1:0] _T_8322; // @[Bitwise.scala 48:55:@8369.4]
  wire [1:0] _GEN_933; // @[Bitwise.scala 48:55:@8370.4]
  wire [2:0] _T_8323; // @[Bitwise.scala 48:55:@8370.4]
  wire [1:0] _T_8324; // @[Bitwise.scala 48:55:@8371.4]
  wire [1:0] _T_8325; // @[Bitwise.scala 48:55:@8372.4]
  wire [2:0] _T_8326; // @[Bitwise.scala 48:55:@8373.4]
  wire [3:0] _T_8327; // @[Bitwise.scala 48:55:@8374.4]
  wire [4:0] _T_8328; // @[Bitwise.scala 48:55:@8375.4]
  wire [1:0] _T_8329; // @[Bitwise.scala 48:55:@8376.4]
  wire [1:0] _GEN_934; // @[Bitwise.scala 48:55:@8377.4]
  wire [2:0] _T_8330; // @[Bitwise.scala 48:55:@8377.4]
  wire [1:0] _T_8331; // @[Bitwise.scala 48:55:@8378.4]
  wire [1:0] _GEN_935; // @[Bitwise.scala 48:55:@8379.4]
  wire [2:0] _T_8332; // @[Bitwise.scala 48:55:@8379.4]
  wire [3:0] _T_8333; // @[Bitwise.scala 48:55:@8380.4]
  wire [1:0] _T_8334; // @[Bitwise.scala 48:55:@8381.4]
  wire [1:0] _GEN_936; // @[Bitwise.scala 48:55:@8382.4]
  wire [2:0] _T_8335; // @[Bitwise.scala 48:55:@8382.4]
  wire [1:0] _T_8336; // @[Bitwise.scala 48:55:@8383.4]
  wire [1:0] _T_8337; // @[Bitwise.scala 48:55:@8384.4]
  wire [2:0] _T_8338; // @[Bitwise.scala 48:55:@8385.4]
  wire [3:0] _T_8339; // @[Bitwise.scala 48:55:@8386.4]
  wire [4:0] _T_8340; // @[Bitwise.scala 48:55:@8387.4]
  wire [5:0] _T_8341; // @[Bitwise.scala 48:55:@8388.4]
  wire [1:0] _T_8342; // @[Bitwise.scala 48:55:@8389.4]
  wire [1:0] _GEN_937; // @[Bitwise.scala 48:55:@8390.4]
  wire [2:0] _T_8343; // @[Bitwise.scala 48:55:@8390.4]
  wire [1:0] _T_8344; // @[Bitwise.scala 48:55:@8391.4]
  wire [1:0] _GEN_938; // @[Bitwise.scala 48:55:@8392.4]
  wire [2:0] _T_8345; // @[Bitwise.scala 48:55:@8392.4]
  wire [3:0] _T_8346; // @[Bitwise.scala 48:55:@8393.4]
  wire [1:0] _T_8347; // @[Bitwise.scala 48:55:@8394.4]
  wire [1:0] _GEN_939; // @[Bitwise.scala 48:55:@8395.4]
  wire [2:0] _T_8348; // @[Bitwise.scala 48:55:@8395.4]
  wire [1:0] _T_8349; // @[Bitwise.scala 48:55:@8396.4]
  wire [1:0] _T_8350; // @[Bitwise.scala 48:55:@8397.4]
  wire [2:0] _T_8351; // @[Bitwise.scala 48:55:@8398.4]
  wire [3:0] _T_8352; // @[Bitwise.scala 48:55:@8399.4]
  wire [4:0] _T_8353; // @[Bitwise.scala 48:55:@8400.4]
  wire [1:0] _T_8354; // @[Bitwise.scala 48:55:@8401.4]
  wire [1:0] _GEN_940; // @[Bitwise.scala 48:55:@8402.4]
  wire [2:0] _T_8355; // @[Bitwise.scala 48:55:@8402.4]
  wire [1:0] _T_8356; // @[Bitwise.scala 48:55:@8403.4]
  wire [1:0] _T_8357; // @[Bitwise.scala 48:55:@8404.4]
  wire [2:0] _T_8358; // @[Bitwise.scala 48:55:@8405.4]
  wire [3:0] _T_8359; // @[Bitwise.scala 48:55:@8406.4]
  wire [1:0] _T_8360; // @[Bitwise.scala 48:55:@8407.4]
  wire [1:0] _GEN_941; // @[Bitwise.scala 48:55:@8408.4]
  wire [2:0] _T_8361; // @[Bitwise.scala 48:55:@8408.4]
  wire [1:0] _T_8362; // @[Bitwise.scala 48:55:@8409.4]
  wire [1:0] _T_8363; // @[Bitwise.scala 48:55:@8410.4]
  wire [2:0] _T_8364; // @[Bitwise.scala 48:55:@8411.4]
  wire [3:0] _T_8365; // @[Bitwise.scala 48:55:@8412.4]
  wire [4:0] _T_8366; // @[Bitwise.scala 48:55:@8413.4]
  wire [5:0] _T_8367; // @[Bitwise.scala 48:55:@8414.4]
  wire [6:0] _T_8368; // @[Bitwise.scala 48:55:@8415.4]
  wire [53:0] _T_8432; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@8480.4]
  wire  _T_8433; // @[Bitwise.scala 50:65:@8481.4]
  wire  _T_8434; // @[Bitwise.scala 50:65:@8482.4]
  wire  _T_8435; // @[Bitwise.scala 50:65:@8483.4]
  wire  _T_8436; // @[Bitwise.scala 50:65:@8484.4]
  wire  _T_8437; // @[Bitwise.scala 50:65:@8485.4]
  wire  _T_8438; // @[Bitwise.scala 50:65:@8486.4]
  wire  _T_8439; // @[Bitwise.scala 50:65:@8487.4]
  wire  _T_8440; // @[Bitwise.scala 50:65:@8488.4]
  wire  _T_8441; // @[Bitwise.scala 50:65:@8489.4]
  wire  _T_8442; // @[Bitwise.scala 50:65:@8490.4]
  wire  _T_8443; // @[Bitwise.scala 50:65:@8491.4]
  wire  _T_8444; // @[Bitwise.scala 50:65:@8492.4]
  wire  _T_8445; // @[Bitwise.scala 50:65:@8493.4]
  wire  _T_8446; // @[Bitwise.scala 50:65:@8494.4]
  wire  _T_8447; // @[Bitwise.scala 50:65:@8495.4]
  wire  _T_8448; // @[Bitwise.scala 50:65:@8496.4]
  wire  _T_8449; // @[Bitwise.scala 50:65:@8497.4]
  wire  _T_8450; // @[Bitwise.scala 50:65:@8498.4]
  wire  _T_8451; // @[Bitwise.scala 50:65:@8499.4]
  wire  _T_8452; // @[Bitwise.scala 50:65:@8500.4]
  wire  _T_8453; // @[Bitwise.scala 50:65:@8501.4]
  wire  _T_8454; // @[Bitwise.scala 50:65:@8502.4]
  wire  _T_8455; // @[Bitwise.scala 50:65:@8503.4]
  wire  _T_8456; // @[Bitwise.scala 50:65:@8504.4]
  wire  _T_8457; // @[Bitwise.scala 50:65:@8505.4]
  wire  _T_8458; // @[Bitwise.scala 50:65:@8506.4]
  wire  _T_8459; // @[Bitwise.scala 50:65:@8507.4]
  wire  _T_8460; // @[Bitwise.scala 50:65:@8508.4]
  wire  _T_8461; // @[Bitwise.scala 50:65:@8509.4]
  wire  _T_8462; // @[Bitwise.scala 50:65:@8510.4]
  wire  _T_8463; // @[Bitwise.scala 50:65:@8511.4]
  wire  _T_8464; // @[Bitwise.scala 50:65:@8512.4]
  wire  _T_8465; // @[Bitwise.scala 50:65:@8513.4]
  wire  _T_8466; // @[Bitwise.scala 50:65:@8514.4]
  wire  _T_8467; // @[Bitwise.scala 50:65:@8515.4]
  wire  _T_8468; // @[Bitwise.scala 50:65:@8516.4]
  wire  _T_8469; // @[Bitwise.scala 50:65:@8517.4]
  wire  _T_8470; // @[Bitwise.scala 50:65:@8518.4]
  wire  _T_8471; // @[Bitwise.scala 50:65:@8519.4]
  wire  _T_8472; // @[Bitwise.scala 50:65:@8520.4]
  wire  _T_8473; // @[Bitwise.scala 50:65:@8521.4]
  wire  _T_8474; // @[Bitwise.scala 50:65:@8522.4]
  wire  _T_8475; // @[Bitwise.scala 50:65:@8523.4]
  wire  _T_8476; // @[Bitwise.scala 50:65:@8524.4]
  wire  _T_8477; // @[Bitwise.scala 50:65:@8525.4]
  wire  _T_8478; // @[Bitwise.scala 50:65:@8526.4]
  wire  _T_8479; // @[Bitwise.scala 50:65:@8527.4]
  wire  _T_8480; // @[Bitwise.scala 50:65:@8528.4]
  wire  _T_8481; // @[Bitwise.scala 50:65:@8529.4]
  wire  _T_8482; // @[Bitwise.scala 50:65:@8530.4]
  wire  _T_8483; // @[Bitwise.scala 50:65:@8531.4]
  wire  _T_8484; // @[Bitwise.scala 50:65:@8532.4]
  wire  _T_8485; // @[Bitwise.scala 50:65:@8533.4]
  wire  _T_8486; // @[Bitwise.scala 50:65:@8534.4]
  wire [1:0] _T_8487; // @[Bitwise.scala 48:55:@8535.4]
  wire [1:0] _GEN_942; // @[Bitwise.scala 48:55:@8536.4]
  wire [2:0] _T_8488; // @[Bitwise.scala 48:55:@8536.4]
  wire [1:0] _T_8489; // @[Bitwise.scala 48:55:@8537.4]
  wire [1:0] _GEN_943; // @[Bitwise.scala 48:55:@8538.4]
  wire [2:0] _T_8490; // @[Bitwise.scala 48:55:@8538.4]
  wire [3:0] _T_8491; // @[Bitwise.scala 48:55:@8539.4]
  wire [1:0] _T_8492; // @[Bitwise.scala 48:55:@8540.4]
  wire [1:0] _GEN_944; // @[Bitwise.scala 48:55:@8541.4]
  wire [2:0] _T_8493; // @[Bitwise.scala 48:55:@8541.4]
  wire [1:0] _T_8494; // @[Bitwise.scala 48:55:@8542.4]
  wire [1:0] _T_8495; // @[Bitwise.scala 48:55:@8543.4]
  wire [2:0] _T_8496; // @[Bitwise.scala 48:55:@8544.4]
  wire [3:0] _T_8497; // @[Bitwise.scala 48:55:@8545.4]
  wire [4:0] _T_8498; // @[Bitwise.scala 48:55:@8546.4]
  wire [1:0] _T_8499; // @[Bitwise.scala 48:55:@8547.4]
  wire [1:0] _GEN_945; // @[Bitwise.scala 48:55:@8548.4]
  wire [2:0] _T_8500; // @[Bitwise.scala 48:55:@8548.4]
  wire [1:0] _T_8501; // @[Bitwise.scala 48:55:@8549.4]
  wire [1:0] _T_8502; // @[Bitwise.scala 48:55:@8550.4]
  wire [2:0] _T_8503; // @[Bitwise.scala 48:55:@8551.4]
  wire [3:0] _T_8504; // @[Bitwise.scala 48:55:@8552.4]
  wire [1:0] _T_8505; // @[Bitwise.scala 48:55:@8553.4]
  wire [1:0] _GEN_946; // @[Bitwise.scala 48:55:@8554.4]
  wire [2:0] _T_8506; // @[Bitwise.scala 48:55:@8554.4]
  wire [1:0] _T_8507; // @[Bitwise.scala 48:55:@8555.4]
  wire [1:0] _T_8508; // @[Bitwise.scala 48:55:@8556.4]
  wire [2:0] _T_8509; // @[Bitwise.scala 48:55:@8557.4]
  wire [3:0] _T_8510; // @[Bitwise.scala 48:55:@8558.4]
  wire [4:0] _T_8511; // @[Bitwise.scala 48:55:@8559.4]
  wire [5:0] _T_8512; // @[Bitwise.scala 48:55:@8560.4]
  wire [1:0] _T_8513; // @[Bitwise.scala 48:55:@8561.4]
  wire [1:0] _GEN_947; // @[Bitwise.scala 48:55:@8562.4]
  wire [2:0] _T_8514; // @[Bitwise.scala 48:55:@8562.4]
  wire [1:0] _T_8515; // @[Bitwise.scala 48:55:@8563.4]
  wire [1:0] _GEN_948; // @[Bitwise.scala 48:55:@8564.4]
  wire [2:0] _T_8516; // @[Bitwise.scala 48:55:@8564.4]
  wire [3:0] _T_8517; // @[Bitwise.scala 48:55:@8565.4]
  wire [1:0] _T_8518; // @[Bitwise.scala 48:55:@8566.4]
  wire [1:0] _GEN_949; // @[Bitwise.scala 48:55:@8567.4]
  wire [2:0] _T_8519; // @[Bitwise.scala 48:55:@8567.4]
  wire [1:0] _T_8520; // @[Bitwise.scala 48:55:@8568.4]
  wire [1:0] _T_8521; // @[Bitwise.scala 48:55:@8569.4]
  wire [2:0] _T_8522; // @[Bitwise.scala 48:55:@8570.4]
  wire [3:0] _T_8523; // @[Bitwise.scala 48:55:@8571.4]
  wire [4:0] _T_8524; // @[Bitwise.scala 48:55:@8572.4]
  wire [1:0] _T_8525; // @[Bitwise.scala 48:55:@8573.4]
  wire [1:0] _GEN_950; // @[Bitwise.scala 48:55:@8574.4]
  wire [2:0] _T_8526; // @[Bitwise.scala 48:55:@8574.4]
  wire [1:0] _T_8527; // @[Bitwise.scala 48:55:@8575.4]
  wire [1:0] _T_8528; // @[Bitwise.scala 48:55:@8576.4]
  wire [2:0] _T_8529; // @[Bitwise.scala 48:55:@8577.4]
  wire [3:0] _T_8530; // @[Bitwise.scala 48:55:@8578.4]
  wire [1:0] _T_8531; // @[Bitwise.scala 48:55:@8579.4]
  wire [1:0] _GEN_951; // @[Bitwise.scala 48:55:@8580.4]
  wire [2:0] _T_8532; // @[Bitwise.scala 48:55:@8580.4]
  wire [1:0] _T_8533; // @[Bitwise.scala 48:55:@8581.4]
  wire [1:0] _T_8534; // @[Bitwise.scala 48:55:@8582.4]
  wire [2:0] _T_8535; // @[Bitwise.scala 48:55:@8583.4]
  wire [3:0] _T_8536; // @[Bitwise.scala 48:55:@8584.4]
  wire [4:0] _T_8537; // @[Bitwise.scala 48:55:@8585.4]
  wire [5:0] _T_8538; // @[Bitwise.scala 48:55:@8586.4]
  wire [6:0] _T_8539; // @[Bitwise.scala 48:55:@8587.4]
  wire [54:0] _T_8603; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@8652.4]
  wire  _T_8604; // @[Bitwise.scala 50:65:@8653.4]
  wire  _T_8605; // @[Bitwise.scala 50:65:@8654.4]
  wire  _T_8606; // @[Bitwise.scala 50:65:@8655.4]
  wire  _T_8607; // @[Bitwise.scala 50:65:@8656.4]
  wire  _T_8608; // @[Bitwise.scala 50:65:@8657.4]
  wire  _T_8609; // @[Bitwise.scala 50:65:@8658.4]
  wire  _T_8610; // @[Bitwise.scala 50:65:@8659.4]
  wire  _T_8611; // @[Bitwise.scala 50:65:@8660.4]
  wire  _T_8612; // @[Bitwise.scala 50:65:@8661.4]
  wire  _T_8613; // @[Bitwise.scala 50:65:@8662.4]
  wire  _T_8614; // @[Bitwise.scala 50:65:@8663.4]
  wire  _T_8615; // @[Bitwise.scala 50:65:@8664.4]
  wire  _T_8616; // @[Bitwise.scala 50:65:@8665.4]
  wire  _T_8617; // @[Bitwise.scala 50:65:@8666.4]
  wire  _T_8618; // @[Bitwise.scala 50:65:@8667.4]
  wire  _T_8619; // @[Bitwise.scala 50:65:@8668.4]
  wire  _T_8620; // @[Bitwise.scala 50:65:@8669.4]
  wire  _T_8621; // @[Bitwise.scala 50:65:@8670.4]
  wire  _T_8622; // @[Bitwise.scala 50:65:@8671.4]
  wire  _T_8623; // @[Bitwise.scala 50:65:@8672.4]
  wire  _T_8624; // @[Bitwise.scala 50:65:@8673.4]
  wire  _T_8625; // @[Bitwise.scala 50:65:@8674.4]
  wire  _T_8626; // @[Bitwise.scala 50:65:@8675.4]
  wire  _T_8627; // @[Bitwise.scala 50:65:@8676.4]
  wire  _T_8628; // @[Bitwise.scala 50:65:@8677.4]
  wire  _T_8629; // @[Bitwise.scala 50:65:@8678.4]
  wire  _T_8630; // @[Bitwise.scala 50:65:@8679.4]
  wire  _T_8631; // @[Bitwise.scala 50:65:@8680.4]
  wire  _T_8632; // @[Bitwise.scala 50:65:@8681.4]
  wire  _T_8633; // @[Bitwise.scala 50:65:@8682.4]
  wire  _T_8634; // @[Bitwise.scala 50:65:@8683.4]
  wire  _T_8635; // @[Bitwise.scala 50:65:@8684.4]
  wire  _T_8636; // @[Bitwise.scala 50:65:@8685.4]
  wire  _T_8637; // @[Bitwise.scala 50:65:@8686.4]
  wire  _T_8638; // @[Bitwise.scala 50:65:@8687.4]
  wire  _T_8639; // @[Bitwise.scala 50:65:@8688.4]
  wire  _T_8640; // @[Bitwise.scala 50:65:@8689.4]
  wire  _T_8641; // @[Bitwise.scala 50:65:@8690.4]
  wire  _T_8642; // @[Bitwise.scala 50:65:@8691.4]
  wire  _T_8643; // @[Bitwise.scala 50:65:@8692.4]
  wire  _T_8644; // @[Bitwise.scala 50:65:@8693.4]
  wire  _T_8645; // @[Bitwise.scala 50:65:@8694.4]
  wire  _T_8646; // @[Bitwise.scala 50:65:@8695.4]
  wire  _T_8647; // @[Bitwise.scala 50:65:@8696.4]
  wire  _T_8648; // @[Bitwise.scala 50:65:@8697.4]
  wire  _T_8649; // @[Bitwise.scala 50:65:@8698.4]
  wire  _T_8650; // @[Bitwise.scala 50:65:@8699.4]
  wire  _T_8651; // @[Bitwise.scala 50:65:@8700.4]
  wire  _T_8652; // @[Bitwise.scala 50:65:@8701.4]
  wire  _T_8653; // @[Bitwise.scala 50:65:@8702.4]
  wire  _T_8654; // @[Bitwise.scala 50:65:@8703.4]
  wire  _T_8655; // @[Bitwise.scala 50:65:@8704.4]
  wire  _T_8656; // @[Bitwise.scala 50:65:@8705.4]
  wire  _T_8657; // @[Bitwise.scala 50:65:@8706.4]
  wire  _T_8658; // @[Bitwise.scala 50:65:@8707.4]
  wire [1:0] _T_8659; // @[Bitwise.scala 48:55:@8708.4]
  wire [1:0] _GEN_952; // @[Bitwise.scala 48:55:@8709.4]
  wire [2:0] _T_8660; // @[Bitwise.scala 48:55:@8709.4]
  wire [1:0] _T_8661; // @[Bitwise.scala 48:55:@8710.4]
  wire [1:0] _GEN_953; // @[Bitwise.scala 48:55:@8711.4]
  wire [2:0] _T_8662; // @[Bitwise.scala 48:55:@8711.4]
  wire [3:0] _T_8663; // @[Bitwise.scala 48:55:@8712.4]
  wire [1:0] _T_8664; // @[Bitwise.scala 48:55:@8713.4]
  wire [1:0] _GEN_954; // @[Bitwise.scala 48:55:@8714.4]
  wire [2:0] _T_8665; // @[Bitwise.scala 48:55:@8714.4]
  wire [1:0] _T_8666; // @[Bitwise.scala 48:55:@8715.4]
  wire [1:0] _T_8667; // @[Bitwise.scala 48:55:@8716.4]
  wire [2:0] _T_8668; // @[Bitwise.scala 48:55:@8717.4]
  wire [3:0] _T_8669; // @[Bitwise.scala 48:55:@8718.4]
  wire [4:0] _T_8670; // @[Bitwise.scala 48:55:@8719.4]
  wire [1:0] _T_8671; // @[Bitwise.scala 48:55:@8720.4]
  wire [1:0] _GEN_955; // @[Bitwise.scala 48:55:@8721.4]
  wire [2:0] _T_8672; // @[Bitwise.scala 48:55:@8721.4]
  wire [1:0] _T_8673; // @[Bitwise.scala 48:55:@8722.4]
  wire [1:0] _T_8674; // @[Bitwise.scala 48:55:@8723.4]
  wire [2:0] _T_8675; // @[Bitwise.scala 48:55:@8724.4]
  wire [3:0] _T_8676; // @[Bitwise.scala 48:55:@8725.4]
  wire [1:0] _T_8677; // @[Bitwise.scala 48:55:@8726.4]
  wire [1:0] _GEN_956; // @[Bitwise.scala 48:55:@8727.4]
  wire [2:0] _T_8678; // @[Bitwise.scala 48:55:@8727.4]
  wire [1:0] _T_8679; // @[Bitwise.scala 48:55:@8728.4]
  wire [1:0] _T_8680; // @[Bitwise.scala 48:55:@8729.4]
  wire [2:0] _T_8681; // @[Bitwise.scala 48:55:@8730.4]
  wire [3:0] _T_8682; // @[Bitwise.scala 48:55:@8731.4]
  wire [4:0] _T_8683; // @[Bitwise.scala 48:55:@8732.4]
  wire [5:0] _T_8684; // @[Bitwise.scala 48:55:@8733.4]
  wire [1:0] _T_8685; // @[Bitwise.scala 48:55:@8734.4]
  wire [1:0] _GEN_957; // @[Bitwise.scala 48:55:@8735.4]
  wire [2:0] _T_8686; // @[Bitwise.scala 48:55:@8735.4]
  wire [1:0] _T_8687; // @[Bitwise.scala 48:55:@8736.4]
  wire [1:0] _T_8688; // @[Bitwise.scala 48:55:@8737.4]
  wire [2:0] _T_8689; // @[Bitwise.scala 48:55:@8738.4]
  wire [3:0] _T_8690; // @[Bitwise.scala 48:55:@8739.4]
  wire [1:0] _T_8691; // @[Bitwise.scala 48:55:@8740.4]
  wire [1:0] _GEN_958; // @[Bitwise.scala 48:55:@8741.4]
  wire [2:0] _T_8692; // @[Bitwise.scala 48:55:@8741.4]
  wire [1:0] _T_8693; // @[Bitwise.scala 48:55:@8742.4]
  wire [1:0] _T_8694; // @[Bitwise.scala 48:55:@8743.4]
  wire [2:0] _T_8695; // @[Bitwise.scala 48:55:@8744.4]
  wire [3:0] _T_8696; // @[Bitwise.scala 48:55:@8745.4]
  wire [4:0] _T_8697; // @[Bitwise.scala 48:55:@8746.4]
  wire [1:0] _T_8698; // @[Bitwise.scala 48:55:@8747.4]
  wire [1:0] _GEN_959; // @[Bitwise.scala 48:55:@8748.4]
  wire [2:0] _T_8699; // @[Bitwise.scala 48:55:@8748.4]
  wire [1:0] _T_8700; // @[Bitwise.scala 48:55:@8749.4]
  wire [1:0] _T_8701; // @[Bitwise.scala 48:55:@8750.4]
  wire [2:0] _T_8702; // @[Bitwise.scala 48:55:@8751.4]
  wire [3:0] _T_8703; // @[Bitwise.scala 48:55:@8752.4]
  wire [1:0] _T_8704; // @[Bitwise.scala 48:55:@8753.4]
  wire [1:0] _GEN_960; // @[Bitwise.scala 48:55:@8754.4]
  wire [2:0] _T_8705; // @[Bitwise.scala 48:55:@8754.4]
  wire [1:0] _T_8706; // @[Bitwise.scala 48:55:@8755.4]
  wire [1:0] _T_8707; // @[Bitwise.scala 48:55:@8756.4]
  wire [2:0] _T_8708; // @[Bitwise.scala 48:55:@8757.4]
  wire [3:0] _T_8709; // @[Bitwise.scala 48:55:@8758.4]
  wire [4:0] _T_8710; // @[Bitwise.scala 48:55:@8759.4]
  wire [5:0] _T_8711; // @[Bitwise.scala 48:55:@8760.4]
  wire [6:0] _T_8712; // @[Bitwise.scala 48:55:@8761.4]
  wire [55:0] _T_8776; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@8826.4]
  wire  _T_8777; // @[Bitwise.scala 50:65:@8827.4]
  wire  _T_8778; // @[Bitwise.scala 50:65:@8828.4]
  wire  _T_8779; // @[Bitwise.scala 50:65:@8829.4]
  wire  _T_8780; // @[Bitwise.scala 50:65:@8830.4]
  wire  _T_8781; // @[Bitwise.scala 50:65:@8831.4]
  wire  _T_8782; // @[Bitwise.scala 50:65:@8832.4]
  wire  _T_8783; // @[Bitwise.scala 50:65:@8833.4]
  wire  _T_8784; // @[Bitwise.scala 50:65:@8834.4]
  wire  _T_8785; // @[Bitwise.scala 50:65:@8835.4]
  wire  _T_8786; // @[Bitwise.scala 50:65:@8836.4]
  wire  _T_8787; // @[Bitwise.scala 50:65:@8837.4]
  wire  _T_8788; // @[Bitwise.scala 50:65:@8838.4]
  wire  _T_8789; // @[Bitwise.scala 50:65:@8839.4]
  wire  _T_8790; // @[Bitwise.scala 50:65:@8840.4]
  wire  _T_8791; // @[Bitwise.scala 50:65:@8841.4]
  wire  _T_8792; // @[Bitwise.scala 50:65:@8842.4]
  wire  _T_8793; // @[Bitwise.scala 50:65:@8843.4]
  wire  _T_8794; // @[Bitwise.scala 50:65:@8844.4]
  wire  _T_8795; // @[Bitwise.scala 50:65:@8845.4]
  wire  _T_8796; // @[Bitwise.scala 50:65:@8846.4]
  wire  _T_8797; // @[Bitwise.scala 50:65:@8847.4]
  wire  _T_8798; // @[Bitwise.scala 50:65:@8848.4]
  wire  _T_8799; // @[Bitwise.scala 50:65:@8849.4]
  wire  _T_8800; // @[Bitwise.scala 50:65:@8850.4]
  wire  _T_8801; // @[Bitwise.scala 50:65:@8851.4]
  wire  _T_8802; // @[Bitwise.scala 50:65:@8852.4]
  wire  _T_8803; // @[Bitwise.scala 50:65:@8853.4]
  wire  _T_8804; // @[Bitwise.scala 50:65:@8854.4]
  wire  _T_8805; // @[Bitwise.scala 50:65:@8855.4]
  wire  _T_8806; // @[Bitwise.scala 50:65:@8856.4]
  wire  _T_8807; // @[Bitwise.scala 50:65:@8857.4]
  wire  _T_8808; // @[Bitwise.scala 50:65:@8858.4]
  wire  _T_8809; // @[Bitwise.scala 50:65:@8859.4]
  wire  _T_8810; // @[Bitwise.scala 50:65:@8860.4]
  wire  _T_8811; // @[Bitwise.scala 50:65:@8861.4]
  wire  _T_8812; // @[Bitwise.scala 50:65:@8862.4]
  wire  _T_8813; // @[Bitwise.scala 50:65:@8863.4]
  wire  _T_8814; // @[Bitwise.scala 50:65:@8864.4]
  wire  _T_8815; // @[Bitwise.scala 50:65:@8865.4]
  wire  _T_8816; // @[Bitwise.scala 50:65:@8866.4]
  wire  _T_8817; // @[Bitwise.scala 50:65:@8867.4]
  wire  _T_8818; // @[Bitwise.scala 50:65:@8868.4]
  wire  _T_8819; // @[Bitwise.scala 50:65:@8869.4]
  wire  _T_8820; // @[Bitwise.scala 50:65:@8870.4]
  wire  _T_8821; // @[Bitwise.scala 50:65:@8871.4]
  wire  _T_8822; // @[Bitwise.scala 50:65:@8872.4]
  wire  _T_8823; // @[Bitwise.scala 50:65:@8873.4]
  wire  _T_8824; // @[Bitwise.scala 50:65:@8874.4]
  wire  _T_8825; // @[Bitwise.scala 50:65:@8875.4]
  wire  _T_8826; // @[Bitwise.scala 50:65:@8876.4]
  wire  _T_8827; // @[Bitwise.scala 50:65:@8877.4]
  wire  _T_8828; // @[Bitwise.scala 50:65:@8878.4]
  wire  _T_8829; // @[Bitwise.scala 50:65:@8879.4]
  wire  _T_8830; // @[Bitwise.scala 50:65:@8880.4]
  wire  _T_8831; // @[Bitwise.scala 50:65:@8881.4]
  wire  _T_8832; // @[Bitwise.scala 50:65:@8882.4]
  wire [1:0] _T_8833; // @[Bitwise.scala 48:55:@8883.4]
  wire [1:0] _GEN_961; // @[Bitwise.scala 48:55:@8884.4]
  wire [2:0] _T_8834; // @[Bitwise.scala 48:55:@8884.4]
  wire [1:0] _T_8835; // @[Bitwise.scala 48:55:@8885.4]
  wire [1:0] _T_8836; // @[Bitwise.scala 48:55:@8886.4]
  wire [2:0] _T_8837; // @[Bitwise.scala 48:55:@8887.4]
  wire [3:0] _T_8838; // @[Bitwise.scala 48:55:@8888.4]
  wire [1:0] _T_8839; // @[Bitwise.scala 48:55:@8889.4]
  wire [1:0] _GEN_962; // @[Bitwise.scala 48:55:@8890.4]
  wire [2:0] _T_8840; // @[Bitwise.scala 48:55:@8890.4]
  wire [1:0] _T_8841; // @[Bitwise.scala 48:55:@8891.4]
  wire [1:0] _T_8842; // @[Bitwise.scala 48:55:@8892.4]
  wire [2:0] _T_8843; // @[Bitwise.scala 48:55:@8893.4]
  wire [3:0] _T_8844; // @[Bitwise.scala 48:55:@8894.4]
  wire [4:0] _T_8845; // @[Bitwise.scala 48:55:@8895.4]
  wire [1:0] _T_8846; // @[Bitwise.scala 48:55:@8896.4]
  wire [1:0] _GEN_963; // @[Bitwise.scala 48:55:@8897.4]
  wire [2:0] _T_8847; // @[Bitwise.scala 48:55:@8897.4]
  wire [1:0] _T_8848; // @[Bitwise.scala 48:55:@8898.4]
  wire [1:0] _T_8849; // @[Bitwise.scala 48:55:@8899.4]
  wire [2:0] _T_8850; // @[Bitwise.scala 48:55:@8900.4]
  wire [3:0] _T_8851; // @[Bitwise.scala 48:55:@8901.4]
  wire [1:0] _T_8852; // @[Bitwise.scala 48:55:@8902.4]
  wire [1:0] _GEN_964; // @[Bitwise.scala 48:55:@8903.4]
  wire [2:0] _T_8853; // @[Bitwise.scala 48:55:@8903.4]
  wire [1:0] _T_8854; // @[Bitwise.scala 48:55:@8904.4]
  wire [1:0] _T_8855; // @[Bitwise.scala 48:55:@8905.4]
  wire [2:0] _T_8856; // @[Bitwise.scala 48:55:@8906.4]
  wire [3:0] _T_8857; // @[Bitwise.scala 48:55:@8907.4]
  wire [4:0] _T_8858; // @[Bitwise.scala 48:55:@8908.4]
  wire [5:0] _T_8859; // @[Bitwise.scala 48:55:@8909.4]
  wire [1:0] _T_8860; // @[Bitwise.scala 48:55:@8910.4]
  wire [1:0] _GEN_965; // @[Bitwise.scala 48:55:@8911.4]
  wire [2:0] _T_8861; // @[Bitwise.scala 48:55:@8911.4]
  wire [1:0] _T_8862; // @[Bitwise.scala 48:55:@8912.4]
  wire [1:0] _T_8863; // @[Bitwise.scala 48:55:@8913.4]
  wire [2:0] _T_8864; // @[Bitwise.scala 48:55:@8914.4]
  wire [3:0] _T_8865; // @[Bitwise.scala 48:55:@8915.4]
  wire [1:0] _T_8866; // @[Bitwise.scala 48:55:@8916.4]
  wire [1:0] _GEN_966; // @[Bitwise.scala 48:55:@8917.4]
  wire [2:0] _T_8867; // @[Bitwise.scala 48:55:@8917.4]
  wire [1:0] _T_8868; // @[Bitwise.scala 48:55:@8918.4]
  wire [1:0] _T_8869; // @[Bitwise.scala 48:55:@8919.4]
  wire [2:0] _T_8870; // @[Bitwise.scala 48:55:@8920.4]
  wire [3:0] _T_8871; // @[Bitwise.scala 48:55:@8921.4]
  wire [4:0] _T_8872; // @[Bitwise.scala 48:55:@8922.4]
  wire [1:0] _T_8873; // @[Bitwise.scala 48:55:@8923.4]
  wire [1:0] _GEN_967; // @[Bitwise.scala 48:55:@8924.4]
  wire [2:0] _T_8874; // @[Bitwise.scala 48:55:@8924.4]
  wire [1:0] _T_8875; // @[Bitwise.scala 48:55:@8925.4]
  wire [1:0] _T_8876; // @[Bitwise.scala 48:55:@8926.4]
  wire [2:0] _T_8877; // @[Bitwise.scala 48:55:@8927.4]
  wire [3:0] _T_8878; // @[Bitwise.scala 48:55:@8928.4]
  wire [1:0] _T_8879; // @[Bitwise.scala 48:55:@8929.4]
  wire [1:0] _GEN_968; // @[Bitwise.scala 48:55:@8930.4]
  wire [2:0] _T_8880; // @[Bitwise.scala 48:55:@8930.4]
  wire [1:0] _T_8881; // @[Bitwise.scala 48:55:@8931.4]
  wire [1:0] _T_8882; // @[Bitwise.scala 48:55:@8932.4]
  wire [2:0] _T_8883; // @[Bitwise.scala 48:55:@8933.4]
  wire [3:0] _T_8884; // @[Bitwise.scala 48:55:@8934.4]
  wire [4:0] _T_8885; // @[Bitwise.scala 48:55:@8935.4]
  wire [5:0] _T_8886; // @[Bitwise.scala 48:55:@8936.4]
  wire [6:0] _T_8887; // @[Bitwise.scala 48:55:@8937.4]
  wire [56:0] _T_8951; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@9002.4]
  wire  _T_8952; // @[Bitwise.scala 50:65:@9003.4]
  wire  _T_8953; // @[Bitwise.scala 50:65:@9004.4]
  wire  _T_8954; // @[Bitwise.scala 50:65:@9005.4]
  wire  _T_8955; // @[Bitwise.scala 50:65:@9006.4]
  wire  _T_8956; // @[Bitwise.scala 50:65:@9007.4]
  wire  _T_8957; // @[Bitwise.scala 50:65:@9008.4]
  wire  _T_8958; // @[Bitwise.scala 50:65:@9009.4]
  wire  _T_8959; // @[Bitwise.scala 50:65:@9010.4]
  wire  _T_8960; // @[Bitwise.scala 50:65:@9011.4]
  wire  _T_8961; // @[Bitwise.scala 50:65:@9012.4]
  wire  _T_8962; // @[Bitwise.scala 50:65:@9013.4]
  wire  _T_8963; // @[Bitwise.scala 50:65:@9014.4]
  wire  _T_8964; // @[Bitwise.scala 50:65:@9015.4]
  wire  _T_8965; // @[Bitwise.scala 50:65:@9016.4]
  wire  _T_8966; // @[Bitwise.scala 50:65:@9017.4]
  wire  _T_8967; // @[Bitwise.scala 50:65:@9018.4]
  wire  _T_8968; // @[Bitwise.scala 50:65:@9019.4]
  wire  _T_8969; // @[Bitwise.scala 50:65:@9020.4]
  wire  _T_8970; // @[Bitwise.scala 50:65:@9021.4]
  wire  _T_8971; // @[Bitwise.scala 50:65:@9022.4]
  wire  _T_8972; // @[Bitwise.scala 50:65:@9023.4]
  wire  _T_8973; // @[Bitwise.scala 50:65:@9024.4]
  wire  _T_8974; // @[Bitwise.scala 50:65:@9025.4]
  wire  _T_8975; // @[Bitwise.scala 50:65:@9026.4]
  wire  _T_8976; // @[Bitwise.scala 50:65:@9027.4]
  wire  _T_8977; // @[Bitwise.scala 50:65:@9028.4]
  wire  _T_8978; // @[Bitwise.scala 50:65:@9029.4]
  wire  _T_8979; // @[Bitwise.scala 50:65:@9030.4]
  wire  _T_8980; // @[Bitwise.scala 50:65:@9031.4]
  wire  _T_8981; // @[Bitwise.scala 50:65:@9032.4]
  wire  _T_8982; // @[Bitwise.scala 50:65:@9033.4]
  wire  _T_8983; // @[Bitwise.scala 50:65:@9034.4]
  wire  _T_8984; // @[Bitwise.scala 50:65:@9035.4]
  wire  _T_8985; // @[Bitwise.scala 50:65:@9036.4]
  wire  _T_8986; // @[Bitwise.scala 50:65:@9037.4]
  wire  _T_8987; // @[Bitwise.scala 50:65:@9038.4]
  wire  _T_8988; // @[Bitwise.scala 50:65:@9039.4]
  wire  _T_8989; // @[Bitwise.scala 50:65:@9040.4]
  wire  _T_8990; // @[Bitwise.scala 50:65:@9041.4]
  wire  _T_8991; // @[Bitwise.scala 50:65:@9042.4]
  wire  _T_8992; // @[Bitwise.scala 50:65:@9043.4]
  wire  _T_8993; // @[Bitwise.scala 50:65:@9044.4]
  wire  _T_8994; // @[Bitwise.scala 50:65:@9045.4]
  wire  _T_8995; // @[Bitwise.scala 50:65:@9046.4]
  wire  _T_8996; // @[Bitwise.scala 50:65:@9047.4]
  wire  _T_8997; // @[Bitwise.scala 50:65:@9048.4]
  wire  _T_8998; // @[Bitwise.scala 50:65:@9049.4]
  wire  _T_8999; // @[Bitwise.scala 50:65:@9050.4]
  wire  _T_9000; // @[Bitwise.scala 50:65:@9051.4]
  wire  _T_9001; // @[Bitwise.scala 50:65:@9052.4]
  wire  _T_9002; // @[Bitwise.scala 50:65:@9053.4]
  wire  _T_9003; // @[Bitwise.scala 50:65:@9054.4]
  wire  _T_9004; // @[Bitwise.scala 50:65:@9055.4]
  wire  _T_9005; // @[Bitwise.scala 50:65:@9056.4]
  wire  _T_9006; // @[Bitwise.scala 50:65:@9057.4]
  wire  _T_9007; // @[Bitwise.scala 50:65:@9058.4]
  wire  _T_9008; // @[Bitwise.scala 50:65:@9059.4]
  wire [1:0] _T_9009; // @[Bitwise.scala 48:55:@9060.4]
  wire [1:0] _GEN_969; // @[Bitwise.scala 48:55:@9061.4]
  wire [2:0] _T_9010; // @[Bitwise.scala 48:55:@9061.4]
  wire [1:0] _T_9011; // @[Bitwise.scala 48:55:@9062.4]
  wire [1:0] _T_9012; // @[Bitwise.scala 48:55:@9063.4]
  wire [2:0] _T_9013; // @[Bitwise.scala 48:55:@9064.4]
  wire [3:0] _T_9014; // @[Bitwise.scala 48:55:@9065.4]
  wire [1:0] _T_9015; // @[Bitwise.scala 48:55:@9066.4]
  wire [1:0] _GEN_970; // @[Bitwise.scala 48:55:@9067.4]
  wire [2:0] _T_9016; // @[Bitwise.scala 48:55:@9067.4]
  wire [1:0] _T_9017; // @[Bitwise.scala 48:55:@9068.4]
  wire [1:0] _T_9018; // @[Bitwise.scala 48:55:@9069.4]
  wire [2:0] _T_9019; // @[Bitwise.scala 48:55:@9070.4]
  wire [3:0] _T_9020; // @[Bitwise.scala 48:55:@9071.4]
  wire [4:0] _T_9021; // @[Bitwise.scala 48:55:@9072.4]
  wire [1:0] _T_9022; // @[Bitwise.scala 48:55:@9073.4]
  wire [1:0] _GEN_971; // @[Bitwise.scala 48:55:@9074.4]
  wire [2:0] _T_9023; // @[Bitwise.scala 48:55:@9074.4]
  wire [1:0] _T_9024; // @[Bitwise.scala 48:55:@9075.4]
  wire [1:0] _T_9025; // @[Bitwise.scala 48:55:@9076.4]
  wire [2:0] _T_9026; // @[Bitwise.scala 48:55:@9077.4]
  wire [3:0] _T_9027; // @[Bitwise.scala 48:55:@9078.4]
  wire [1:0] _T_9028; // @[Bitwise.scala 48:55:@9079.4]
  wire [1:0] _GEN_972; // @[Bitwise.scala 48:55:@9080.4]
  wire [2:0] _T_9029; // @[Bitwise.scala 48:55:@9080.4]
  wire [1:0] _T_9030; // @[Bitwise.scala 48:55:@9081.4]
  wire [1:0] _T_9031; // @[Bitwise.scala 48:55:@9082.4]
  wire [2:0] _T_9032; // @[Bitwise.scala 48:55:@9083.4]
  wire [3:0] _T_9033; // @[Bitwise.scala 48:55:@9084.4]
  wire [4:0] _T_9034; // @[Bitwise.scala 48:55:@9085.4]
  wire [5:0] _T_9035; // @[Bitwise.scala 48:55:@9086.4]
  wire [1:0] _T_9036; // @[Bitwise.scala 48:55:@9087.4]
  wire [1:0] _GEN_973; // @[Bitwise.scala 48:55:@9088.4]
  wire [2:0] _T_9037; // @[Bitwise.scala 48:55:@9088.4]
  wire [1:0] _T_9038; // @[Bitwise.scala 48:55:@9089.4]
  wire [1:0] _T_9039; // @[Bitwise.scala 48:55:@9090.4]
  wire [2:0] _T_9040; // @[Bitwise.scala 48:55:@9091.4]
  wire [3:0] _T_9041; // @[Bitwise.scala 48:55:@9092.4]
  wire [1:0] _T_9042; // @[Bitwise.scala 48:55:@9093.4]
  wire [1:0] _GEN_974; // @[Bitwise.scala 48:55:@9094.4]
  wire [2:0] _T_9043; // @[Bitwise.scala 48:55:@9094.4]
  wire [1:0] _T_9044; // @[Bitwise.scala 48:55:@9095.4]
  wire [1:0] _T_9045; // @[Bitwise.scala 48:55:@9096.4]
  wire [2:0] _T_9046; // @[Bitwise.scala 48:55:@9097.4]
  wire [3:0] _T_9047; // @[Bitwise.scala 48:55:@9098.4]
  wire [4:0] _T_9048; // @[Bitwise.scala 48:55:@9099.4]
  wire [1:0] _T_9049; // @[Bitwise.scala 48:55:@9100.4]
  wire [1:0] _GEN_975; // @[Bitwise.scala 48:55:@9101.4]
  wire [2:0] _T_9050; // @[Bitwise.scala 48:55:@9101.4]
  wire [1:0] _T_9051; // @[Bitwise.scala 48:55:@9102.4]
  wire [1:0] _T_9052; // @[Bitwise.scala 48:55:@9103.4]
  wire [2:0] _T_9053; // @[Bitwise.scala 48:55:@9104.4]
  wire [3:0] _T_9054; // @[Bitwise.scala 48:55:@9105.4]
  wire [1:0] _T_9055; // @[Bitwise.scala 48:55:@9106.4]
  wire [1:0] _T_9056; // @[Bitwise.scala 48:55:@9107.4]
  wire [2:0] _T_9057; // @[Bitwise.scala 48:55:@9108.4]
  wire [1:0] _T_9058; // @[Bitwise.scala 48:55:@9109.4]
  wire [1:0] _T_9059; // @[Bitwise.scala 48:55:@9110.4]
  wire [2:0] _T_9060; // @[Bitwise.scala 48:55:@9111.4]
  wire [3:0] _T_9061; // @[Bitwise.scala 48:55:@9112.4]
  wire [4:0] _T_9062; // @[Bitwise.scala 48:55:@9113.4]
  wire [5:0] _T_9063; // @[Bitwise.scala 48:55:@9114.4]
  wire [6:0] _T_9064; // @[Bitwise.scala 48:55:@9115.4]
  wire [57:0] _T_9128; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@9180.4]
  wire  _T_9129; // @[Bitwise.scala 50:65:@9181.4]
  wire  _T_9130; // @[Bitwise.scala 50:65:@9182.4]
  wire  _T_9131; // @[Bitwise.scala 50:65:@9183.4]
  wire  _T_9132; // @[Bitwise.scala 50:65:@9184.4]
  wire  _T_9133; // @[Bitwise.scala 50:65:@9185.4]
  wire  _T_9134; // @[Bitwise.scala 50:65:@9186.4]
  wire  _T_9135; // @[Bitwise.scala 50:65:@9187.4]
  wire  _T_9136; // @[Bitwise.scala 50:65:@9188.4]
  wire  _T_9137; // @[Bitwise.scala 50:65:@9189.4]
  wire  _T_9138; // @[Bitwise.scala 50:65:@9190.4]
  wire  _T_9139; // @[Bitwise.scala 50:65:@9191.4]
  wire  _T_9140; // @[Bitwise.scala 50:65:@9192.4]
  wire  _T_9141; // @[Bitwise.scala 50:65:@9193.4]
  wire  _T_9142; // @[Bitwise.scala 50:65:@9194.4]
  wire  _T_9143; // @[Bitwise.scala 50:65:@9195.4]
  wire  _T_9144; // @[Bitwise.scala 50:65:@9196.4]
  wire  _T_9145; // @[Bitwise.scala 50:65:@9197.4]
  wire  _T_9146; // @[Bitwise.scala 50:65:@9198.4]
  wire  _T_9147; // @[Bitwise.scala 50:65:@9199.4]
  wire  _T_9148; // @[Bitwise.scala 50:65:@9200.4]
  wire  _T_9149; // @[Bitwise.scala 50:65:@9201.4]
  wire  _T_9150; // @[Bitwise.scala 50:65:@9202.4]
  wire  _T_9151; // @[Bitwise.scala 50:65:@9203.4]
  wire  _T_9152; // @[Bitwise.scala 50:65:@9204.4]
  wire  _T_9153; // @[Bitwise.scala 50:65:@9205.4]
  wire  _T_9154; // @[Bitwise.scala 50:65:@9206.4]
  wire  _T_9155; // @[Bitwise.scala 50:65:@9207.4]
  wire  _T_9156; // @[Bitwise.scala 50:65:@9208.4]
  wire  _T_9157; // @[Bitwise.scala 50:65:@9209.4]
  wire  _T_9158; // @[Bitwise.scala 50:65:@9210.4]
  wire  _T_9159; // @[Bitwise.scala 50:65:@9211.4]
  wire  _T_9160; // @[Bitwise.scala 50:65:@9212.4]
  wire  _T_9161; // @[Bitwise.scala 50:65:@9213.4]
  wire  _T_9162; // @[Bitwise.scala 50:65:@9214.4]
  wire  _T_9163; // @[Bitwise.scala 50:65:@9215.4]
  wire  _T_9164; // @[Bitwise.scala 50:65:@9216.4]
  wire  _T_9165; // @[Bitwise.scala 50:65:@9217.4]
  wire  _T_9166; // @[Bitwise.scala 50:65:@9218.4]
  wire  _T_9167; // @[Bitwise.scala 50:65:@9219.4]
  wire  _T_9168; // @[Bitwise.scala 50:65:@9220.4]
  wire  _T_9169; // @[Bitwise.scala 50:65:@9221.4]
  wire  _T_9170; // @[Bitwise.scala 50:65:@9222.4]
  wire  _T_9171; // @[Bitwise.scala 50:65:@9223.4]
  wire  _T_9172; // @[Bitwise.scala 50:65:@9224.4]
  wire  _T_9173; // @[Bitwise.scala 50:65:@9225.4]
  wire  _T_9174; // @[Bitwise.scala 50:65:@9226.4]
  wire  _T_9175; // @[Bitwise.scala 50:65:@9227.4]
  wire  _T_9176; // @[Bitwise.scala 50:65:@9228.4]
  wire  _T_9177; // @[Bitwise.scala 50:65:@9229.4]
  wire  _T_9178; // @[Bitwise.scala 50:65:@9230.4]
  wire  _T_9179; // @[Bitwise.scala 50:65:@9231.4]
  wire  _T_9180; // @[Bitwise.scala 50:65:@9232.4]
  wire  _T_9181; // @[Bitwise.scala 50:65:@9233.4]
  wire  _T_9182; // @[Bitwise.scala 50:65:@9234.4]
  wire  _T_9183; // @[Bitwise.scala 50:65:@9235.4]
  wire  _T_9184; // @[Bitwise.scala 50:65:@9236.4]
  wire  _T_9185; // @[Bitwise.scala 50:65:@9237.4]
  wire  _T_9186; // @[Bitwise.scala 50:65:@9238.4]
  wire [1:0] _T_9187; // @[Bitwise.scala 48:55:@9239.4]
  wire [1:0] _GEN_976; // @[Bitwise.scala 48:55:@9240.4]
  wire [2:0] _T_9188; // @[Bitwise.scala 48:55:@9240.4]
  wire [1:0] _T_9189; // @[Bitwise.scala 48:55:@9241.4]
  wire [1:0] _T_9190; // @[Bitwise.scala 48:55:@9242.4]
  wire [2:0] _T_9191; // @[Bitwise.scala 48:55:@9243.4]
  wire [3:0] _T_9192; // @[Bitwise.scala 48:55:@9244.4]
  wire [1:0] _T_9193; // @[Bitwise.scala 48:55:@9245.4]
  wire [1:0] _GEN_977; // @[Bitwise.scala 48:55:@9246.4]
  wire [2:0] _T_9194; // @[Bitwise.scala 48:55:@9246.4]
  wire [1:0] _T_9195; // @[Bitwise.scala 48:55:@9247.4]
  wire [1:0] _T_9196; // @[Bitwise.scala 48:55:@9248.4]
  wire [2:0] _T_9197; // @[Bitwise.scala 48:55:@9249.4]
  wire [3:0] _T_9198; // @[Bitwise.scala 48:55:@9250.4]
  wire [4:0] _T_9199; // @[Bitwise.scala 48:55:@9251.4]
  wire [1:0] _T_9200; // @[Bitwise.scala 48:55:@9252.4]
  wire [1:0] _GEN_978; // @[Bitwise.scala 48:55:@9253.4]
  wire [2:0] _T_9201; // @[Bitwise.scala 48:55:@9253.4]
  wire [1:0] _T_9202; // @[Bitwise.scala 48:55:@9254.4]
  wire [1:0] _T_9203; // @[Bitwise.scala 48:55:@9255.4]
  wire [2:0] _T_9204; // @[Bitwise.scala 48:55:@9256.4]
  wire [3:0] _T_9205; // @[Bitwise.scala 48:55:@9257.4]
  wire [1:0] _T_9206; // @[Bitwise.scala 48:55:@9258.4]
  wire [1:0] _T_9207; // @[Bitwise.scala 48:55:@9259.4]
  wire [2:0] _T_9208; // @[Bitwise.scala 48:55:@9260.4]
  wire [1:0] _T_9209; // @[Bitwise.scala 48:55:@9261.4]
  wire [1:0] _T_9210; // @[Bitwise.scala 48:55:@9262.4]
  wire [2:0] _T_9211; // @[Bitwise.scala 48:55:@9263.4]
  wire [3:0] _T_9212; // @[Bitwise.scala 48:55:@9264.4]
  wire [4:0] _T_9213; // @[Bitwise.scala 48:55:@9265.4]
  wire [5:0] _T_9214; // @[Bitwise.scala 48:55:@9266.4]
  wire [1:0] _T_9215; // @[Bitwise.scala 48:55:@9267.4]
  wire [1:0] _GEN_979; // @[Bitwise.scala 48:55:@9268.4]
  wire [2:0] _T_9216; // @[Bitwise.scala 48:55:@9268.4]
  wire [1:0] _T_9217; // @[Bitwise.scala 48:55:@9269.4]
  wire [1:0] _T_9218; // @[Bitwise.scala 48:55:@9270.4]
  wire [2:0] _T_9219; // @[Bitwise.scala 48:55:@9271.4]
  wire [3:0] _T_9220; // @[Bitwise.scala 48:55:@9272.4]
  wire [1:0] _T_9221; // @[Bitwise.scala 48:55:@9273.4]
  wire [1:0] _GEN_980; // @[Bitwise.scala 48:55:@9274.4]
  wire [2:0] _T_9222; // @[Bitwise.scala 48:55:@9274.4]
  wire [1:0] _T_9223; // @[Bitwise.scala 48:55:@9275.4]
  wire [1:0] _T_9224; // @[Bitwise.scala 48:55:@9276.4]
  wire [2:0] _T_9225; // @[Bitwise.scala 48:55:@9277.4]
  wire [3:0] _T_9226; // @[Bitwise.scala 48:55:@9278.4]
  wire [4:0] _T_9227; // @[Bitwise.scala 48:55:@9279.4]
  wire [1:0] _T_9228; // @[Bitwise.scala 48:55:@9280.4]
  wire [1:0] _GEN_981; // @[Bitwise.scala 48:55:@9281.4]
  wire [2:0] _T_9229; // @[Bitwise.scala 48:55:@9281.4]
  wire [1:0] _T_9230; // @[Bitwise.scala 48:55:@9282.4]
  wire [1:0] _T_9231; // @[Bitwise.scala 48:55:@9283.4]
  wire [2:0] _T_9232; // @[Bitwise.scala 48:55:@9284.4]
  wire [3:0] _T_9233; // @[Bitwise.scala 48:55:@9285.4]
  wire [1:0] _T_9234; // @[Bitwise.scala 48:55:@9286.4]
  wire [1:0] _T_9235; // @[Bitwise.scala 48:55:@9287.4]
  wire [2:0] _T_9236; // @[Bitwise.scala 48:55:@9288.4]
  wire [1:0] _T_9237; // @[Bitwise.scala 48:55:@9289.4]
  wire [1:0] _T_9238; // @[Bitwise.scala 48:55:@9290.4]
  wire [2:0] _T_9239; // @[Bitwise.scala 48:55:@9291.4]
  wire [3:0] _T_9240; // @[Bitwise.scala 48:55:@9292.4]
  wire [4:0] _T_9241; // @[Bitwise.scala 48:55:@9293.4]
  wire [5:0] _T_9242; // @[Bitwise.scala 48:55:@9294.4]
  wire [6:0] _T_9243; // @[Bitwise.scala 48:55:@9295.4]
  wire [58:0] _T_9307; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@9360.4]
  wire  _T_9308; // @[Bitwise.scala 50:65:@9361.4]
  wire  _T_9309; // @[Bitwise.scala 50:65:@9362.4]
  wire  _T_9310; // @[Bitwise.scala 50:65:@9363.4]
  wire  _T_9311; // @[Bitwise.scala 50:65:@9364.4]
  wire  _T_9312; // @[Bitwise.scala 50:65:@9365.4]
  wire  _T_9313; // @[Bitwise.scala 50:65:@9366.4]
  wire  _T_9314; // @[Bitwise.scala 50:65:@9367.4]
  wire  _T_9315; // @[Bitwise.scala 50:65:@9368.4]
  wire  _T_9316; // @[Bitwise.scala 50:65:@9369.4]
  wire  _T_9317; // @[Bitwise.scala 50:65:@9370.4]
  wire  _T_9318; // @[Bitwise.scala 50:65:@9371.4]
  wire  _T_9319; // @[Bitwise.scala 50:65:@9372.4]
  wire  _T_9320; // @[Bitwise.scala 50:65:@9373.4]
  wire  _T_9321; // @[Bitwise.scala 50:65:@9374.4]
  wire  _T_9322; // @[Bitwise.scala 50:65:@9375.4]
  wire  _T_9323; // @[Bitwise.scala 50:65:@9376.4]
  wire  _T_9324; // @[Bitwise.scala 50:65:@9377.4]
  wire  _T_9325; // @[Bitwise.scala 50:65:@9378.4]
  wire  _T_9326; // @[Bitwise.scala 50:65:@9379.4]
  wire  _T_9327; // @[Bitwise.scala 50:65:@9380.4]
  wire  _T_9328; // @[Bitwise.scala 50:65:@9381.4]
  wire  _T_9329; // @[Bitwise.scala 50:65:@9382.4]
  wire  _T_9330; // @[Bitwise.scala 50:65:@9383.4]
  wire  _T_9331; // @[Bitwise.scala 50:65:@9384.4]
  wire  _T_9332; // @[Bitwise.scala 50:65:@9385.4]
  wire  _T_9333; // @[Bitwise.scala 50:65:@9386.4]
  wire  _T_9334; // @[Bitwise.scala 50:65:@9387.4]
  wire  _T_9335; // @[Bitwise.scala 50:65:@9388.4]
  wire  _T_9336; // @[Bitwise.scala 50:65:@9389.4]
  wire  _T_9337; // @[Bitwise.scala 50:65:@9390.4]
  wire  _T_9338; // @[Bitwise.scala 50:65:@9391.4]
  wire  _T_9339; // @[Bitwise.scala 50:65:@9392.4]
  wire  _T_9340; // @[Bitwise.scala 50:65:@9393.4]
  wire  _T_9341; // @[Bitwise.scala 50:65:@9394.4]
  wire  _T_9342; // @[Bitwise.scala 50:65:@9395.4]
  wire  _T_9343; // @[Bitwise.scala 50:65:@9396.4]
  wire  _T_9344; // @[Bitwise.scala 50:65:@9397.4]
  wire  _T_9345; // @[Bitwise.scala 50:65:@9398.4]
  wire  _T_9346; // @[Bitwise.scala 50:65:@9399.4]
  wire  _T_9347; // @[Bitwise.scala 50:65:@9400.4]
  wire  _T_9348; // @[Bitwise.scala 50:65:@9401.4]
  wire  _T_9349; // @[Bitwise.scala 50:65:@9402.4]
  wire  _T_9350; // @[Bitwise.scala 50:65:@9403.4]
  wire  _T_9351; // @[Bitwise.scala 50:65:@9404.4]
  wire  _T_9352; // @[Bitwise.scala 50:65:@9405.4]
  wire  _T_9353; // @[Bitwise.scala 50:65:@9406.4]
  wire  _T_9354; // @[Bitwise.scala 50:65:@9407.4]
  wire  _T_9355; // @[Bitwise.scala 50:65:@9408.4]
  wire  _T_9356; // @[Bitwise.scala 50:65:@9409.4]
  wire  _T_9357; // @[Bitwise.scala 50:65:@9410.4]
  wire  _T_9358; // @[Bitwise.scala 50:65:@9411.4]
  wire  _T_9359; // @[Bitwise.scala 50:65:@9412.4]
  wire  _T_9360; // @[Bitwise.scala 50:65:@9413.4]
  wire  _T_9361; // @[Bitwise.scala 50:65:@9414.4]
  wire  _T_9362; // @[Bitwise.scala 50:65:@9415.4]
  wire  _T_9363; // @[Bitwise.scala 50:65:@9416.4]
  wire  _T_9364; // @[Bitwise.scala 50:65:@9417.4]
  wire  _T_9365; // @[Bitwise.scala 50:65:@9418.4]
  wire  _T_9366; // @[Bitwise.scala 50:65:@9419.4]
  wire [1:0] _T_9367; // @[Bitwise.scala 48:55:@9420.4]
  wire [1:0] _GEN_982; // @[Bitwise.scala 48:55:@9421.4]
  wire [2:0] _T_9368; // @[Bitwise.scala 48:55:@9421.4]
  wire [1:0] _T_9369; // @[Bitwise.scala 48:55:@9422.4]
  wire [1:0] _T_9370; // @[Bitwise.scala 48:55:@9423.4]
  wire [2:0] _T_9371; // @[Bitwise.scala 48:55:@9424.4]
  wire [3:0] _T_9372; // @[Bitwise.scala 48:55:@9425.4]
  wire [1:0] _T_9373; // @[Bitwise.scala 48:55:@9426.4]
  wire [1:0] _GEN_983; // @[Bitwise.scala 48:55:@9427.4]
  wire [2:0] _T_9374; // @[Bitwise.scala 48:55:@9427.4]
  wire [1:0] _T_9375; // @[Bitwise.scala 48:55:@9428.4]
  wire [1:0] _T_9376; // @[Bitwise.scala 48:55:@9429.4]
  wire [2:0] _T_9377; // @[Bitwise.scala 48:55:@9430.4]
  wire [3:0] _T_9378; // @[Bitwise.scala 48:55:@9431.4]
  wire [4:0] _T_9379; // @[Bitwise.scala 48:55:@9432.4]
  wire [1:0] _T_9380; // @[Bitwise.scala 48:55:@9433.4]
  wire [1:0] _GEN_984; // @[Bitwise.scala 48:55:@9434.4]
  wire [2:0] _T_9381; // @[Bitwise.scala 48:55:@9434.4]
  wire [1:0] _T_9382; // @[Bitwise.scala 48:55:@9435.4]
  wire [1:0] _T_9383; // @[Bitwise.scala 48:55:@9436.4]
  wire [2:0] _T_9384; // @[Bitwise.scala 48:55:@9437.4]
  wire [3:0] _T_9385; // @[Bitwise.scala 48:55:@9438.4]
  wire [1:0] _T_9386; // @[Bitwise.scala 48:55:@9439.4]
  wire [1:0] _T_9387; // @[Bitwise.scala 48:55:@9440.4]
  wire [2:0] _T_9388; // @[Bitwise.scala 48:55:@9441.4]
  wire [1:0] _T_9389; // @[Bitwise.scala 48:55:@9442.4]
  wire [1:0] _T_9390; // @[Bitwise.scala 48:55:@9443.4]
  wire [2:0] _T_9391; // @[Bitwise.scala 48:55:@9444.4]
  wire [3:0] _T_9392; // @[Bitwise.scala 48:55:@9445.4]
  wire [4:0] _T_9393; // @[Bitwise.scala 48:55:@9446.4]
  wire [5:0] _T_9394; // @[Bitwise.scala 48:55:@9447.4]
  wire [1:0] _T_9395; // @[Bitwise.scala 48:55:@9448.4]
  wire [1:0] _GEN_985; // @[Bitwise.scala 48:55:@9449.4]
  wire [2:0] _T_9396; // @[Bitwise.scala 48:55:@9449.4]
  wire [1:0] _T_9397; // @[Bitwise.scala 48:55:@9450.4]
  wire [1:0] _T_9398; // @[Bitwise.scala 48:55:@9451.4]
  wire [2:0] _T_9399; // @[Bitwise.scala 48:55:@9452.4]
  wire [3:0] _T_9400; // @[Bitwise.scala 48:55:@9453.4]
  wire [1:0] _T_9401; // @[Bitwise.scala 48:55:@9454.4]
  wire [1:0] _T_9402; // @[Bitwise.scala 48:55:@9455.4]
  wire [2:0] _T_9403; // @[Bitwise.scala 48:55:@9456.4]
  wire [1:0] _T_9404; // @[Bitwise.scala 48:55:@9457.4]
  wire [1:0] _T_9405; // @[Bitwise.scala 48:55:@9458.4]
  wire [2:0] _T_9406; // @[Bitwise.scala 48:55:@9459.4]
  wire [3:0] _T_9407; // @[Bitwise.scala 48:55:@9460.4]
  wire [4:0] _T_9408; // @[Bitwise.scala 48:55:@9461.4]
  wire [1:0] _T_9409; // @[Bitwise.scala 48:55:@9462.4]
  wire [1:0] _GEN_986; // @[Bitwise.scala 48:55:@9463.4]
  wire [2:0] _T_9410; // @[Bitwise.scala 48:55:@9463.4]
  wire [1:0] _T_9411; // @[Bitwise.scala 48:55:@9464.4]
  wire [1:0] _T_9412; // @[Bitwise.scala 48:55:@9465.4]
  wire [2:0] _T_9413; // @[Bitwise.scala 48:55:@9466.4]
  wire [3:0] _T_9414; // @[Bitwise.scala 48:55:@9467.4]
  wire [1:0] _T_9415; // @[Bitwise.scala 48:55:@9468.4]
  wire [1:0] _T_9416; // @[Bitwise.scala 48:55:@9469.4]
  wire [2:0] _T_9417; // @[Bitwise.scala 48:55:@9470.4]
  wire [1:0] _T_9418; // @[Bitwise.scala 48:55:@9471.4]
  wire [1:0] _T_9419; // @[Bitwise.scala 48:55:@9472.4]
  wire [2:0] _T_9420; // @[Bitwise.scala 48:55:@9473.4]
  wire [3:0] _T_9421; // @[Bitwise.scala 48:55:@9474.4]
  wire [4:0] _T_9422; // @[Bitwise.scala 48:55:@9475.4]
  wire [5:0] _T_9423; // @[Bitwise.scala 48:55:@9476.4]
  wire [6:0] _T_9424; // @[Bitwise.scala 48:55:@9477.4]
  wire [59:0] _T_9488; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@9542.4]
  wire  _T_9489; // @[Bitwise.scala 50:65:@9543.4]
  wire  _T_9490; // @[Bitwise.scala 50:65:@9544.4]
  wire  _T_9491; // @[Bitwise.scala 50:65:@9545.4]
  wire  _T_9492; // @[Bitwise.scala 50:65:@9546.4]
  wire  _T_9493; // @[Bitwise.scala 50:65:@9547.4]
  wire  _T_9494; // @[Bitwise.scala 50:65:@9548.4]
  wire  _T_9495; // @[Bitwise.scala 50:65:@9549.4]
  wire  _T_9496; // @[Bitwise.scala 50:65:@9550.4]
  wire  _T_9497; // @[Bitwise.scala 50:65:@9551.4]
  wire  _T_9498; // @[Bitwise.scala 50:65:@9552.4]
  wire  _T_9499; // @[Bitwise.scala 50:65:@9553.4]
  wire  _T_9500; // @[Bitwise.scala 50:65:@9554.4]
  wire  _T_9501; // @[Bitwise.scala 50:65:@9555.4]
  wire  _T_9502; // @[Bitwise.scala 50:65:@9556.4]
  wire  _T_9503; // @[Bitwise.scala 50:65:@9557.4]
  wire  _T_9504; // @[Bitwise.scala 50:65:@9558.4]
  wire  _T_9505; // @[Bitwise.scala 50:65:@9559.4]
  wire  _T_9506; // @[Bitwise.scala 50:65:@9560.4]
  wire  _T_9507; // @[Bitwise.scala 50:65:@9561.4]
  wire  _T_9508; // @[Bitwise.scala 50:65:@9562.4]
  wire  _T_9509; // @[Bitwise.scala 50:65:@9563.4]
  wire  _T_9510; // @[Bitwise.scala 50:65:@9564.4]
  wire  _T_9511; // @[Bitwise.scala 50:65:@9565.4]
  wire  _T_9512; // @[Bitwise.scala 50:65:@9566.4]
  wire  _T_9513; // @[Bitwise.scala 50:65:@9567.4]
  wire  _T_9514; // @[Bitwise.scala 50:65:@9568.4]
  wire  _T_9515; // @[Bitwise.scala 50:65:@9569.4]
  wire  _T_9516; // @[Bitwise.scala 50:65:@9570.4]
  wire  _T_9517; // @[Bitwise.scala 50:65:@9571.4]
  wire  _T_9518; // @[Bitwise.scala 50:65:@9572.4]
  wire  _T_9519; // @[Bitwise.scala 50:65:@9573.4]
  wire  _T_9520; // @[Bitwise.scala 50:65:@9574.4]
  wire  _T_9521; // @[Bitwise.scala 50:65:@9575.4]
  wire  _T_9522; // @[Bitwise.scala 50:65:@9576.4]
  wire  _T_9523; // @[Bitwise.scala 50:65:@9577.4]
  wire  _T_9524; // @[Bitwise.scala 50:65:@9578.4]
  wire  _T_9525; // @[Bitwise.scala 50:65:@9579.4]
  wire  _T_9526; // @[Bitwise.scala 50:65:@9580.4]
  wire  _T_9527; // @[Bitwise.scala 50:65:@9581.4]
  wire  _T_9528; // @[Bitwise.scala 50:65:@9582.4]
  wire  _T_9529; // @[Bitwise.scala 50:65:@9583.4]
  wire  _T_9530; // @[Bitwise.scala 50:65:@9584.4]
  wire  _T_9531; // @[Bitwise.scala 50:65:@9585.4]
  wire  _T_9532; // @[Bitwise.scala 50:65:@9586.4]
  wire  _T_9533; // @[Bitwise.scala 50:65:@9587.4]
  wire  _T_9534; // @[Bitwise.scala 50:65:@9588.4]
  wire  _T_9535; // @[Bitwise.scala 50:65:@9589.4]
  wire  _T_9536; // @[Bitwise.scala 50:65:@9590.4]
  wire  _T_9537; // @[Bitwise.scala 50:65:@9591.4]
  wire  _T_9538; // @[Bitwise.scala 50:65:@9592.4]
  wire  _T_9539; // @[Bitwise.scala 50:65:@9593.4]
  wire  _T_9540; // @[Bitwise.scala 50:65:@9594.4]
  wire  _T_9541; // @[Bitwise.scala 50:65:@9595.4]
  wire  _T_9542; // @[Bitwise.scala 50:65:@9596.4]
  wire  _T_9543; // @[Bitwise.scala 50:65:@9597.4]
  wire  _T_9544; // @[Bitwise.scala 50:65:@9598.4]
  wire  _T_9545; // @[Bitwise.scala 50:65:@9599.4]
  wire  _T_9546; // @[Bitwise.scala 50:65:@9600.4]
  wire  _T_9547; // @[Bitwise.scala 50:65:@9601.4]
  wire  _T_9548; // @[Bitwise.scala 50:65:@9602.4]
  wire [1:0] _T_9549; // @[Bitwise.scala 48:55:@9603.4]
  wire [1:0] _GEN_987; // @[Bitwise.scala 48:55:@9604.4]
  wire [2:0] _T_9550; // @[Bitwise.scala 48:55:@9604.4]
  wire [1:0] _T_9551; // @[Bitwise.scala 48:55:@9605.4]
  wire [1:0] _T_9552; // @[Bitwise.scala 48:55:@9606.4]
  wire [2:0] _T_9553; // @[Bitwise.scala 48:55:@9607.4]
  wire [3:0] _T_9554; // @[Bitwise.scala 48:55:@9608.4]
  wire [1:0] _T_9555; // @[Bitwise.scala 48:55:@9609.4]
  wire [1:0] _T_9556; // @[Bitwise.scala 48:55:@9610.4]
  wire [2:0] _T_9557; // @[Bitwise.scala 48:55:@9611.4]
  wire [1:0] _T_9558; // @[Bitwise.scala 48:55:@9612.4]
  wire [1:0] _T_9559; // @[Bitwise.scala 48:55:@9613.4]
  wire [2:0] _T_9560; // @[Bitwise.scala 48:55:@9614.4]
  wire [3:0] _T_9561; // @[Bitwise.scala 48:55:@9615.4]
  wire [4:0] _T_9562; // @[Bitwise.scala 48:55:@9616.4]
  wire [1:0] _T_9563; // @[Bitwise.scala 48:55:@9617.4]
  wire [1:0] _GEN_988; // @[Bitwise.scala 48:55:@9618.4]
  wire [2:0] _T_9564; // @[Bitwise.scala 48:55:@9618.4]
  wire [1:0] _T_9565; // @[Bitwise.scala 48:55:@9619.4]
  wire [1:0] _T_9566; // @[Bitwise.scala 48:55:@9620.4]
  wire [2:0] _T_9567; // @[Bitwise.scala 48:55:@9621.4]
  wire [3:0] _T_9568; // @[Bitwise.scala 48:55:@9622.4]
  wire [1:0] _T_9569; // @[Bitwise.scala 48:55:@9623.4]
  wire [1:0] _T_9570; // @[Bitwise.scala 48:55:@9624.4]
  wire [2:0] _T_9571; // @[Bitwise.scala 48:55:@9625.4]
  wire [1:0] _T_9572; // @[Bitwise.scala 48:55:@9626.4]
  wire [1:0] _T_9573; // @[Bitwise.scala 48:55:@9627.4]
  wire [2:0] _T_9574; // @[Bitwise.scala 48:55:@9628.4]
  wire [3:0] _T_9575; // @[Bitwise.scala 48:55:@9629.4]
  wire [4:0] _T_9576; // @[Bitwise.scala 48:55:@9630.4]
  wire [5:0] _T_9577; // @[Bitwise.scala 48:55:@9631.4]
  wire [1:0] _T_9578; // @[Bitwise.scala 48:55:@9632.4]
  wire [1:0] _GEN_989; // @[Bitwise.scala 48:55:@9633.4]
  wire [2:0] _T_9579; // @[Bitwise.scala 48:55:@9633.4]
  wire [1:0] _T_9580; // @[Bitwise.scala 48:55:@9634.4]
  wire [1:0] _T_9581; // @[Bitwise.scala 48:55:@9635.4]
  wire [2:0] _T_9582; // @[Bitwise.scala 48:55:@9636.4]
  wire [3:0] _T_9583; // @[Bitwise.scala 48:55:@9637.4]
  wire [1:0] _T_9584; // @[Bitwise.scala 48:55:@9638.4]
  wire [1:0] _T_9585; // @[Bitwise.scala 48:55:@9639.4]
  wire [2:0] _T_9586; // @[Bitwise.scala 48:55:@9640.4]
  wire [1:0] _T_9587; // @[Bitwise.scala 48:55:@9641.4]
  wire [1:0] _T_9588; // @[Bitwise.scala 48:55:@9642.4]
  wire [2:0] _T_9589; // @[Bitwise.scala 48:55:@9643.4]
  wire [3:0] _T_9590; // @[Bitwise.scala 48:55:@9644.4]
  wire [4:0] _T_9591; // @[Bitwise.scala 48:55:@9645.4]
  wire [1:0] _T_9592; // @[Bitwise.scala 48:55:@9646.4]
  wire [1:0] _GEN_990; // @[Bitwise.scala 48:55:@9647.4]
  wire [2:0] _T_9593; // @[Bitwise.scala 48:55:@9647.4]
  wire [1:0] _T_9594; // @[Bitwise.scala 48:55:@9648.4]
  wire [1:0] _T_9595; // @[Bitwise.scala 48:55:@9649.4]
  wire [2:0] _T_9596; // @[Bitwise.scala 48:55:@9650.4]
  wire [3:0] _T_9597; // @[Bitwise.scala 48:55:@9651.4]
  wire [1:0] _T_9598; // @[Bitwise.scala 48:55:@9652.4]
  wire [1:0] _T_9599; // @[Bitwise.scala 48:55:@9653.4]
  wire [2:0] _T_9600; // @[Bitwise.scala 48:55:@9654.4]
  wire [1:0] _T_9601; // @[Bitwise.scala 48:55:@9655.4]
  wire [1:0] _T_9602; // @[Bitwise.scala 48:55:@9656.4]
  wire [2:0] _T_9603; // @[Bitwise.scala 48:55:@9657.4]
  wire [3:0] _T_9604; // @[Bitwise.scala 48:55:@9658.4]
  wire [4:0] _T_9605; // @[Bitwise.scala 48:55:@9659.4]
  wire [5:0] _T_9606; // @[Bitwise.scala 48:55:@9660.4]
  wire [6:0] _T_9607; // @[Bitwise.scala 48:55:@9661.4]
  wire [60:0] _T_9671; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@9726.4]
  wire  _T_9672; // @[Bitwise.scala 50:65:@9727.4]
  wire  _T_9673; // @[Bitwise.scala 50:65:@9728.4]
  wire  _T_9674; // @[Bitwise.scala 50:65:@9729.4]
  wire  _T_9675; // @[Bitwise.scala 50:65:@9730.4]
  wire  _T_9676; // @[Bitwise.scala 50:65:@9731.4]
  wire  _T_9677; // @[Bitwise.scala 50:65:@9732.4]
  wire  _T_9678; // @[Bitwise.scala 50:65:@9733.4]
  wire  _T_9679; // @[Bitwise.scala 50:65:@9734.4]
  wire  _T_9680; // @[Bitwise.scala 50:65:@9735.4]
  wire  _T_9681; // @[Bitwise.scala 50:65:@9736.4]
  wire  _T_9682; // @[Bitwise.scala 50:65:@9737.4]
  wire  _T_9683; // @[Bitwise.scala 50:65:@9738.4]
  wire  _T_9684; // @[Bitwise.scala 50:65:@9739.4]
  wire  _T_9685; // @[Bitwise.scala 50:65:@9740.4]
  wire  _T_9686; // @[Bitwise.scala 50:65:@9741.4]
  wire  _T_9687; // @[Bitwise.scala 50:65:@9742.4]
  wire  _T_9688; // @[Bitwise.scala 50:65:@9743.4]
  wire  _T_9689; // @[Bitwise.scala 50:65:@9744.4]
  wire  _T_9690; // @[Bitwise.scala 50:65:@9745.4]
  wire  _T_9691; // @[Bitwise.scala 50:65:@9746.4]
  wire  _T_9692; // @[Bitwise.scala 50:65:@9747.4]
  wire  _T_9693; // @[Bitwise.scala 50:65:@9748.4]
  wire  _T_9694; // @[Bitwise.scala 50:65:@9749.4]
  wire  _T_9695; // @[Bitwise.scala 50:65:@9750.4]
  wire  _T_9696; // @[Bitwise.scala 50:65:@9751.4]
  wire  _T_9697; // @[Bitwise.scala 50:65:@9752.4]
  wire  _T_9698; // @[Bitwise.scala 50:65:@9753.4]
  wire  _T_9699; // @[Bitwise.scala 50:65:@9754.4]
  wire  _T_9700; // @[Bitwise.scala 50:65:@9755.4]
  wire  _T_9701; // @[Bitwise.scala 50:65:@9756.4]
  wire  _T_9702; // @[Bitwise.scala 50:65:@9757.4]
  wire  _T_9703; // @[Bitwise.scala 50:65:@9758.4]
  wire  _T_9704; // @[Bitwise.scala 50:65:@9759.4]
  wire  _T_9705; // @[Bitwise.scala 50:65:@9760.4]
  wire  _T_9706; // @[Bitwise.scala 50:65:@9761.4]
  wire  _T_9707; // @[Bitwise.scala 50:65:@9762.4]
  wire  _T_9708; // @[Bitwise.scala 50:65:@9763.4]
  wire  _T_9709; // @[Bitwise.scala 50:65:@9764.4]
  wire  _T_9710; // @[Bitwise.scala 50:65:@9765.4]
  wire  _T_9711; // @[Bitwise.scala 50:65:@9766.4]
  wire  _T_9712; // @[Bitwise.scala 50:65:@9767.4]
  wire  _T_9713; // @[Bitwise.scala 50:65:@9768.4]
  wire  _T_9714; // @[Bitwise.scala 50:65:@9769.4]
  wire  _T_9715; // @[Bitwise.scala 50:65:@9770.4]
  wire  _T_9716; // @[Bitwise.scala 50:65:@9771.4]
  wire  _T_9717; // @[Bitwise.scala 50:65:@9772.4]
  wire  _T_9718; // @[Bitwise.scala 50:65:@9773.4]
  wire  _T_9719; // @[Bitwise.scala 50:65:@9774.4]
  wire  _T_9720; // @[Bitwise.scala 50:65:@9775.4]
  wire  _T_9721; // @[Bitwise.scala 50:65:@9776.4]
  wire  _T_9722; // @[Bitwise.scala 50:65:@9777.4]
  wire  _T_9723; // @[Bitwise.scala 50:65:@9778.4]
  wire  _T_9724; // @[Bitwise.scala 50:65:@9779.4]
  wire  _T_9725; // @[Bitwise.scala 50:65:@9780.4]
  wire  _T_9726; // @[Bitwise.scala 50:65:@9781.4]
  wire  _T_9727; // @[Bitwise.scala 50:65:@9782.4]
  wire  _T_9728; // @[Bitwise.scala 50:65:@9783.4]
  wire  _T_9729; // @[Bitwise.scala 50:65:@9784.4]
  wire  _T_9730; // @[Bitwise.scala 50:65:@9785.4]
  wire  _T_9731; // @[Bitwise.scala 50:65:@9786.4]
  wire  _T_9732; // @[Bitwise.scala 50:65:@9787.4]
  wire [1:0] _T_9733; // @[Bitwise.scala 48:55:@9788.4]
  wire [1:0] _GEN_991; // @[Bitwise.scala 48:55:@9789.4]
  wire [2:0] _T_9734; // @[Bitwise.scala 48:55:@9789.4]
  wire [1:0] _T_9735; // @[Bitwise.scala 48:55:@9790.4]
  wire [1:0] _T_9736; // @[Bitwise.scala 48:55:@9791.4]
  wire [2:0] _T_9737; // @[Bitwise.scala 48:55:@9792.4]
  wire [3:0] _T_9738; // @[Bitwise.scala 48:55:@9793.4]
  wire [1:0] _T_9739; // @[Bitwise.scala 48:55:@9794.4]
  wire [1:0] _T_9740; // @[Bitwise.scala 48:55:@9795.4]
  wire [2:0] _T_9741; // @[Bitwise.scala 48:55:@9796.4]
  wire [1:0] _T_9742; // @[Bitwise.scala 48:55:@9797.4]
  wire [1:0] _T_9743; // @[Bitwise.scala 48:55:@9798.4]
  wire [2:0] _T_9744; // @[Bitwise.scala 48:55:@9799.4]
  wire [3:0] _T_9745; // @[Bitwise.scala 48:55:@9800.4]
  wire [4:0] _T_9746; // @[Bitwise.scala 48:55:@9801.4]
  wire [1:0] _T_9747; // @[Bitwise.scala 48:55:@9802.4]
  wire [1:0] _GEN_992; // @[Bitwise.scala 48:55:@9803.4]
  wire [2:0] _T_9748; // @[Bitwise.scala 48:55:@9803.4]
  wire [1:0] _T_9749; // @[Bitwise.scala 48:55:@9804.4]
  wire [1:0] _T_9750; // @[Bitwise.scala 48:55:@9805.4]
  wire [2:0] _T_9751; // @[Bitwise.scala 48:55:@9806.4]
  wire [3:0] _T_9752; // @[Bitwise.scala 48:55:@9807.4]
  wire [1:0] _T_9753; // @[Bitwise.scala 48:55:@9808.4]
  wire [1:0] _T_9754; // @[Bitwise.scala 48:55:@9809.4]
  wire [2:0] _T_9755; // @[Bitwise.scala 48:55:@9810.4]
  wire [1:0] _T_9756; // @[Bitwise.scala 48:55:@9811.4]
  wire [1:0] _T_9757; // @[Bitwise.scala 48:55:@9812.4]
  wire [2:0] _T_9758; // @[Bitwise.scala 48:55:@9813.4]
  wire [3:0] _T_9759; // @[Bitwise.scala 48:55:@9814.4]
  wire [4:0] _T_9760; // @[Bitwise.scala 48:55:@9815.4]
  wire [5:0] _T_9761; // @[Bitwise.scala 48:55:@9816.4]
  wire [1:0] _T_9762; // @[Bitwise.scala 48:55:@9817.4]
  wire [1:0] _GEN_993; // @[Bitwise.scala 48:55:@9818.4]
  wire [2:0] _T_9763; // @[Bitwise.scala 48:55:@9818.4]
  wire [1:0] _T_9764; // @[Bitwise.scala 48:55:@9819.4]
  wire [1:0] _T_9765; // @[Bitwise.scala 48:55:@9820.4]
  wire [2:0] _T_9766; // @[Bitwise.scala 48:55:@9821.4]
  wire [3:0] _T_9767; // @[Bitwise.scala 48:55:@9822.4]
  wire [1:0] _T_9768; // @[Bitwise.scala 48:55:@9823.4]
  wire [1:0] _T_9769; // @[Bitwise.scala 48:55:@9824.4]
  wire [2:0] _T_9770; // @[Bitwise.scala 48:55:@9825.4]
  wire [1:0] _T_9771; // @[Bitwise.scala 48:55:@9826.4]
  wire [1:0] _T_9772; // @[Bitwise.scala 48:55:@9827.4]
  wire [2:0] _T_9773; // @[Bitwise.scala 48:55:@9828.4]
  wire [3:0] _T_9774; // @[Bitwise.scala 48:55:@9829.4]
  wire [4:0] _T_9775; // @[Bitwise.scala 48:55:@9830.4]
  wire [1:0] _T_9776; // @[Bitwise.scala 48:55:@9831.4]
  wire [1:0] _T_9777; // @[Bitwise.scala 48:55:@9832.4]
  wire [2:0] _T_9778; // @[Bitwise.scala 48:55:@9833.4]
  wire [1:0] _T_9779; // @[Bitwise.scala 48:55:@9834.4]
  wire [1:0] _T_9780; // @[Bitwise.scala 48:55:@9835.4]
  wire [2:0] _T_9781; // @[Bitwise.scala 48:55:@9836.4]
  wire [3:0] _T_9782; // @[Bitwise.scala 48:55:@9837.4]
  wire [1:0] _T_9783; // @[Bitwise.scala 48:55:@9838.4]
  wire [1:0] _T_9784; // @[Bitwise.scala 48:55:@9839.4]
  wire [2:0] _T_9785; // @[Bitwise.scala 48:55:@9840.4]
  wire [1:0] _T_9786; // @[Bitwise.scala 48:55:@9841.4]
  wire [1:0] _T_9787; // @[Bitwise.scala 48:55:@9842.4]
  wire [2:0] _T_9788; // @[Bitwise.scala 48:55:@9843.4]
  wire [3:0] _T_9789; // @[Bitwise.scala 48:55:@9844.4]
  wire [4:0] _T_9790; // @[Bitwise.scala 48:55:@9845.4]
  wire [5:0] _T_9791; // @[Bitwise.scala 48:55:@9846.4]
  wire [6:0] _T_9792; // @[Bitwise.scala 48:55:@9847.4]
  wire [61:0] _T_9856; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@9912.4]
  wire  _T_9857; // @[Bitwise.scala 50:65:@9913.4]
  wire  _T_9858; // @[Bitwise.scala 50:65:@9914.4]
  wire  _T_9859; // @[Bitwise.scala 50:65:@9915.4]
  wire  _T_9860; // @[Bitwise.scala 50:65:@9916.4]
  wire  _T_9861; // @[Bitwise.scala 50:65:@9917.4]
  wire  _T_9862; // @[Bitwise.scala 50:65:@9918.4]
  wire  _T_9863; // @[Bitwise.scala 50:65:@9919.4]
  wire  _T_9864; // @[Bitwise.scala 50:65:@9920.4]
  wire  _T_9865; // @[Bitwise.scala 50:65:@9921.4]
  wire  _T_9866; // @[Bitwise.scala 50:65:@9922.4]
  wire  _T_9867; // @[Bitwise.scala 50:65:@9923.4]
  wire  _T_9868; // @[Bitwise.scala 50:65:@9924.4]
  wire  _T_9869; // @[Bitwise.scala 50:65:@9925.4]
  wire  _T_9870; // @[Bitwise.scala 50:65:@9926.4]
  wire  _T_9871; // @[Bitwise.scala 50:65:@9927.4]
  wire  _T_9872; // @[Bitwise.scala 50:65:@9928.4]
  wire  _T_9873; // @[Bitwise.scala 50:65:@9929.4]
  wire  _T_9874; // @[Bitwise.scala 50:65:@9930.4]
  wire  _T_9875; // @[Bitwise.scala 50:65:@9931.4]
  wire  _T_9876; // @[Bitwise.scala 50:65:@9932.4]
  wire  _T_9877; // @[Bitwise.scala 50:65:@9933.4]
  wire  _T_9878; // @[Bitwise.scala 50:65:@9934.4]
  wire  _T_9879; // @[Bitwise.scala 50:65:@9935.4]
  wire  _T_9880; // @[Bitwise.scala 50:65:@9936.4]
  wire  _T_9881; // @[Bitwise.scala 50:65:@9937.4]
  wire  _T_9882; // @[Bitwise.scala 50:65:@9938.4]
  wire  _T_9883; // @[Bitwise.scala 50:65:@9939.4]
  wire  _T_9884; // @[Bitwise.scala 50:65:@9940.4]
  wire  _T_9885; // @[Bitwise.scala 50:65:@9941.4]
  wire  _T_9886; // @[Bitwise.scala 50:65:@9942.4]
  wire  _T_9887; // @[Bitwise.scala 50:65:@9943.4]
  wire  _T_9888; // @[Bitwise.scala 50:65:@9944.4]
  wire  _T_9889; // @[Bitwise.scala 50:65:@9945.4]
  wire  _T_9890; // @[Bitwise.scala 50:65:@9946.4]
  wire  _T_9891; // @[Bitwise.scala 50:65:@9947.4]
  wire  _T_9892; // @[Bitwise.scala 50:65:@9948.4]
  wire  _T_9893; // @[Bitwise.scala 50:65:@9949.4]
  wire  _T_9894; // @[Bitwise.scala 50:65:@9950.4]
  wire  _T_9895; // @[Bitwise.scala 50:65:@9951.4]
  wire  _T_9896; // @[Bitwise.scala 50:65:@9952.4]
  wire  _T_9897; // @[Bitwise.scala 50:65:@9953.4]
  wire  _T_9898; // @[Bitwise.scala 50:65:@9954.4]
  wire  _T_9899; // @[Bitwise.scala 50:65:@9955.4]
  wire  _T_9900; // @[Bitwise.scala 50:65:@9956.4]
  wire  _T_9901; // @[Bitwise.scala 50:65:@9957.4]
  wire  _T_9902; // @[Bitwise.scala 50:65:@9958.4]
  wire  _T_9903; // @[Bitwise.scala 50:65:@9959.4]
  wire  _T_9904; // @[Bitwise.scala 50:65:@9960.4]
  wire  _T_9905; // @[Bitwise.scala 50:65:@9961.4]
  wire  _T_9906; // @[Bitwise.scala 50:65:@9962.4]
  wire  _T_9907; // @[Bitwise.scala 50:65:@9963.4]
  wire  _T_9908; // @[Bitwise.scala 50:65:@9964.4]
  wire  _T_9909; // @[Bitwise.scala 50:65:@9965.4]
  wire  _T_9910; // @[Bitwise.scala 50:65:@9966.4]
  wire  _T_9911; // @[Bitwise.scala 50:65:@9967.4]
  wire  _T_9912; // @[Bitwise.scala 50:65:@9968.4]
  wire  _T_9913; // @[Bitwise.scala 50:65:@9969.4]
  wire  _T_9914; // @[Bitwise.scala 50:65:@9970.4]
  wire  _T_9915; // @[Bitwise.scala 50:65:@9971.4]
  wire  _T_9916; // @[Bitwise.scala 50:65:@9972.4]
  wire  _T_9917; // @[Bitwise.scala 50:65:@9973.4]
  wire  _T_9918; // @[Bitwise.scala 50:65:@9974.4]
  wire [1:0] _T_9919; // @[Bitwise.scala 48:55:@9975.4]
  wire [1:0] _GEN_994; // @[Bitwise.scala 48:55:@9976.4]
  wire [2:0] _T_9920; // @[Bitwise.scala 48:55:@9976.4]
  wire [1:0] _T_9921; // @[Bitwise.scala 48:55:@9977.4]
  wire [1:0] _T_9922; // @[Bitwise.scala 48:55:@9978.4]
  wire [2:0] _T_9923; // @[Bitwise.scala 48:55:@9979.4]
  wire [3:0] _T_9924; // @[Bitwise.scala 48:55:@9980.4]
  wire [1:0] _T_9925; // @[Bitwise.scala 48:55:@9981.4]
  wire [1:0] _T_9926; // @[Bitwise.scala 48:55:@9982.4]
  wire [2:0] _T_9927; // @[Bitwise.scala 48:55:@9983.4]
  wire [1:0] _T_9928; // @[Bitwise.scala 48:55:@9984.4]
  wire [1:0] _T_9929; // @[Bitwise.scala 48:55:@9985.4]
  wire [2:0] _T_9930; // @[Bitwise.scala 48:55:@9986.4]
  wire [3:0] _T_9931; // @[Bitwise.scala 48:55:@9987.4]
  wire [4:0] _T_9932; // @[Bitwise.scala 48:55:@9988.4]
  wire [1:0] _T_9933; // @[Bitwise.scala 48:55:@9989.4]
  wire [1:0] _T_9934; // @[Bitwise.scala 48:55:@9990.4]
  wire [2:0] _T_9935; // @[Bitwise.scala 48:55:@9991.4]
  wire [1:0] _T_9936; // @[Bitwise.scala 48:55:@9992.4]
  wire [1:0] _T_9937; // @[Bitwise.scala 48:55:@9993.4]
  wire [2:0] _T_9938; // @[Bitwise.scala 48:55:@9994.4]
  wire [3:0] _T_9939; // @[Bitwise.scala 48:55:@9995.4]
  wire [1:0] _T_9940; // @[Bitwise.scala 48:55:@9996.4]
  wire [1:0] _T_9941; // @[Bitwise.scala 48:55:@9997.4]
  wire [2:0] _T_9942; // @[Bitwise.scala 48:55:@9998.4]
  wire [1:0] _T_9943; // @[Bitwise.scala 48:55:@9999.4]
  wire [1:0] _T_9944; // @[Bitwise.scala 48:55:@10000.4]
  wire [2:0] _T_9945; // @[Bitwise.scala 48:55:@10001.4]
  wire [3:0] _T_9946; // @[Bitwise.scala 48:55:@10002.4]
  wire [4:0] _T_9947; // @[Bitwise.scala 48:55:@10003.4]
  wire [5:0] _T_9948; // @[Bitwise.scala 48:55:@10004.4]
  wire [1:0] _T_9949; // @[Bitwise.scala 48:55:@10005.4]
  wire [1:0] _GEN_995; // @[Bitwise.scala 48:55:@10006.4]
  wire [2:0] _T_9950; // @[Bitwise.scala 48:55:@10006.4]
  wire [1:0] _T_9951; // @[Bitwise.scala 48:55:@10007.4]
  wire [1:0] _T_9952; // @[Bitwise.scala 48:55:@10008.4]
  wire [2:0] _T_9953; // @[Bitwise.scala 48:55:@10009.4]
  wire [3:0] _T_9954; // @[Bitwise.scala 48:55:@10010.4]
  wire [1:0] _T_9955; // @[Bitwise.scala 48:55:@10011.4]
  wire [1:0] _T_9956; // @[Bitwise.scala 48:55:@10012.4]
  wire [2:0] _T_9957; // @[Bitwise.scala 48:55:@10013.4]
  wire [1:0] _T_9958; // @[Bitwise.scala 48:55:@10014.4]
  wire [1:0] _T_9959; // @[Bitwise.scala 48:55:@10015.4]
  wire [2:0] _T_9960; // @[Bitwise.scala 48:55:@10016.4]
  wire [3:0] _T_9961; // @[Bitwise.scala 48:55:@10017.4]
  wire [4:0] _T_9962; // @[Bitwise.scala 48:55:@10018.4]
  wire [1:0] _T_9963; // @[Bitwise.scala 48:55:@10019.4]
  wire [1:0] _T_9964; // @[Bitwise.scala 48:55:@10020.4]
  wire [2:0] _T_9965; // @[Bitwise.scala 48:55:@10021.4]
  wire [1:0] _T_9966; // @[Bitwise.scala 48:55:@10022.4]
  wire [1:0] _T_9967; // @[Bitwise.scala 48:55:@10023.4]
  wire [2:0] _T_9968; // @[Bitwise.scala 48:55:@10024.4]
  wire [3:0] _T_9969; // @[Bitwise.scala 48:55:@10025.4]
  wire [1:0] _T_9970; // @[Bitwise.scala 48:55:@10026.4]
  wire [1:0] _T_9971; // @[Bitwise.scala 48:55:@10027.4]
  wire [2:0] _T_9972; // @[Bitwise.scala 48:55:@10028.4]
  wire [1:0] _T_9973; // @[Bitwise.scala 48:55:@10029.4]
  wire [1:0] _T_9974; // @[Bitwise.scala 48:55:@10030.4]
  wire [2:0] _T_9975; // @[Bitwise.scala 48:55:@10031.4]
  wire [3:0] _T_9976; // @[Bitwise.scala 48:55:@10032.4]
  wire [4:0] _T_9977; // @[Bitwise.scala 48:55:@10033.4]
  wire [5:0] _T_9978; // @[Bitwise.scala 48:55:@10034.4]
  wire [6:0] _T_9979; // @[Bitwise.scala 48:55:@10035.4]
  wire [62:0] _T_10043; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@10100.4]
  wire  _T_10044; // @[Bitwise.scala 50:65:@10101.4]
  wire  _T_10045; // @[Bitwise.scala 50:65:@10102.4]
  wire  _T_10046; // @[Bitwise.scala 50:65:@10103.4]
  wire  _T_10047; // @[Bitwise.scala 50:65:@10104.4]
  wire  _T_10048; // @[Bitwise.scala 50:65:@10105.4]
  wire  _T_10049; // @[Bitwise.scala 50:65:@10106.4]
  wire  _T_10050; // @[Bitwise.scala 50:65:@10107.4]
  wire  _T_10051; // @[Bitwise.scala 50:65:@10108.4]
  wire  _T_10052; // @[Bitwise.scala 50:65:@10109.4]
  wire  _T_10053; // @[Bitwise.scala 50:65:@10110.4]
  wire  _T_10054; // @[Bitwise.scala 50:65:@10111.4]
  wire  _T_10055; // @[Bitwise.scala 50:65:@10112.4]
  wire  _T_10056; // @[Bitwise.scala 50:65:@10113.4]
  wire  _T_10057; // @[Bitwise.scala 50:65:@10114.4]
  wire  _T_10058; // @[Bitwise.scala 50:65:@10115.4]
  wire  _T_10059; // @[Bitwise.scala 50:65:@10116.4]
  wire  _T_10060; // @[Bitwise.scala 50:65:@10117.4]
  wire  _T_10061; // @[Bitwise.scala 50:65:@10118.4]
  wire  _T_10062; // @[Bitwise.scala 50:65:@10119.4]
  wire  _T_10063; // @[Bitwise.scala 50:65:@10120.4]
  wire  _T_10064; // @[Bitwise.scala 50:65:@10121.4]
  wire  _T_10065; // @[Bitwise.scala 50:65:@10122.4]
  wire  _T_10066; // @[Bitwise.scala 50:65:@10123.4]
  wire  _T_10067; // @[Bitwise.scala 50:65:@10124.4]
  wire  _T_10068; // @[Bitwise.scala 50:65:@10125.4]
  wire  _T_10069; // @[Bitwise.scala 50:65:@10126.4]
  wire  _T_10070; // @[Bitwise.scala 50:65:@10127.4]
  wire  _T_10071; // @[Bitwise.scala 50:65:@10128.4]
  wire  _T_10072; // @[Bitwise.scala 50:65:@10129.4]
  wire  _T_10073; // @[Bitwise.scala 50:65:@10130.4]
  wire  _T_10074; // @[Bitwise.scala 50:65:@10131.4]
  wire  _T_10075; // @[Bitwise.scala 50:65:@10132.4]
  wire  _T_10076; // @[Bitwise.scala 50:65:@10133.4]
  wire  _T_10077; // @[Bitwise.scala 50:65:@10134.4]
  wire  _T_10078; // @[Bitwise.scala 50:65:@10135.4]
  wire  _T_10079; // @[Bitwise.scala 50:65:@10136.4]
  wire  _T_10080; // @[Bitwise.scala 50:65:@10137.4]
  wire  _T_10081; // @[Bitwise.scala 50:65:@10138.4]
  wire  _T_10082; // @[Bitwise.scala 50:65:@10139.4]
  wire  _T_10083; // @[Bitwise.scala 50:65:@10140.4]
  wire  _T_10084; // @[Bitwise.scala 50:65:@10141.4]
  wire  _T_10085; // @[Bitwise.scala 50:65:@10142.4]
  wire  _T_10086; // @[Bitwise.scala 50:65:@10143.4]
  wire  _T_10087; // @[Bitwise.scala 50:65:@10144.4]
  wire  _T_10088; // @[Bitwise.scala 50:65:@10145.4]
  wire  _T_10089; // @[Bitwise.scala 50:65:@10146.4]
  wire  _T_10090; // @[Bitwise.scala 50:65:@10147.4]
  wire  _T_10091; // @[Bitwise.scala 50:65:@10148.4]
  wire  _T_10092; // @[Bitwise.scala 50:65:@10149.4]
  wire  _T_10093; // @[Bitwise.scala 50:65:@10150.4]
  wire  _T_10094; // @[Bitwise.scala 50:65:@10151.4]
  wire  _T_10095; // @[Bitwise.scala 50:65:@10152.4]
  wire  _T_10096; // @[Bitwise.scala 50:65:@10153.4]
  wire  _T_10097; // @[Bitwise.scala 50:65:@10154.4]
  wire  _T_10098; // @[Bitwise.scala 50:65:@10155.4]
  wire  _T_10099; // @[Bitwise.scala 50:65:@10156.4]
  wire  _T_10100; // @[Bitwise.scala 50:65:@10157.4]
  wire  _T_10101; // @[Bitwise.scala 50:65:@10158.4]
  wire  _T_10102; // @[Bitwise.scala 50:65:@10159.4]
  wire  _T_10103; // @[Bitwise.scala 50:65:@10160.4]
  wire  _T_10104; // @[Bitwise.scala 50:65:@10161.4]
  wire  _T_10105; // @[Bitwise.scala 50:65:@10162.4]
  wire  _T_10106; // @[Bitwise.scala 50:65:@10163.4]
  wire [1:0] _T_10107; // @[Bitwise.scala 48:55:@10164.4]
  wire [1:0] _GEN_996; // @[Bitwise.scala 48:55:@10165.4]
  wire [2:0] _T_10108; // @[Bitwise.scala 48:55:@10165.4]
  wire [1:0] _T_10109; // @[Bitwise.scala 48:55:@10166.4]
  wire [1:0] _T_10110; // @[Bitwise.scala 48:55:@10167.4]
  wire [2:0] _T_10111; // @[Bitwise.scala 48:55:@10168.4]
  wire [3:0] _T_10112; // @[Bitwise.scala 48:55:@10169.4]
  wire [1:0] _T_10113; // @[Bitwise.scala 48:55:@10170.4]
  wire [1:0] _T_10114; // @[Bitwise.scala 48:55:@10171.4]
  wire [2:0] _T_10115; // @[Bitwise.scala 48:55:@10172.4]
  wire [1:0] _T_10116; // @[Bitwise.scala 48:55:@10173.4]
  wire [1:0] _T_10117; // @[Bitwise.scala 48:55:@10174.4]
  wire [2:0] _T_10118; // @[Bitwise.scala 48:55:@10175.4]
  wire [3:0] _T_10119; // @[Bitwise.scala 48:55:@10176.4]
  wire [4:0] _T_10120; // @[Bitwise.scala 48:55:@10177.4]
  wire [1:0] _T_10121; // @[Bitwise.scala 48:55:@10178.4]
  wire [1:0] _T_10122; // @[Bitwise.scala 48:55:@10179.4]
  wire [2:0] _T_10123; // @[Bitwise.scala 48:55:@10180.4]
  wire [1:0] _T_10124; // @[Bitwise.scala 48:55:@10181.4]
  wire [1:0] _T_10125; // @[Bitwise.scala 48:55:@10182.4]
  wire [2:0] _T_10126; // @[Bitwise.scala 48:55:@10183.4]
  wire [3:0] _T_10127; // @[Bitwise.scala 48:55:@10184.4]
  wire [1:0] _T_10128; // @[Bitwise.scala 48:55:@10185.4]
  wire [1:0] _T_10129; // @[Bitwise.scala 48:55:@10186.4]
  wire [2:0] _T_10130; // @[Bitwise.scala 48:55:@10187.4]
  wire [1:0] _T_10131; // @[Bitwise.scala 48:55:@10188.4]
  wire [1:0] _T_10132; // @[Bitwise.scala 48:55:@10189.4]
  wire [2:0] _T_10133; // @[Bitwise.scala 48:55:@10190.4]
  wire [3:0] _T_10134; // @[Bitwise.scala 48:55:@10191.4]
  wire [4:0] _T_10135; // @[Bitwise.scala 48:55:@10192.4]
  wire [5:0] _T_10136; // @[Bitwise.scala 48:55:@10193.4]
  wire [1:0] _T_10137; // @[Bitwise.scala 48:55:@10194.4]
  wire [1:0] _T_10138; // @[Bitwise.scala 48:55:@10195.4]
  wire [2:0] _T_10139; // @[Bitwise.scala 48:55:@10196.4]
  wire [1:0] _T_10140; // @[Bitwise.scala 48:55:@10197.4]
  wire [1:0] _T_10141; // @[Bitwise.scala 48:55:@10198.4]
  wire [2:0] _T_10142; // @[Bitwise.scala 48:55:@10199.4]
  wire [3:0] _T_10143; // @[Bitwise.scala 48:55:@10200.4]
  wire [1:0] _T_10144; // @[Bitwise.scala 48:55:@10201.4]
  wire [1:0] _T_10145; // @[Bitwise.scala 48:55:@10202.4]
  wire [2:0] _T_10146; // @[Bitwise.scala 48:55:@10203.4]
  wire [1:0] _T_10147; // @[Bitwise.scala 48:55:@10204.4]
  wire [1:0] _T_10148; // @[Bitwise.scala 48:55:@10205.4]
  wire [2:0] _T_10149; // @[Bitwise.scala 48:55:@10206.4]
  wire [3:0] _T_10150; // @[Bitwise.scala 48:55:@10207.4]
  wire [4:0] _T_10151; // @[Bitwise.scala 48:55:@10208.4]
  wire [1:0] _T_10152; // @[Bitwise.scala 48:55:@10209.4]
  wire [1:0] _T_10153; // @[Bitwise.scala 48:55:@10210.4]
  wire [2:0] _T_10154; // @[Bitwise.scala 48:55:@10211.4]
  wire [1:0] _T_10155; // @[Bitwise.scala 48:55:@10212.4]
  wire [1:0] _T_10156; // @[Bitwise.scala 48:55:@10213.4]
  wire [2:0] _T_10157; // @[Bitwise.scala 48:55:@10214.4]
  wire [3:0] _T_10158; // @[Bitwise.scala 48:55:@10215.4]
  wire [1:0] _T_10159; // @[Bitwise.scala 48:55:@10216.4]
  wire [1:0] _T_10160; // @[Bitwise.scala 48:55:@10217.4]
  wire [2:0] _T_10161; // @[Bitwise.scala 48:55:@10218.4]
  wire [1:0] _T_10162; // @[Bitwise.scala 48:55:@10219.4]
  wire [1:0] _T_10163; // @[Bitwise.scala 48:55:@10220.4]
  wire [2:0] _T_10164; // @[Bitwise.scala 48:55:@10221.4]
  wire [3:0] _T_10165; // @[Bitwise.scala 48:55:@10222.4]
  wire [4:0] _T_10166; // @[Bitwise.scala 48:55:@10223.4]
  wire [5:0] _T_10167; // @[Bitwise.scala 48:55:@10224.4]
  wire [6:0] _T_10168; // @[Bitwise.scala 48:55:@10225.4]
  wire  _T_10234; // @[Bitwise.scala 50:65:@10292.4]
  wire  _T_10235; // @[Bitwise.scala 50:65:@10293.4]
  wire  _T_10236; // @[Bitwise.scala 50:65:@10294.4]
  wire  _T_10237; // @[Bitwise.scala 50:65:@10295.4]
  wire  _T_10238; // @[Bitwise.scala 50:65:@10296.4]
  wire  _T_10239; // @[Bitwise.scala 50:65:@10297.4]
  wire  _T_10240; // @[Bitwise.scala 50:65:@10298.4]
  wire  _T_10241; // @[Bitwise.scala 50:65:@10299.4]
  wire  _T_10242; // @[Bitwise.scala 50:65:@10300.4]
  wire  _T_10243; // @[Bitwise.scala 50:65:@10301.4]
  wire  _T_10244; // @[Bitwise.scala 50:65:@10302.4]
  wire  _T_10245; // @[Bitwise.scala 50:65:@10303.4]
  wire  _T_10246; // @[Bitwise.scala 50:65:@10304.4]
  wire  _T_10247; // @[Bitwise.scala 50:65:@10305.4]
  wire  _T_10248; // @[Bitwise.scala 50:65:@10306.4]
  wire  _T_10249; // @[Bitwise.scala 50:65:@10307.4]
  wire  _T_10250; // @[Bitwise.scala 50:65:@10308.4]
  wire  _T_10251; // @[Bitwise.scala 50:65:@10309.4]
  wire  _T_10252; // @[Bitwise.scala 50:65:@10310.4]
  wire  _T_10253; // @[Bitwise.scala 50:65:@10311.4]
  wire  _T_10254; // @[Bitwise.scala 50:65:@10312.4]
  wire  _T_10255; // @[Bitwise.scala 50:65:@10313.4]
  wire  _T_10256; // @[Bitwise.scala 50:65:@10314.4]
  wire  _T_10257; // @[Bitwise.scala 50:65:@10315.4]
  wire  _T_10258; // @[Bitwise.scala 50:65:@10316.4]
  wire  _T_10259; // @[Bitwise.scala 50:65:@10317.4]
  wire  _T_10260; // @[Bitwise.scala 50:65:@10318.4]
  wire  _T_10261; // @[Bitwise.scala 50:65:@10319.4]
  wire  _T_10262; // @[Bitwise.scala 50:65:@10320.4]
  wire  _T_10263; // @[Bitwise.scala 50:65:@10321.4]
  wire  _T_10264; // @[Bitwise.scala 50:65:@10322.4]
  wire  _T_10265; // @[Bitwise.scala 50:65:@10323.4]
  wire  _T_10266; // @[Bitwise.scala 50:65:@10324.4]
  wire  _T_10267; // @[Bitwise.scala 50:65:@10325.4]
  wire  _T_10268; // @[Bitwise.scala 50:65:@10326.4]
  wire  _T_10269; // @[Bitwise.scala 50:65:@10327.4]
  wire  _T_10270; // @[Bitwise.scala 50:65:@10328.4]
  wire  _T_10271; // @[Bitwise.scala 50:65:@10329.4]
  wire  _T_10272; // @[Bitwise.scala 50:65:@10330.4]
  wire  _T_10273; // @[Bitwise.scala 50:65:@10331.4]
  wire  _T_10274; // @[Bitwise.scala 50:65:@10332.4]
  wire  _T_10275; // @[Bitwise.scala 50:65:@10333.4]
  wire  _T_10276; // @[Bitwise.scala 50:65:@10334.4]
  wire  _T_10277; // @[Bitwise.scala 50:65:@10335.4]
  wire  _T_10278; // @[Bitwise.scala 50:65:@10336.4]
  wire  _T_10279; // @[Bitwise.scala 50:65:@10337.4]
  wire  _T_10280; // @[Bitwise.scala 50:65:@10338.4]
  wire  _T_10281; // @[Bitwise.scala 50:65:@10339.4]
  wire  _T_10282; // @[Bitwise.scala 50:65:@10340.4]
  wire  _T_10283; // @[Bitwise.scala 50:65:@10341.4]
  wire  _T_10284; // @[Bitwise.scala 50:65:@10342.4]
  wire  _T_10285; // @[Bitwise.scala 50:65:@10343.4]
  wire  _T_10286; // @[Bitwise.scala 50:65:@10344.4]
  wire  _T_10287; // @[Bitwise.scala 50:65:@10345.4]
  wire  _T_10288; // @[Bitwise.scala 50:65:@10346.4]
  wire  _T_10289; // @[Bitwise.scala 50:65:@10347.4]
  wire  _T_10290; // @[Bitwise.scala 50:65:@10348.4]
  wire  _T_10291; // @[Bitwise.scala 50:65:@10349.4]
  wire  _T_10292; // @[Bitwise.scala 50:65:@10350.4]
  wire  _T_10293; // @[Bitwise.scala 50:65:@10351.4]
  wire  _T_10294; // @[Bitwise.scala 50:65:@10352.4]
  wire  _T_10295; // @[Bitwise.scala 50:65:@10353.4]
  wire  _T_10296; // @[Bitwise.scala 50:65:@10354.4]
  wire [1:0] _T_10297; // @[Bitwise.scala 48:55:@10355.4]
  wire [1:0] _T_10298; // @[Bitwise.scala 48:55:@10356.4]
  wire [2:0] _T_10299; // @[Bitwise.scala 48:55:@10357.4]
  wire [1:0] _T_10300; // @[Bitwise.scala 48:55:@10358.4]
  wire [1:0] _T_10301; // @[Bitwise.scala 48:55:@10359.4]
  wire [2:0] _T_10302; // @[Bitwise.scala 48:55:@10360.4]
  wire [3:0] _T_10303; // @[Bitwise.scala 48:55:@10361.4]
  wire [1:0] _T_10304; // @[Bitwise.scala 48:55:@10362.4]
  wire [1:0] _T_10305; // @[Bitwise.scala 48:55:@10363.4]
  wire [2:0] _T_10306; // @[Bitwise.scala 48:55:@10364.4]
  wire [1:0] _T_10307; // @[Bitwise.scala 48:55:@10365.4]
  wire [1:0] _T_10308; // @[Bitwise.scala 48:55:@10366.4]
  wire [2:0] _T_10309; // @[Bitwise.scala 48:55:@10367.4]
  wire [3:0] _T_10310; // @[Bitwise.scala 48:55:@10368.4]
  wire [4:0] _T_10311; // @[Bitwise.scala 48:55:@10369.4]
  wire [1:0] _T_10312; // @[Bitwise.scala 48:55:@10370.4]
  wire [1:0] _T_10313; // @[Bitwise.scala 48:55:@10371.4]
  wire [2:0] _T_10314; // @[Bitwise.scala 48:55:@10372.4]
  wire [1:0] _T_10315; // @[Bitwise.scala 48:55:@10373.4]
  wire [1:0] _T_10316; // @[Bitwise.scala 48:55:@10374.4]
  wire [2:0] _T_10317; // @[Bitwise.scala 48:55:@10375.4]
  wire [3:0] _T_10318; // @[Bitwise.scala 48:55:@10376.4]
  wire [1:0] _T_10319; // @[Bitwise.scala 48:55:@10377.4]
  wire [1:0] _T_10320; // @[Bitwise.scala 48:55:@10378.4]
  wire [2:0] _T_10321; // @[Bitwise.scala 48:55:@10379.4]
  wire [1:0] _T_10322; // @[Bitwise.scala 48:55:@10380.4]
  wire [1:0] _T_10323; // @[Bitwise.scala 48:55:@10381.4]
  wire [2:0] _T_10324; // @[Bitwise.scala 48:55:@10382.4]
  wire [3:0] _T_10325; // @[Bitwise.scala 48:55:@10383.4]
  wire [4:0] _T_10326; // @[Bitwise.scala 48:55:@10384.4]
  wire [5:0] _T_10327; // @[Bitwise.scala 48:55:@10385.4]
  wire [1:0] _T_10328; // @[Bitwise.scala 48:55:@10386.4]
  wire [1:0] _T_10329; // @[Bitwise.scala 48:55:@10387.4]
  wire [2:0] _T_10330; // @[Bitwise.scala 48:55:@10388.4]
  wire [1:0] _T_10331; // @[Bitwise.scala 48:55:@10389.4]
  wire [1:0] _T_10332; // @[Bitwise.scala 48:55:@10390.4]
  wire [2:0] _T_10333; // @[Bitwise.scala 48:55:@10391.4]
  wire [3:0] _T_10334; // @[Bitwise.scala 48:55:@10392.4]
  wire [1:0] _T_10335; // @[Bitwise.scala 48:55:@10393.4]
  wire [1:0] _T_10336; // @[Bitwise.scala 48:55:@10394.4]
  wire [2:0] _T_10337; // @[Bitwise.scala 48:55:@10395.4]
  wire [1:0] _T_10338; // @[Bitwise.scala 48:55:@10396.4]
  wire [1:0] _T_10339; // @[Bitwise.scala 48:55:@10397.4]
  wire [2:0] _T_10340; // @[Bitwise.scala 48:55:@10398.4]
  wire [3:0] _T_10341; // @[Bitwise.scala 48:55:@10399.4]
  wire [4:0] _T_10342; // @[Bitwise.scala 48:55:@10400.4]
  wire [1:0] _T_10343; // @[Bitwise.scala 48:55:@10401.4]
  wire [1:0] _T_10344; // @[Bitwise.scala 48:55:@10402.4]
  wire [2:0] _T_10345; // @[Bitwise.scala 48:55:@10403.4]
  wire [1:0] _T_10346; // @[Bitwise.scala 48:55:@10404.4]
  wire [1:0] _T_10347; // @[Bitwise.scala 48:55:@10405.4]
  wire [2:0] _T_10348; // @[Bitwise.scala 48:55:@10406.4]
  wire [3:0] _T_10349; // @[Bitwise.scala 48:55:@10407.4]
  wire [1:0] _T_10350; // @[Bitwise.scala 48:55:@10408.4]
  wire [1:0] _T_10351; // @[Bitwise.scala 48:55:@10409.4]
  wire [2:0] _T_10352; // @[Bitwise.scala 48:55:@10410.4]
  wire [1:0] _T_10353; // @[Bitwise.scala 48:55:@10411.4]
  wire [1:0] _T_10354; // @[Bitwise.scala 48:55:@10412.4]
  wire [2:0] _T_10355; // @[Bitwise.scala 48:55:@10413.4]
  wire [3:0] _T_10356; // @[Bitwise.scala 48:55:@10414.4]
  wire [4:0] _T_10357; // @[Bitwise.scala 48:55:@10415.4]
  wire [5:0] _T_10358; // @[Bitwise.scala 48:55:@10416.4]
  wire [6:0] _T_10359; // @[Bitwise.scala 48:55:@10417.4]
  reg  _T_10362; // @[NV_NVDLA_CSC_WL_dec.scala 64:27:@10419.4]
  reg [31:0] _RAND_0;
  reg [7:0] _T_10366_0; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_1;
  reg [7:0] _T_10366_1; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_2;
  reg [7:0] _T_10366_2; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_3;
  reg [7:0] _T_10366_3; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_4;
  reg [7:0] _T_10366_4; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_5;
  reg [7:0] _T_10366_5; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_6;
  reg [7:0] _T_10366_6; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_7;
  reg [7:0] _T_10366_7; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_8;
  reg [7:0] _T_10366_8; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_9;
  reg [7:0] _T_10366_9; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_10;
  reg [7:0] _T_10366_10; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_11;
  reg [7:0] _T_10366_11; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_12;
  reg [7:0] _T_10366_12; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_13;
  reg [7:0] _T_10366_13; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_14;
  reg [7:0] _T_10366_14; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_15;
  reg [7:0] _T_10366_15; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_16;
  reg [7:0] _T_10366_16; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_17;
  reg [7:0] _T_10366_17; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_18;
  reg [7:0] _T_10366_18; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_19;
  reg [7:0] _T_10366_19; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_20;
  reg [7:0] _T_10366_20; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_21;
  reg [7:0] _T_10366_21; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_22;
  reg [7:0] _T_10366_22; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_23;
  reg [7:0] _T_10366_23; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_24;
  reg [7:0] _T_10366_24; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_25;
  reg [7:0] _T_10366_25; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_26;
  reg [7:0] _T_10366_26; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_27;
  reg [7:0] _T_10366_27; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_28;
  reg [7:0] _T_10366_28; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_29;
  reg [7:0] _T_10366_29; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_30;
  reg [7:0] _T_10366_30; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_31;
  reg [7:0] _T_10366_31; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_32;
  reg [7:0] _T_10366_32; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_33;
  reg [7:0] _T_10366_33; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_34;
  reg [7:0] _T_10366_34; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_35;
  reg [7:0] _T_10366_35; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_36;
  reg [7:0] _T_10366_36; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_37;
  reg [7:0] _T_10366_37; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_38;
  reg [7:0] _T_10366_38; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_39;
  reg [7:0] _T_10366_39; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_40;
  reg [7:0] _T_10366_40; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_41;
  reg [7:0] _T_10366_41; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_42;
  reg [7:0] _T_10366_42; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_43;
  reg [7:0] _T_10366_43; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_44;
  reg [7:0] _T_10366_44; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_45;
  reg [7:0] _T_10366_45; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_46;
  reg [7:0] _T_10366_46; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_47;
  reg [7:0] _T_10366_47; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_48;
  reg [7:0] _T_10366_48; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_49;
  reg [7:0] _T_10366_49; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_50;
  reg [7:0] _T_10366_50; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_51;
  reg [7:0] _T_10366_51; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_52;
  reg [7:0] _T_10366_52; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_53;
  reg [7:0] _T_10366_53; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_54;
  reg [7:0] _T_10366_54; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_55;
  reg [7:0] _T_10366_55; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_56;
  reg [7:0] _T_10366_56; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_57;
  reg [7:0] _T_10366_57; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_58;
  reg [7:0] _T_10366_58; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_59;
  reg [7:0] _T_10366_59; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_60;
  reg [7:0] _T_10366_60; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_61;
  reg [7:0] _T_10366_61; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_62;
  reg [7:0] _T_10366_62; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_63;
  reg [7:0] _T_10366_63; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@10420.4]
  reg [31:0] _RAND_64;
  reg  _T_10436_0; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_65;
  reg  _T_10436_1; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_66;
  reg  _T_10436_2; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_67;
  reg  _T_10436_3; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_68;
  reg  _T_10436_4; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_69;
  reg  _T_10436_5; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_70;
  reg  _T_10436_6; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_71;
  reg  _T_10436_7; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_72;
  reg  _T_10436_8; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_73;
  reg  _T_10436_9; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_74;
  reg  _T_10436_10; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_75;
  reg  _T_10436_11; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_76;
  reg  _T_10436_12; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_77;
  reg  _T_10436_13; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_78;
  reg  _T_10436_14; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_79;
  reg  _T_10436_15; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_80;
  reg  _T_10436_16; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_81;
  reg  _T_10436_17; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_82;
  reg  _T_10436_18; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_83;
  reg  _T_10436_19; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_84;
  reg  _T_10436_20; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_85;
  reg  _T_10436_21; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_86;
  reg  _T_10436_22; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_87;
  reg  _T_10436_23; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_88;
  reg  _T_10436_24; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_89;
  reg  _T_10436_25; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_90;
  reg  _T_10436_26; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_91;
  reg  _T_10436_27; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_92;
  reg  _T_10436_28; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_93;
  reg  _T_10436_29; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_94;
  reg  _T_10436_30; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_95;
  reg  _T_10436_31; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_96;
  reg  _T_10436_32; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_97;
  reg  _T_10436_33; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_98;
  reg  _T_10436_34; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_99;
  reg  _T_10436_35; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_100;
  reg  _T_10436_36; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_101;
  reg  _T_10436_37; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_102;
  reg  _T_10436_38; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_103;
  reg  _T_10436_39; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_104;
  reg  _T_10436_40; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_105;
  reg  _T_10436_41; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_106;
  reg  _T_10436_42; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_107;
  reg  _T_10436_43; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_108;
  reg  _T_10436_44; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_109;
  reg  _T_10436_45; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_110;
  reg  _T_10436_46; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_111;
  reg  _T_10436_47; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_112;
  reg  _T_10436_48; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_113;
  reg  _T_10436_49; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_114;
  reg  _T_10436_50; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_115;
  reg  _T_10436_51; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_116;
  reg  _T_10436_52; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_117;
  reg  _T_10436_53; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_118;
  reg  _T_10436_54; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_119;
  reg  _T_10436_55; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_120;
  reg  _T_10436_56; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_121;
  reg  _T_10436_57; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_122;
  reg  _T_10436_58; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_123;
  reg  _T_10436_59; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_124;
  reg  _T_10436_60; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_125;
  reg  _T_10436_61; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_126;
  reg  _T_10436_62; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_127;
  reg  _T_10436_63; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@10421.4]
  reg [31:0] _RAND_128;
  reg  _T_10641_0; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_129;
  reg  _T_10641_1; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_130;
  reg  _T_10641_2; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_131;
  reg  _T_10641_3; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_132;
  reg  _T_10641_4; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_133;
  reg  _T_10641_5; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_134;
  reg  _T_10641_6; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_135;
  reg  _T_10641_7; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_136;
  reg  _T_10641_8; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_137;
  reg  _T_10641_9; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_138;
  reg  _T_10641_10; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_139;
  reg  _T_10641_11; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_140;
  reg  _T_10641_12; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_141;
  reg  _T_10641_13; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_142;
  reg  _T_10641_14; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_143;
  reg  _T_10641_15; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_144;
  reg  _T_10641_16; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_145;
  reg  _T_10641_17; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_146;
  reg  _T_10641_18; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_147;
  reg  _T_10641_19; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_148;
  reg  _T_10641_20; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_149;
  reg  _T_10641_21; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_150;
  reg  _T_10641_22; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_151;
  reg  _T_10641_23; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_152;
  reg  _T_10641_24; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_153;
  reg  _T_10641_25; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_154;
  reg  _T_10641_26; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_155;
  reg  _T_10641_27; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_156;
  reg  _T_10641_28; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_157;
  reg  _T_10641_29; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_158;
  reg  _T_10641_30; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_159;
  reg  _T_10641_31; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@10455.4]
  reg [31:0] _RAND_160;
  reg [6:0] _T_11317_63; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_161;
  reg [5:0] _T_11317_62; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_162;
  reg [5:0] _T_11317_61; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_163;
  reg [5:0] _T_11317_60; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_164;
  reg [5:0] _T_11317_59; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_165;
  reg [5:0] _T_11317_58; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_166;
  reg [5:0] _T_11317_57; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_167;
  reg [5:0] _T_11317_56; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_168;
  reg [5:0] _T_11317_55; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_169;
  reg [5:0] _T_11317_54; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_170;
  reg [5:0] _T_11317_53; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_171;
  reg [5:0] _T_11317_52; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_172;
  reg [5:0] _T_11317_51; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_173;
  reg [5:0] _T_11317_50; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_174;
  reg [5:0] _T_11317_49; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_175;
  reg [5:0] _T_11317_48; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_176;
  reg [5:0] _T_11317_47; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_177;
  reg [5:0] _T_11317_46; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_178;
  reg [5:0] _T_11317_45; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_179;
  reg [5:0] _T_11317_44; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_180;
  reg [5:0] _T_11317_43; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_181;
  reg [5:0] _T_11317_42; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_182;
  reg [5:0] _T_11317_41; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_183;
  reg [5:0] _T_11317_40; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_184;
  reg [5:0] _T_11317_39; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_185;
  reg [5:0] _T_11317_38; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_186;
  reg [5:0] _T_11317_37; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_187;
  reg [5:0] _T_11317_36; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_188;
  reg [5:0] _T_11317_35; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_189;
  reg [5:0] _T_11317_34; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_190;
  reg [5:0] _T_11317_33; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_191;
  reg [5:0] _T_11317_32; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_192;
  reg [5:0] _T_11317_31; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_193;
  reg [4:0] _T_11317_30; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_194;
  reg [4:0] _T_11317_29; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_195;
  reg [4:0] _T_11317_28; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_196;
  reg [4:0] _T_11317_27; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_197;
  reg [4:0] _T_11317_26; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_198;
  reg [4:0] _T_11317_25; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_199;
  reg [4:0] _T_11317_24; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_200;
  reg [4:0] _T_11317_23; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_201;
  reg [4:0] _T_11317_22; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_202;
  reg [4:0] _T_11317_21; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_203;
  reg [4:0] _T_11317_20; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_204;
  reg [4:0] _T_11317_19; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_205;
  reg [4:0] _T_11317_18; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_206;
  reg [4:0] _T_11317_17; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_207;
  reg [4:0] _T_11317_16; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_208;
  reg [4:0] _T_11317_15; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_209;
  reg [3:0] _T_11317_14; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_210;
  reg [3:0] _T_11317_13; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_211;
  reg [3:0] _T_11317_12; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_212;
  reg [3:0] _T_11317_11; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_213;
  reg [3:0] _T_11317_10; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_214;
  reg [3:0] _T_11317_9; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_215;
  reg [3:0] _T_11317_8; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_216;
  reg [3:0] _T_11317_7; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_217;
  reg [2:0] _T_11317_6; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_218;
  reg [2:0] _T_11317_5; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_219;
  reg [2:0] _T_11317_4; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_220;
  reg [2:0] _T_11317_3; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_221;
  reg [1:0] _T_11317_2; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_222;
  reg [1:0] _T_11317_1; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_223;
  reg  _T_11317_0; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@10584.4]
  reg [31:0] _RAND_224;
  wire  _GEN_128; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_129; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_130; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_131; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_132; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_133; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_134; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_135; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_136; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_137; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_138; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_139; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_140; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_141; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_142; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_143; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_144; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_145; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_146; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_147; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_148; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_149; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_150; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_151; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_152; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_153; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_154; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_155; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_156; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_157; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_158; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _GEN_159; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  wire  _T_11318; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@10748.4]
  wire  _T_11319; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@10749.4]
  wire  _GEN_160; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10750.4]
  wire [1:0] _GEN_161; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10755.4]
  wire [1:0] _T_2167_2; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2366.4]
  wire [1:0] _GEN_162; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10760.4]
  wire [2:0] _GEN_163; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10765.4]
  wire [2:0] _T_2167_4; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2512.4]
  wire [2:0] _GEN_164; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10770.4]
  wire [2:0] _T_2167_5; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2588.4]
  wire [2:0] _GEN_165; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10775.4]
  wire [2:0] _T_2167_6; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2666.4]
  wire [2:0] _GEN_166; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10780.4]
  wire [3:0] _GEN_167; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10785.4]
  wire  _T_11334; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@10788.4]
  wire  _T_11335; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@10789.4]
  wire [3:0] _T_2167_8; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2828.4]
  wire [3:0] _GEN_168; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10790.4]
  wire [3:0] _T_2167_9; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2912.4]
  wire [3:0] _GEN_169; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10795.4]
  wire [3:0] _T_2167_10; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2998.4]
  wire [3:0] _GEN_170; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10800.4]
  wire [3:0] _T_2167_11; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3086.4]
  wire [3:0] _GEN_171; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10805.4]
  wire [3:0] _T_2167_12; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3176.4]
  wire [3:0] _GEN_172; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10810.4]
  wire [3:0] _T_2167_13; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3268.4]
  wire [3:0] _GEN_173; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10815.4]
  wire [3:0] _T_2167_14; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3362.4]
  wire [3:0] _GEN_174; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10820.4]
  wire [4:0] _GEN_175; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10825.4]
  wire  _T_11350; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@10828.4]
  wire  _T_11351; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@10829.4]
  wire [4:0] _T_2167_16; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3556.4]
  wire [4:0] _GEN_176; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10830.4]
  wire [4:0] _T_2167_17; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3656.4]
  wire [4:0] _GEN_177; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10835.4]
  wire [4:0] _T_2167_18; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3758.4]
  wire [4:0] _GEN_178; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10840.4]
  wire [4:0] _T_2167_19; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3862.4]
  wire [4:0] _GEN_179; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10845.4]
  wire [4:0] _T_2167_20; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3968.4]
  wire [4:0] _GEN_180; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10850.4]
  wire [4:0] _T_2167_21; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4076.4]
  wire [4:0] _GEN_181; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10855.4]
  wire [4:0] _T_2167_22; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4186.4]
  wire [4:0] _GEN_182; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10860.4]
  wire [4:0] _T_2167_23; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4298.4]
  wire [4:0] _GEN_183; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10865.4]
  wire  _T_11366; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@10868.4]
  wire  _T_11367; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@10869.4]
  wire [4:0] _T_2167_24; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4412.4]
  wire [4:0] _GEN_184; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10870.4]
  wire [4:0] _T_2167_25; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4528.4]
  wire [4:0] _GEN_185; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10875.4]
  wire [4:0] _T_2167_26; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4646.4]
  wire [4:0] _GEN_186; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10880.4]
  wire [4:0] _T_2167_27; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4766.4]
  wire [4:0] _GEN_187; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10885.4]
  wire [4:0] _T_2167_28; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4888.4]
  wire [4:0] _GEN_188; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10890.4]
  wire [4:0] _T_2167_29; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5012.4]
  wire [4:0] _GEN_189; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10895.4]
  wire [4:0] _T_2167_30; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5138.4]
  wire [4:0] _GEN_190; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10900.4]
  wire [5:0] _GEN_191; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10905.4]
  wire  _T_11382; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@10908.4]
  wire  _T_11383; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@10909.4]
  wire [5:0] _T_2167_32; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5396.4]
  wire [5:0] _GEN_192; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10910.4]
  wire [5:0] _T_2167_33; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5528.4]
  wire [5:0] _GEN_193; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10915.4]
  wire [5:0] _T_2167_34; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5662.4]
  wire [5:0] _GEN_194; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10920.4]
  wire [5:0] _T_2167_35; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5798.4]
  wire [5:0] _GEN_195; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10925.4]
  wire [5:0] _T_2167_36; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5936.4]
  wire [5:0] _GEN_196; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10930.4]
  wire [5:0] _T_2167_37; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6076.4]
  wire [5:0] _GEN_197; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10935.4]
  wire [5:0] _T_2167_38; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6218.4]
  wire [5:0] _GEN_198; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10940.4]
  wire [5:0] _T_2167_39; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6362.4]
  wire [5:0] _GEN_199; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10945.4]
  wire  _T_11398; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@10948.4]
  wire  _T_11399; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@10949.4]
  wire [5:0] _T_2167_40; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6508.4]
  wire [5:0] _GEN_200; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10950.4]
  wire [5:0] _T_2167_41; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6656.4]
  wire [5:0] _GEN_201; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10955.4]
  wire [5:0] _T_2167_42; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6806.4]
  wire [5:0] _GEN_202; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10960.4]
  wire [5:0] _T_2167_43; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6958.4]
  wire [5:0] _GEN_203; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10965.4]
  wire [5:0] _T_2167_44; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7112.4]
  wire [5:0] _GEN_204; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10970.4]
  wire [5:0] _T_2167_45; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7268.4]
  wire [5:0] _GEN_205; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10975.4]
  wire [5:0] _T_2167_46; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7426.4]
  wire [5:0] _GEN_206; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10980.4]
  wire [5:0] _T_2167_47; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7586.4]
  wire [5:0] _GEN_207; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10985.4]
  wire  _T_11414; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@10988.4]
  wire  _T_11415; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@10989.4]
  wire [5:0] _T_2167_48; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7748.4]
  wire [5:0] _GEN_208; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10990.4]
  wire [5:0] _T_2167_49; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7912.4]
  wire [5:0] _GEN_209; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10995.4]
  wire [5:0] _T_2167_50; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@8078.4]
  wire [5:0] _GEN_210; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11000.4]
  wire [5:0] _T_2167_51; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@8246.4]
  wire [5:0] _GEN_211; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11005.4]
  wire [5:0] _T_2167_52; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@8416.4]
  wire [5:0] _GEN_212; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11010.4]
  wire [5:0] _T_2167_53; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@8588.4]
  wire [5:0] _GEN_213; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11015.4]
  wire [5:0] _T_2167_54; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@8762.4]
  wire [5:0] _GEN_214; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11020.4]
  wire [5:0] _T_2167_55; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@8938.4]
  wire [5:0] _GEN_215; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11025.4]
  wire  _T_11430; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@11028.4]
  wire  _T_11431; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@11029.4]
  wire [5:0] _T_2167_56; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@9116.4]
  wire [5:0] _GEN_216; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11030.4]
  wire [5:0] _T_2167_57; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@9296.4]
  wire [5:0] _GEN_217; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11035.4]
  wire [5:0] _T_2167_58; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@9478.4]
  wire [5:0] _GEN_218; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11040.4]
  wire [5:0] _T_2167_59; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@9662.4]
  wire [5:0] _GEN_219; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11045.4]
  wire [5:0] _T_2167_60; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@9848.4]
  wire [5:0] _GEN_220; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11050.4]
  wire [5:0] _T_2167_61; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@10036.4]
  wire [5:0] _GEN_221; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11055.4]
  wire [5:0] _T_2167_62; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@10226.4]
  wire [5:0] _GEN_222; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11060.4]
  wire [6:0] _GEN_223; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11065.4]
  wire [7:0] _T_11519; // @[Mux.scala 46:16:@11070.4]
  wire  _T_11523; // @[Mux.scala 46:19:@11072.4]
  wire [7:0] _T_11524; // @[Mux.scala 46:16:@11073.4]
  wire  _T_11525; // @[Mux.scala 46:19:@11074.4]
  wire [7:0] _T_11526; // @[Mux.scala 46:16:@11075.4]
  wire  _T_11531; // @[Mux.scala 46:19:@11077.4]
  wire [7:0] _T_11532; // @[Mux.scala 46:16:@11078.4]
  wire  _T_11533; // @[Mux.scala 46:19:@11079.4]
  wire [7:0] _T_11534; // @[Mux.scala 46:16:@11080.4]
  wire  _T_11535; // @[Mux.scala 46:19:@11081.4]
  wire [7:0] _T_11536; // @[Mux.scala 46:16:@11082.4]
  wire  _T_11542; // @[Mux.scala 46:19:@11084.4]
  wire [7:0] _T_11543; // @[Mux.scala 46:16:@11085.4]
  wire  _T_11544; // @[Mux.scala 46:19:@11086.4]
  wire [7:0] _T_11545; // @[Mux.scala 46:16:@11087.4]
  wire  _T_11546; // @[Mux.scala 46:19:@11088.4]
  wire [7:0] _T_11547; // @[Mux.scala 46:16:@11089.4]
  wire  _T_11548; // @[Mux.scala 46:19:@11090.4]
  wire [7:0] _T_11549; // @[Mux.scala 46:16:@11091.4]
  wire  _T_11556; // @[Mux.scala 46:19:@11093.4]
  wire [7:0] _T_11557; // @[Mux.scala 46:16:@11094.4]
  wire  _T_11558; // @[Mux.scala 46:19:@11095.4]
  wire [7:0] _T_11559; // @[Mux.scala 46:16:@11096.4]
  wire  _T_11560; // @[Mux.scala 46:19:@11097.4]
  wire [7:0] _T_11561; // @[Mux.scala 46:16:@11098.4]
  wire  _T_11562; // @[Mux.scala 46:19:@11099.4]
  wire [7:0] _T_11563; // @[Mux.scala 46:16:@11100.4]
  wire  _T_11564; // @[Mux.scala 46:19:@11101.4]
  wire [7:0] _T_11565; // @[Mux.scala 46:16:@11102.4]
  wire  _T_11573; // @[Mux.scala 46:19:@11104.4]
  wire [7:0] _T_11574; // @[Mux.scala 46:16:@11105.4]
  wire  _T_11575; // @[Mux.scala 46:19:@11106.4]
  wire [7:0] _T_11576; // @[Mux.scala 46:16:@11107.4]
  wire  _T_11577; // @[Mux.scala 46:19:@11108.4]
  wire [7:0] _T_11578; // @[Mux.scala 46:16:@11109.4]
  wire  _T_11579; // @[Mux.scala 46:19:@11110.4]
  wire [7:0] _T_11580; // @[Mux.scala 46:16:@11111.4]
  wire  _T_11581; // @[Mux.scala 46:19:@11112.4]
  wire [7:0] _T_11582; // @[Mux.scala 46:16:@11113.4]
  wire  _T_11583; // @[Mux.scala 46:19:@11114.4]
  wire [7:0] _T_11584; // @[Mux.scala 46:16:@11115.4]
  wire  _T_11593; // @[Mux.scala 46:19:@11117.4]
  wire [7:0] _T_11594; // @[Mux.scala 46:16:@11118.4]
  wire  _T_11595; // @[Mux.scala 46:19:@11119.4]
  wire [7:0] _T_11596; // @[Mux.scala 46:16:@11120.4]
  wire  _T_11597; // @[Mux.scala 46:19:@11121.4]
  wire [7:0] _T_11598; // @[Mux.scala 46:16:@11122.4]
  wire  _T_11599; // @[Mux.scala 46:19:@11123.4]
  wire [7:0] _T_11600; // @[Mux.scala 46:16:@11124.4]
  wire  _T_11601; // @[Mux.scala 46:19:@11125.4]
  wire [7:0] _T_11602; // @[Mux.scala 46:16:@11126.4]
  wire  _T_11603; // @[Mux.scala 46:19:@11127.4]
  wire [7:0] _T_11604; // @[Mux.scala 46:16:@11128.4]
  wire  _T_11605; // @[Mux.scala 46:19:@11129.4]
  wire [7:0] _T_11606; // @[Mux.scala 46:16:@11130.4]
  wire  _T_11616; // @[Mux.scala 46:19:@11132.4]
  wire [7:0] _T_11617; // @[Mux.scala 46:16:@11133.4]
  wire  _T_11618; // @[Mux.scala 46:19:@11134.4]
  wire [7:0] _T_11619; // @[Mux.scala 46:16:@11135.4]
  wire  _T_11620; // @[Mux.scala 46:19:@11136.4]
  wire [7:0] _T_11621; // @[Mux.scala 46:16:@11137.4]
  wire  _T_11622; // @[Mux.scala 46:19:@11138.4]
  wire [7:0] _T_11623; // @[Mux.scala 46:16:@11139.4]
  wire  _T_11624; // @[Mux.scala 46:19:@11140.4]
  wire [7:0] _T_11625; // @[Mux.scala 46:16:@11141.4]
  wire  _T_11626; // @[Mux.scala 46:19:@11142.4]
  wire [7:0] _T_11627; // @[Mux.scala 46:16:@11143.4]
  wire  _T_11628; // @[Mux.scala 46:19:@11144.4]
  wire [7:0] _T_11629; // @[Mux.scala 46:16:@11145.4]
  wire  _T_11630; // @[Mux.scala 46:19:@11146.4]
  wire [7:0] _T_11631; // @[Mux.scala 46:16:@11147.4]
  wire  _T_11642; // @[Mux.scala 46:19:@11149.4]
  wire [7:0] _T_11643; // @[Mux.scala 46:16:@11150.4]
  wire  _T_11644; // @[Mux.scala 46:19:@11151.4]
  wire [7:0] _T_11645; // @[Mux.scala 46:16:@11152.4]
  wire  _T_11646; // @[Mux.scala 46:19:@11153.4]
  wire [7:0] _T_11647; // @[Mux.scala 46:16:@11154.4]
  wire  _T_11648; // @[Mux.scala 46:19:@11155.4]
  wire [7:0] _T_11649; // @[Mux.scala 46:16:@11156.4]
  wire  _T_11650; // @[Mux.scala 46:19:@11157.4]
  wire [7:0] _T_11651; // @[Mux.scala 46:16:@11158.4]
  wire  _T_11652; // @[Mux.scala 46:19:@11159.4]
  wire [7:0] _T_11653; // @[Mux.scala 46:16:@11160.4]
  wire  _T_11654; // @[Mux.scala 46:19:@11161.4]
  wire [7:0] _T_11655; // @[Mux.scala 46:16:@11162.4]
  wire  _T_11656; // @[Mux.scala 46:19:@11163.4]
  wire [7:0] _T_11657; // @[Mux.scala 46:16:@11164.4]
  wire  _T_11658; // @[Mux.scala 46:19:@11165.4]
  wire [7:0] _T_11659; // @[Mux.scala 46:16:@11166.4]
  wire  _T_11671; // @[Mux.scala 46:19:@11168.4]
  wire [7:0] _T_11672; // @[Mux.scala 46:16:@11169.4]
  wire  _T_11673; // @[Mux.scala 46:19:@11170.4]
  wire [7:0] _T_11674; // @[Mux.scala 46:16:@11171.4]
  wire  _T_11675; // @[Mux.scala 46:19:@11172.4]
  wire [7:0] _T_11676; // @[Mux.scala 46:16:@11173.4]
  wire  _T_11677; // @[Mux.scala 46:19:@11174.4]
  wire [7:0] _T_11678; // @[Mux.scala 46:16:@11175.4]
  wire  _T_11679; // @[Mux.scala 46:19:@11176.4]
  wire [7:0] _T_11680; // @[Mux.scala 46:16:@11177.4]
  wire  _T_11681; // @[Mux.scala 46:19:@11178.4]
  wire [7:0] _T_11682; // @[Mux.scala 46:16:@11179.4]
  wire  _T_11683; // @[Mux.scala 46:19:@11180.4]
  wire [7:0] _T_11684; // @[Mux.scala 46:16:@11181.4]
  wire  _T_11685; // @[Mux.scala 46:19:@11182.4]
  wire [7:0] _T_11686; // @[Mux.scala 46:16:@11183.4]
  wire  _T_11687; // @[Mux.scala 46:19:@11184.4]
  wire [7:0] _T_11688; // @[Mux.scala 46:16:@11185.4]
  wire  _T_11689; // @[Mux.scala 46:19:@11186.4]
  wire [7:0] _T_11690; // @[Mux.scala 46:16:@11187.4]
  wire  _T_11703; // @[Mux.scala 46:19:@11189.4]
  wire [7:0] _T_11704; // @[Mux.scala 46:16:@11190.4]
  wire  _T_11705; // @[Mux.scala 46:19:@11191.4]
  wire [7:0] _T_11706; // @[Mux.scala 46:16:@11192.4]
  wire  _T_11707; // @[Mux.scala 46:19:@11193.4]
  wire [7:0] _T_11708; // @[Mux.scala 46:16:@11194.4]
  wire  _T_11709; // @[Mux.scala 46:19:@11195.4]
  wire [7:0] _T_11710; // @[Mux.scala 46:16:@11196.4]
  wire  _T_11711; // @[Mux.scala 46:19:@11197.4]
  wire [7:0] _T_11712; // @[Mux.scala 46:16:@11198.4]
  wire  _T_11713; // @[Mux.scala 46:19:@11199.4]
  wire [7:0] _T_11714; // @[Mux.scala 46:16:@11200.4]
  wire  _T_11715; // @[Mux.scala 46:19:@11201.4]
  wire [7:0] _T_11716; // @[Mux.scala 46:16:@11202.4]
  wire  _T_11717; // @[Mux.scala 46:19:@11203.4]
  wire [7:0] _T_11718; // @[Mux.scala 46:16:@11204.4]
  wire  _T_11719; // @[Mux.scala 46:19:@11205.4]
  wire [7:0] _T_11720; // @[Mux.scala 46:16:@11206.4]
  wire  _T_11721; // @[Mux.scala 46:19:@11207.4]
  wire [7:0] _T_11722; // @[Mux.scala 46:16:@11208.4]
  wire  _T_11723; // @[Mux.scala 46:19:@11209.4]
  wire [7:0] _T_11724; // @[Mux.scala 46:16:@11210.4]
  wire  _T_11738; // @[Mux.scala 46:19:@11212.4]
  wire [7:0] _T_11739; // @[Mux.scala 46:16:@11213.4]
  wire  _T_11740; // @[Mux.scala 46:19:@11214.4]
  wire [7:0] _T_11741; // @[Mux.scala 46:16:@11215.4]
  wire  _T_11742; // @[Mux.scala 46:19:@11216.4]
  wire [7:0] _T_11743; // @[Mux.scala 46:16:@11217.4]
  wire  _T_11744; // @[Mux.scala 46:19:@11218.4]
  wire [7:0] _T_11745; // @[Mux.scala 46:16:@11219.4]
  wire  _T_11746; // @[Mux.scala 46:19:@11220.4]
  wire [7:0] _T_11747; // @[Mux.scala 46:16:@11221.4]
  wire  _T_11748; // @[Mux.scala 46:19:@11222.4]
  wire [7:0] _T_11749; // @[Mux.scala 46:16:@11223.4]
  wire  _T_11750; // @[Mux.scala 46:19:@11224.4]
  wire [7:0] _T_11751; // @[Mux.scala 46:16:@11225.4]
  wire  _T_11752; // @[Mux.scala 46:19:@11226.4]
  wire [7:0] _T_11753; // @[Mux.scala 46:16:@11227.4]
  wire  _T_11754; // @[Mux.scala 46:19:@11228.4]
  wire [7:0] _T_11755; // @[Mux.scala 46:16:@11229.4]
  wire  _T_11756; // @[Mux.scala 46:19:@11230.4]
  wire [7:0] _T_11757; // @[Mux.scala 46:16:@11231.4]
  wire  _T_11758; // @[Mux.scala 46:19:@11232.4]
  wire [7:0] _T_11759; // @[Mux.scala 46:16:@11233.4]
  wire  _T_11760; // @[Mux.scala 46:19:@11234.4]
  wire [7:0] _T_11761; // @[Mux.scala 46:16:@11235.4]
  wire  _T_11776; // @[Mux.scala 46:19:@11237.4]
  wire [7:0] _T_11777; // @[Mux.scala 46:16:@11238.4]
  wire  _T_11778; // @[Mux.scala 46:19:@11239.4]
  wire [7:0] _T_11779; // @[Mux.scala 46:16:@11240.4]
  wire  _T_11780; // @[Mux.scala 46:19:@11241.4]
  wire [7:0] _T_11781; // @[Mux.scala 46:16:@11242.4]
  wire  _T_11782; // @[Mux.scala 46:19:@11243.4]
  wire [7:0] _T_11783; // @[Mux.scala 46:16:@11244.4]
  wire  _T_11784; // @[Mux.scala 46:19:@11245.4]
  wire [7:0] _T_11785; // @[Mux.scala 46:16:@11246.4]
  wire  _T_11786; // @[Mux.scala 46:19:@11247.4]
  wire [7:0] _T_11787; // @[Mux.scala 46:16:@11248.4]
  wire  _T_11788; // @[Mux.scala 46:19:@11249.4]
  wire [7:0] _T_11789; // @[Mux.scala 46:16:@11250.4]
  wire  _T_11790; // @[Mux.scala 46:19:@11251.4]
  wire [7:0] _T_11791; // @[Mux.scala 46:16:@11252.4]
  wire  _T_11792; // @[Mux.scala 46:19:@11253.4]
  wire [7:0] _T_11793; // @[Mux.scala 46:16:@11254.4]
  wire  _T_11794; // @[Mux.scala 46:19:@11255.4]
  wire [7:0] _T_11795; // @[Mux.scala 46:16:@11256.4]
  wire  _T_11796; // @[Mux.scala 46:19:@11257.4]
  wire [7:0] _T_11797; // @[Mux.scala 46:16:@11258.4]
  wire  _T_11798; // @[Mux.scala 46:19:@11259.4]
  wire [7:0] _T_11799; // @[Mux.scala 46:16:@11260.4]
  wire  _T_11800; // @[Mux.scala 46:19:@11261.4]
  wire [7:0] _T_11801; // @[Mux.scala 46:16:@11262.4]
  wire  _T_11817; // @[Mux.scala 46:19:@11264.4]
  wire [7:0] _T_11818; // @[Mux.scala 46:16:@11265.4]
  wire  _T_11819; // @[Mux.scala 46:19:@11266.4]
  wire [7:0] _T_11820; // @[Mux.scala 46:16:@11267.4]
  wire  _T_11821; // @[Mux.scala 46:19:@11268.4]
  wire [7:0] _T_11822; // @[Mux.scala 46:16:@11269.4]
  wire  _T_11823; // @[Mux.scala 46:19:@11270.4]
  wire [7:0] _T_11824; // @[Mux.scala 46:16:@11271.4]
  wire  _T_11825; // @[Mux.scala 46:19:@11272.4]
  wire [7:0] _T_11826; // @[Mux.scala 46:16:@11273.4]
  wire  _T_11827; // @[Mux.scala 46:19:@11274.4]
  wire [7:0] _T_11828; // @[Mux.scala 46:16:@11275.4]
  wire  _T_11829; // @[Mux.scala 46:19:@11276.4]
  wire [7:0] _T_11830; // @[Mux.scala 46:16:@11277.4]
  wire  _T_11831; // @[Mux.scala 46:19:@11278.4]
  wire [7:0] _T_11832; // @[Mux.scala 46:16:@11279.4]
  wire  _T_11833; // @[Mux.scala 46:19:@11280.4]
  wire [7:0] _T_11834; // @[Mux.scala 46:16:@11281.4]
  wire  _T_11835; // @[Mux.scala 46:19:@11282.4]
  wire [7:0] _T_11836; // @[Mux.scala 46:16:@11283.4]
  wire  _T_11837; // @[Mux.scala 46:19:@11284.4]
  wire [7:0] _T_11838; // @[Mux.scala 46:16:@11285.4]
  wire  _T_11839; // @[Mux.scala 46:19:@11286.4]
  wire [7:0] _T_11840; // @[Mux.scala 46:16:@11287.4]
  wire  _T_11841; // @[Mux.scala 46:19:@11288.4]
  wire [7:0] _T_11842; // @[Mux.scala 46:16:@11289.4]
  wire  _T_11843; // @[Mux.scala 46:19:@11290.4]
  wire [7:0] _T_11844; // @[Mux.scala 46:16:@11291.4]
  wire  _T_11861; // @[Mux.scala 46:19:@11293.4]
  wire [7:0] _T_11862; // @[Mux.scala 46:16:@11294.4]
  wire  _T_11863; // @[Mux.scala 46:19:@11295.4]
  wire [7:0] _T_11864; // @[Mux.scala 46:16:@11296.4]
  wire  _T_11865; // @[Mux.scala 46:19:@11297.4]
  wire [7:0] _T_11866; // @[Mux.scala 46:16:@11298.4]
  wire  _T_11867; // @[Mux.scala 46:19:@11299.4]
  wire [7:0] _T_11868; // @[Mux.scala 46:16:@11300.4]
  wire  _T_11869; // @[Mux.scala 46:19:@11301.4]
  wire [7:0] _T_11870; // @[Mux.scala 46:16:@11302.4]
  wire  _T_11871; // @[Mux.scala 46:19:@11303.4]
  wire [7:0] _T_11872; // @[Mux.scala 46:16:@11304.4]
  wire  _T_11873; // @[Mux.scala 46:19:@11305.4]
  wire [7:0] _T_11874; // @[Mux.scala 46:16:@11306.4]
  wire  _T_11875; // @[Mux.scala 46:19:@11307.4]
  wire [7:0] _T_11876; // @[Mux.scala 46:16:@11308.4]
  wire  _T_11877; // @[Mux.scala 46:19:@11309.4]
  wire [7:0] _T_11878; // @[Mux.scala 46:16:@11310.4]
  wire  _T_11879; // @[Mux.scala 46:19:@11311.4]
  wire [7:0] _T_11880; // @[Mux.scala 46:16:@11312.4]
  wire  _T_11881; // @[Mux.scala 46:19:@11313.4]
  wire [7:0] _T_11882; // @[Mux.scala 46:16:@11314.4]
  wire  _T_11883; // @[Mux.scala 46:19:@11315.4]
  wire [7:0] _T_11884; // @[Mux.scala 46:16:@11316.4]
  wire  _T_11885; // @[Mux.scala 46:19:@11317.4]
  wire [7:0] _T_11886; // @[Mux.scala 46:16:@11318.4]
  wire  _T_11887; // @[Mux.scala 46:19:@11319.4]
  wire [7:0] _T_11888; // @[Mux.scala 46:16:@11320.4]
  wire  _T_11889; // @[Mux.scala 46:19:@11321.4]
  wire [7:0] _T_11890; // @[Mux.scala 46:16:@11322.4]
  wire  _T_11908; // @[Mux.scala 46:19:@11324.4]
  wire [7:0] _T_11909; // @[Mux.scala 46:16:@11325.4]
  wire  _T_11910; // @[Mux.scala 46:19:@11326.4]
  wire [7:0] _T_11911; // @[Mux.scala 46:16:@11327.4]
  wire  _T_11912; // @[Mux.scala 46:19:@11328.4]
  wire [7:0] _T_11913; // @[Mux.scala 46:16:@11329.4]
  wire  _T_11914; // @[Mux.scala 46:19:@11330.4]
  wire [7:0] _T_11915; // @[Mux.scala 46:16:@11331.4]
  wire  _T_11916; // @[Mux.scala 46:19:@11332.4]
  wire [7:0] _T_11917; // @[Mux.scala 46:16:@11333.4]
  wire  _T_11918; // @[Mux.scala 46:19:@11334.4]
  wire [7:0] _T_11919; // @[Mux.scala 46:16:@11335.4]
  wire  _T_11920; // @[Mux.scala 46:19:@11336.4]
  wire [7:0] _T_11921; // @[Mux.scala 46:16:@11337.4]
  wire  _T_11922; // @[Mux.scala 46:19:@11338.4]
  wire [7:0] _T_11923; // @[Mux.scala 46:16:@11339.4]
  wire  _T_11924; // @[Mux.scala 46:19:@11340.4]
  wire [7:0] _T_11925; // @[Mux.scala 46:16:@11341.4]
  wire  _T_11926; // @[Mux.scala 46:19:@11342.4]
  wire [7:0] _T_11927; // @[Mux.scala 46:16:@11343.4]
  wire  _T_11928; // @[Mux.scala 46:19:@11344.4]
  wire [7:0] _T_11929; // @[Mux.scala 46:16:@11345.4]
  wire  _T_11930; // @[Mux.scala 46:19:@11346.4]
  wire [7:0] _T_11931; // @[Mux.scala 46:16:@11347.4]
  wire  _T_11932; // @[Mux.scala 46:19:@11348.4]
  wire [7:0] _T_11933; // @[Mux.scala 46:16:@11349.4]
  wire  _T_11934; // @[Mux.scala 46:19:@11350.4]
  wire [7:0] _T_11935; // @[Mux.scala 46:16:@11351.4]
  wire  _T_11936; // @[Mux.scala 46:19:@11352.4]
  wire [7:0] _T_11937; // @[Mux.scala 46:16:@11353.4]
  wire  _T_11938; // @[Mux.scala 46:19:@11354.4]
  wire [7:0] _T_11939; // @[Mux.scala 46:16:@11355.4]
  wire  _T_11958; // @[Mux.scala 46:19:@11357.4]
  wire [7:0] _T_11959; // @[Mux.scala 46:16:@11358.4]
  wire  _T_11960; // @[Mux.scala 46:19:@11359.4]
  wire [7:0] _T_11961; // @[Mux.scala 46:16:@11360.4]
  wire  _T_11962; // @[Mux.scala 46:19:@11361.4]
  wire [7:0] _T_11963; // @[Mux.scala 46:16:@11362.4]
  wire  _T_11964; // @[Mux.scala 46:19:@11363.4]
  wire [7:0] _T_11965; // @[Mux.scala 46:16:@11364.4]
  wire  _T_11966; // @[Mux.scala 46:19:@11365.4]
  wire [7:0] _T_11967; // @[Mux.scala 46:16:@11366.4]
  wire  _T_11968; // @[Mux.scala 46:19:@11367.4]
  wire [7:0] _T_11969; // @[Mux.scala 46:16:@11368.4]
  wire  _T_11970; // @[Mux.scala 46:19:@11369.4]
  wire [7:0] _T_11971; // @[Mux.scala 46:16:@11370.4]
  wire  _T_11972; // @[Mux.scala 46:19:@11371.4]
  wire [7:0] _T_11973; // @[Mux.scala 46:16:@11372.4]
  wire  _T_11974; // @[Mux.scala 46:19:@11373.4]
  wire [7:0] _T_11975; // @[Mux.scala 46:16:@11374.4]
  wire  _T_11976; // @[Mux.scala 46:19:@11375.4]
  wire [7:0] _T_11977; // @[Mux.scala 46:16:@11376.4]
  wire  _T_11978; // @[Mux.scala 46:19:@11377.4]
  wire [7:0] _T_11979; // @[Mux.scala 46:16:@11378.4]
  wire  _T_11980; // @[Mux.scala 46:19:@11379.4]
  wire [7:0] _T_11981; // @[Mux.scala 46:16:@11380.4]
  wire  _T_11982; // @[Mux.scala 46:19:@11381.4]
  wire [7:0] _T_11983; // @[Mux.scala 46:16:@11382.4]
  wire  _T_11984; // @[Mux.scala 46:19:@11383.4]
  wire [7:0] _T_11985; // @[Mux.scala 46:16:@11384.4]
  wire  _T_11986; // @[Mux.scala 46:19:@11385.4]
  wire [7:0] _T_11987; // @[Mux.scala 46:16:@11386.4]
  wire  _T_11988; // @[Mux.scala 46:19:@11387.4]
  wire [7:0] _T_11989; // @[Mux.scala 46:16:@11388.4]
  wire  _T_11990; // @[Mux.scala 46:19:@11389.4]
  wire [7:0] _T_11991; // @[Mux.scala 46:16:@11390.4]
  wire  _T_12011; // @[Mux.scala 46:19:@11392.4]
  wire [7:0] _T_12012; // @[Mux.scala 46:16:@11393.4]
  wire  _T_12013; // @[Mux.scala 46:19:@11394.4]
  wire [7:0] _T_12014; // @[Mux.scala 46:16:@11395.4]
  wire  _T_12015; // @[Mux.scala 46:19:@11396.4]
  wire [7:0] _T_12016; // @[Mux.scala 46:16:@11397.4]
  wire  _T_12017; // @[Mux.scala 46:19:@11398.4]
  wire [7:0] _T_12018; // @[Mux.scala 46:16:@11399.4]
  wire  _T_12019; // @[Mux.scala 46:19:@11400.4]
  wire [7:0] _T_12020; // @[Mux.scala 46:16:@11401.4]
  wire  _T_12021; // @[Mux.scala 46:19:@11402.4]
  wire [7:0] _T_12022; // @[Mux.scala 46:16:@11403.4]
  wire  _T_12023; // @[Mux.scala 46:19:@11404.4]
  wire [7:0] _T_12024; // @[Mux.scala 46:16:@11405.4]
  wire  _T_12025; // @[Mux.scala 46:19:@11406.4]
  wire [7:0] _T_12026; // @[Mux.scala 46:16:@11407.4]
  wire  _T_12027; // @[Mux.scala 46:19:@11408.4]
  wire [7:0] _T_12028; // @[Mux.scala 46:16:@11409.4]
  wire  _T_12029; // @[Mux.scala 46:19:@11410.4]
  wire [7:0] _T_12030; // @[Mux.scala 46:16:@11411.4]
  wire  _T_12031; // @[Mux.scala 46:19:@11412.4]
  wire [7:0] _T_12032; // @[Mux.scala 46:16:@11413.4]
  wire  _T_12033; // @[Mux.scala 46:19:@11414.4]
  wire [7:0] _T_12034; // @[Mux.scala 46:16:@11415.4]
  wire  _T_12035; // @[Mux.scala 46:19:@11416.4]
  wire [7:0] _T_12036; // @[Mux.scala 46:16:@11417.4]
  wire  _T_12037; // @[Mux.scala 46:19:@11418.4]
  wire [7:0] _T_12038; // @[Mux.scala 46:16:@11419.4]
  wire  _T_12039; // @[Mux.scala 46:19:@11420.4]
  wire [7:0] _T_12040; // @[Mux.scala 46:16:@11421.4]
  wire  _T_12041; // @[Mux.scala 46:19:@11422.4]
  wire [7:0] _T_12042; // @[Mux.scala 46:16:@11423.4]
  wire  _T_12043; // @[Mux.scala 46:19:@11424.4]
  wire [7:0] _T_12044; // @[Mux.scala 46:16:@11425.4]
  wire  _T_12045; // @[Mux.scala 46:19:@11426.4]
  wire [7:0] _T_12046; // @[Mux.scala 46:16:@11427.4]
  wire  _T_12067; // @[Mux.scala 46:19:@11429.4]
  wire [7:0] _T_12068; // @[Mux.scala 46:16:@11430.4]
  wire  _T_12069; // @[Mux.scala 46:19:@11431.4]
  wire [7:0] _T_12070; // @[Mux.scala 46:16:@11432.4]
  wire  _T_12071; // @[Mux.scala 46:19:@11433.4]
  wire [7:0] _T_12072; // @[Mux.scala 46:16:@11434.4]
  wire  _T_12073; // @[Mux.scala 46:19:@11435.4]
  wire [7:0] _T_12074; // @[Mux.scala 46:16:@11436.4]
  wire  _T_12075; // @[Mux.scala 46:19:@11437.4]
  wire [7:0] _T_12076; // @[Mux.scala 46:16:@11438.4]
  wire  _T_12077; // @[Mux.scala 46:19:@11439.4]
  wire [7:0] _T_12078; // @[Mux.scala 46:16:@11440.4]
  wire  _T_12079; // @[Mux.scala 46:19:@11441.4]
  wire [7:0] _T_12080; // @[Mux.scala 46:16:@11442.4]
  wire  _T_12081; // @[Mux.scala 46:19:@11443.4]
  wire [7:0] _T_12082; // @[Mux.scala 46:16:@11444.4]
  wire  _T_12083; // @[Mux.scala 46:19:@11445.4]
  wire [7:0] _T_12084; // @[Mux.scala 46:16:@11446.4]
  wire  _T_12085; // @[Mux.scala 46:19:@11447.4]
  wire [7:0] _T_12086; // @[Mux.scala 46:16:@11448.4]
  wire  _T_12087; // @[Mux.scala 46:19:@11449.4]
  wire [7:0] _T_12088; // @[Mux.scala 46:16:@11450.4]
  wire  _T_12089; // @[Mux.scala 46:19:@11451.4]
  wire [7:0] _T_12090; // @[Mux.scala 46:16:@11452.4]
  wire  _T_12091; // @[Mux.scala 46:19:@11453.4]
  wire [7:0] _T_12092; // @[Mux.scala 46:16:@11454.4]
  wire  _T_12093; // @[Mux.scala 46:19:@11455.4]
  wire [7:0] _T_12094; // @[Mux.scala 46:16:@11456.4]
  wire  _T_12095; // @[Mux.scala 46:19:@11457.4]
  wire [7:0] _T_12096; // @[Mux.scala 46:16:@11458.4]
  wire  _T_12097; // @[Mux.scala 46:19:@11459.4]
  wire [7:0] _T_12098; // @[Mux.scala 46:16:@11460.4]
  wire  _T_12099; // @[Mux.scala 46:19:@11461.4]
  wire [7:0] _T_12100; // @[Mux.scala 46:16:@11462.4]
  wire  _T_12101; // @[Mux.scala 46:19:@11463.4]
  wire [7:0] _T_12102; // @[Mux.scala 46:16:@11464.4]
  wire  _T_12103; // @[Mux.scala 46:19:@11465.4]
  wire [7:0] _T_12104; // @[Mux.scala 46:16:@11466.4]
  wire  _T_12126; // @[Mux.scala 46:19:@11468.4]
  wire [7:0] _T_12127; // @[Mux.scala 46:16:@11469.4]
  wire  _T_12128; // @[Mux.scala 46:19:@11470.4]
  wire [7:0] _T_12129; // @[Mux.scala 46:16:@11471.4]
  wire  _T_12130; // @[Mux.scala 46:19:@11472.4]
  wire [7:0] _T_12131; // @[Mux.scala 46:16:@11473.4]
  wire  _T_12132; // @[Mux.scala 46:19:@11474.4]
  wire [7:0] _T_12133; // @[Mux.scala 46:16:@11475.4]
  wire  _T_12134; // @[Mux.scala 46:19:@11476.4]
  wire [7:0] _T_12135; // @[Mux.scala 46:16:@11477.4]
  wire  _T_12136; // @[Mux.scala 46:19:@11478.4]
  wire [7:0] _T_12137; // @[Mux.scala 46:16:@11479.4]
  wire  _T_12138; // @[Mux.scala 46:19:@11480.4]
  wire [7:0] _T_12139; // @[Mux.scala 46:16:@11481.4]
  wire  _T_12140; // @[Mux.scala 46:19:@11482.4]
  wire [7:0] _T_12141; // @[Mux.scala 46:16:@11483.4]
  wire  _T_12142; // @[Mux.scala 46:19:@11484.4]
  wire [7:0] _T_12143; // @[Mux.scala 46:16:@11485.4]
  wire  _T_12144; // @[Mux.scala 46:19:@11486.4]
  wire [7:0] _T_12145; // @[Mux.scala 46:16:@11487.4]
  wire  _T_12146; // @[Mux.scala 46:19:@11488.4]
  wire [7:0] _T_12147; // @[Mux.scala 46:16:@11489.4]
  wire  _T_12148; // @[Mux.scala 46:19:@11490.4]
  wire [7:0] _T_12149; // @[Mux.scala 46:16:@11491.4]
  wire  _T_12150; // @[Mux.scala 46:19:@11492.4]
  wire [7:0] _T_12151; // @[Mux.scala 46:16:@11493.4]
  wire  _T_12152; // @[Mux.scala 46:19:@11494.4]
  wire [7:0] _T_12153; // @[Mux.scala 46:16:@11495.4]
  wire  _T_12154; // @[Mux.scala 46:19:@11496.4]
  wire [7:0] _T_12155; // @[Mux.scala 46:16:@11497.4]
  wire  _T_12156; // @[Mux.scala 46:19:@11498.4]
  wire [7:0] _T_12157; // @[Mux.scala 46:16:@11499.4]
  wire  _T_12158; // @[Mux.scala 46:19:@11500.4]
  wire [7:0] _T_12159; // @[Mux.scala 46:16:@11501.4]
  wire  _T_12160; // @[Mux.scala 46:19:@11502.4]
  wire [7:0] _T_12161; // @[Mux.scala 46:16:@11503.4]
  wire  _T_12162; // @[Mux.scala 46:19:@11504.4]
  wire [7:0] _T_12163; // @[Mux.scala 46:16:@11505.4]
  wire  _T_12164; // @[Mux.scala 46:19:@11506.4]
  wire [7:0] _T_12165; // @[Mux.scala 46:16:@11507.4]
  wire  _T_12188; // @[Mux.scala 46:19:@11509.4]
  wire [7:0] _T_12189; // @[Mux.scala 46:16:@11510.4]
  wire  _T_12190; // @[Mux.scala 46:19:@11511.4]
  wire [7:0] _T_12191; // @[Mux.scala 46:16:@11512.4]
  wire  _T_12192; // @[Mux.scala 46:19:@11513.4]
  wire [7:0] _T_12193; // @[Mux.scala 46:16:@11514.4]
  wire  _T_12194; // @[Mux.scala 46:19:@11515.4]
  wire [7:0] _T_12195; // @[Mux.scala 46:16:@11516.4]
  wire  _T_12196; // @[Mux.scala 46:19:@11517.4]
  wire [7:0] _T_12197; // @[Mux.scala 46:16:@11518.4]
  wire  _T_12198; // @[Mux.scala 46:19:@11519.4]
  wire [7:0] _T_12199; // @[Mux.scala 46:16:@11520.4]
  wire  _T_12200; // @[Mux.scala 46:19:@11521.4]
  wire [7:0] _T_12201; // @[Mux.scala 46:16:@11522.4]
  wire  _T_12202; // @[Mux.scala 46:19:@11523.4]
  wire [7:0] _T_12203; // @[Mux.scala 46:16:@11524.4]
  wire  _T_12204; // @[Mux.scala 46:19:@11525.4]
  wire [7:0] _T_12205; // @[Mux.scala 46:16:@11526.4]
  wire  _T_12206; // @[Mux.scala 46:19:@11527.4]
  wire [7:0] _T_12207; // @[Mux.scala 46:16:@11528.4]
  wire  _T_12208; // @[Mux.scala 46:19:@11529.4]
  wire [7:0] _T_12209; // @[Mux.scala 46:16:@11530.4]
  wire  _T_12210; // @[Mux.scala 46:19:@11531.4]
  wire [7:0] _T_12211; // @[Mux.scala 46:16:@11532.4]
  wire  _T_12212; // @[Mux.scala 46:19:@11533.4]
  wire [7:0] _T_12213; // @[Mux.scala 46:16:@11534.4]
  wire  _T_12214; // @[Mux.scala 46:19:@11535.4]
  wire [7:0] _T_12215; // @[Mux.scala 46:16:@11536.4]
  wire  _T_12216; // @[Mux.scala 46:19:@11537.4]
  wire [7:0] _T_12217; // @[Mux.scala 46:16:@11538.4]
  wire  _T_12218; // @[Mux.scala 46:19:@11539.4]
  wire [7:0] _T_12219; // @[Mux.scala 46:16:@11540.4]
  wire  _T_12220; // @[Mux.scala 46:19:@11541.4]
  wire [7:0] _T_12221; // @[Mux.scala 46:16:@11542.4]
  wire  _T_12222; // @[Mux.scala 46:19:@11543.4]
  wire [7:0] _T_12223; // @[Mux.scala 46:16:@11544.4]
  wire  _T_12224; // @[Mux.scala 46:19:@11545.4]
  wire [7:0] _T_12225; // @[Mux.scala 46:16:@11546.4]
  wire  _T_12226; // @[Mux.scala 46:19:@11547.4]
  wire [7:0] _T_12227; // @[Mux.scala 46:16:@11548.4]
  wire  _T_12228; // @[Mux.scala 46:19:@11549.4]
  wire [7:0] _T_12229; // @[Mux.scala 46:16:@11550.4]
  wire  _T_12253; // @[Mux.scala 46:19:@11552.4]
  wire [7:0] _T_12254; // @[Mux.scala 46:16:@11553.4]
  wire  _T_12255; // @[Mux.scala 46:19:@11554.4]
  wire [7:0] _T_12256; // @[Mux.scala 46:16:@11555.4]
  wire  _T_12257; // @[Mux.scala 46:19:@11556.4]
  wire [7:0] _T_12258; // @[Mux.scala 46:16:@11557.4]
  wire  _T_12259; // @[Mux.scala 46:19:@11558.4]
  wire [7:0] _T_12260; // @[Mux.scala 46:16:@11559.4]
  wire  _T_12261; // @[Mux.scala 46:19:@11560.4]
  wire [7:0] _T_12262; // @[Mux.scala 46:16:@11561.4]
  wire  _T_12263; // @[Mux.scala 46:19:@11562.4]
  wire [7:0] _T_12264; // @[Mux.scala 46:16:@11563.4]
  wire  _T_12265; // @[Mux.scala 46:19:@11564.4]
  wire [7:0] _T_12266; // @[Mux.scala 46:16:@11565.4]
  wire  _T_12267; // @[Mux.scala 46:19:@11566.4]
  wire [7:0] _T_12268; // @[Mux.scala 46:16:@11567.4]
  wire  _T_12269; // @[Mux.scala 46:19:@11568.4]
  wire [7:0] _T_12270; // @[Mux.scala 46:16:@11569.4]
  wire  _T_12271; // @[Mux.scala 46:19:@11570.4]
  wire [7:0] _T_12272; // @[Mux.scala 46:16:@11571.4]
  wire  _T_12273; // @[Mux.scala 46:19:@11572.4]
  wire [7:0] _T_12274; // @[Mux.scala 46:16:@11573.4]
  wire  _T_12275; // @[Mux.scala 46:19:@11574.4]
  wire [7:0] _T_12276; // @[Mux.scala 46:16:@11575.4]
  wire  _T_12277; // @[Mux.scala 46:19:@11576.4]
  wire [7:0] _T_12278; // @[Mux.scala 46:16:@11577.4]
  wire  _T_12279; // @[Mux.scala 46:19:@11578.4]
  wire [7:0] _T_12280; // @[Mux.scala 46:16:@11579.4]
  wire  _T_12281; // @[Mux.scala 46:19:@11580.4]
  wire [7:0] _T_12282; // @[Mux.scala 46:16:@11581.4]
  wire  _T_12283; // @[Mux.scala 46:19:@11582.4]
  wire [7:0] _T_12284; // @[Mux.scala 46:16:@11583.4]
  wire  _T_12285; // @[Mux.scala 46:19:@11584.4]
  wire [7:0] _T_12286; // @[Mux.scala 46:16:@11585.4]
  wire  _T_12287; // @[Mux.scala 46:19:@11586.4]
  wire [7:0] _T_12288; // @[Mux.scala 46:16:@11587.4]
  wire  _T_12289; // @[Mux.scala 46:19:@11588.4]
  wire [7:0] _T_12290; // @[Mux.scala 46:16:@11589.4]
  wire  _T_12291; // @[Mux.scala 46:19:@11590.4]
  wire [7:0] _T_12292; // @[Mux.scala 46:16:@11591.4]
  wire  _T_12293; // @[Mux.scala 46:19:@11592.4]
  wire [7:0] _T_12294; // @[Mux.scala 46:16:@11593.4]
  wire  _T_12295; // @[Mux.scala 46:19:@11594.4]
  wire [7:0] _T_12296; // @[Mux.scala 46:16:@11595.4]
  wire  _T_12321; // @[Mux.scala 46:19:@11597.4]
  wire [7:0] _T_12322; // @[Mux.scala 46:16:@11598.4]
  wire  _T_12323; // @[Mux.scala 46:19:@11599.4]
  wire [7:0] _T_12324; // @[Mux.scala 46:16:@11600.4]
  wire  _T_12325; // @[Mux.scala 46:19:@11601.4]
  wire [7:0] _T_12326; // @[Mux.scala 46:16:@11602.4]
  wire  _T_12327; // @[Mux.scala 46:19:@11603.4]
  wire [7:0] _T_12328; // @[Mux.scala 46:16:@11604.4]
  wire  _T_12329; // @[Mux.scala 46:19:@11605.4]
  wire [7:0] _T_12330; // @[Mux.scala 46:16:@11606.4]
  wire  _T_12331; // @[Mux.scala 46:19:@11607.4]
  wire [7:0] _T_12332; // @[Mux.scala 46:16:@11608.4]
  wire  _T_12333; // @[Mux.scala 46:19:@11609.4]
  wire [7:0] _T_12334; // @[Mux.scala 46:16:@11610.4]
  wire  _T_12335; // @[Mux.scala 46:19:@11611.4]
  wire [7:0] _T_12336; // @[Mux.scala 46:16:@11612.4]
  wire  _T_12337; // @[Mux.scala 46:19:@11613.4]
  wire [7:0] _T_12338; // @[Mux.scala 46:16:@11614.4]
  wire  _T_12339; // @[Mux.scala 46:19:@11615.4]
  wire [7:0] _T_12340; // @[Mux.scala 46:16:@11616.4]
  wire  _T_12341; // @[Mux.scala 46:19:@11617.4]
  wire [7:0] _T_12342; // @[Mux.scala 46:16:@11618.4]
  wire  _T_12343; // @[Mux.scala 46:19:@11619.4]
  wire [7:0] _T_12344; // @[Mux.scala 46:16:@11620.4]
  wire  _T_12345; // @[Mux.scala 46:19:@11621.4]
  wire [7:0] _T_12346; // @[Mux.scala 46:16:@11622.4]
  wire  _T_12347; // @[Mux.scala 46:19:@11623.4]
  wire [7:0] _T_12348; // @[Mux.scala 46:16:@11624.4]
  wire  _T_12349; // @[Mux.scala 46:19:@11625.4]
  wire [7:0] _T_12350; // @[Mux.scala 46:16:@11626.4]
  wire  _T_12351; // @[Mux.scala 46:19:@11627.4]
  wire [7:0] _T_12352; // @[Mux.scala 46:16:@11628.4]
  wire  _T_12353; // @[Mux.scala 46:19:@11629.4]
  wire [7:0] _T_12354; // @[Mux.scala 46:16:@11630.4]
  wire  _T_12355; // @[Mux.scala 46:19:@11631.4]
  wire [7:0] _T_12356; // @[Mux.scala 46:16:@11632.4]
  wire  _T_12357; // @[Mux.scala 46:19:@11633.4]
  wire [7:0] _T_12358; // @[Mux.scala 46:16:@11634.4]
  wire  _T_12359; // @[Mux.scala 46:19:@11635.4]
  wire [7:0] _T_12360; // @[Mux.scala 46:16:@11636.4]
  wire  _T_12361; // @[Mux.scala 46:19:@11637.4]
  wire [7:0] _T_12362; // @[Mux.scala 46:16:@11638.4]
  wire  _T_12363; // @[Mux.scala 46:19:@11639.4]
  wire [7:0] _T_12364; // @[Mux.scala 46:16:@11640.4]
  wire  _T_12365; // @[Mux.scala 46:19:@11641.4]
  wire [7:0] _T_12366; // @[Mux.scala 46:16:@11642.4]
  wire  _T_12392; // @[Mux.scala 46:19:@11644.4]
  wire [7:0] _T_12393; // @[Mux.scala 46:16:@11645.4]
  wire  _T_12394; // @[Mux.scala 46:19:@11646.4]
  wire [7:0] _T_12395; // @[Mux.scala 46:16:@11647.4]
  wire  _T_12396; // @[Mux.scala 46:19:@11648.4]
  wire [7:0] _T_12397; // @[Mux.scala 46:16:@11649.4]
  wire  _T_12398; // @[Mux.scala 46:19:@11650.4]
  wire [7:0] _T_12399; // @[Mux.scala 46:16:@11651.4]
  wire  _T_12400; // @[Mux.scala 46:19:@11652.4]
  wire [7:0] _T_12401; // @[Mux.scala 46:16:@11653.4]
  wire  _T_12402; // @[Mux.scala 46:19:@11654.4]
  wire [7:0] _T_12403; // @[Mux.scala 46:16:@11655.4]
  wire  _T_12404; // @[Mux.scala 46:19:@11656.4]
  wire [7:0] _T_12405; // @[Mux.scala 46:16:@11657.4]
  wire  _T_12406; // @[Mux.scala 46:19:@11658.4]
  wire [7:0] _T_12407; // @[Mux.scala 46:16:@11659.4]
  wire  _T_12408; // @[Mux.scala 46:19:@11660.4]
  wire [7:0] _T_12409; // @[Mux.scala 46:16:@11661.4]
  wire  _T_12410; // @[Mux.scala 46:19:@11662.4]
  wire [7:0] _T_12411; // @[Mux.scala 46:16:@11663.4]
  wire  _T_12412; // @[Mux.scala 46:19:@11664.4]
  wire [7:0] _T_12413; // @[Mux.scala 46:16:@11665.4]
  wire  _T_12414; // @[Mux.scala 46:19:@11666.4]
  wire [7:0] _T_12415; // @[Mux.scala 46:16:@11667.4]
  wire  _T_12416; // @[Mux.scala 46:19:@11668.4]
  wire [7:0] _T_12417; // @[Mux.scala 46:16:@11669.4]
  wire  _T_12418; // @[Mux.scala 46:19:@11670.4]
  wire [7:0] _T_12419; // @[Mux.scala 46:16:@11671.4]
  wire  _T_12420; // @[Mux.scala 46:19:@11672.4]
  wire [7:0] _T_12421; // @[Mux.scala 46:16:@11673.4]
  wire  _T_12422; // @[Mux.scala 46:19:@11674.4]
  wire [7:0] _T_12423; // @[Mux.scala 46:16:@11675.4]
  wire  _T_12424; // @[Mux.scala 46:19:@11676.4]
  wire [7:0] _T_12425; // @[Mux.scala 46:16:@11677.4]
  wire  _T_12426; // @[Mux.scala 46:19:@11678.4]
  wire [7:0] _T_12427; // @[Mux.scala 46:16:@11679.4]
  wire  _T_12428; // @[Mux.scala 46:19:@11680.4]
  wire [7:0] _T_12429; // @[Mux.scala 46:16:@11681.4]
  wire  _T_12430; // @[Mux.scala 46:19:@11682.4]
  wire [7:0] _T_12431; // @[Mux.scala 46:16:@11683.4]
  wire  _T_12432; // @[Mux.scala 46:19:@11684.4]
  wire [7:0] _T_12433; // @[Mux.scala 46:16:@11685.4]
  wire  _T_12434; // @[Mux.scala 46:19:@11686.4]
  wire [7:0] _T_12435; // @[Mux.scala 46:16:@11687.4]
  wire  _T_12436; // @[Mux.scala 46:19:@11688.4]
  wire [7:0] _T_12437; // @[Mux.scala 46:16:@11689.4]
  wire  _T_12438; // @[Mux.scala 46:19:@11690.4]
  wire [7:0] _T_12439; // @[Mux.scala 46:16:@11691.4]
  wire  _T_12466; // @[Mux.scala 46:19:@11693.4]
  wire [7:0] _T_12467; // @[Mux.scala 46:16:@11694.4]
  wire  _T_12468; // @[Mux.scala 46:19:@11695.4]
  wire [7:0] _T_12469; // @[Mux.scala 46:16:@11696.4]
  wire  _T_12470; // @[Mux.scala 46:19:@11697.4]
  wire [7:0] _T_12471; // @[Mux.scala 46:16:@11698.4]
  wire  _T_12472; // @[Mux.scala 46:19:@11699.4]
  wire [7:0] _T_12473; // @[Mux.scala 46:16:@11700.4]
  wire  _T_12474; // @[Mux.scala 46:19:@11701.4]
  wire [7:0] _T_12475; // @[Mux.scala 46:16:@11702.4]
  wire  _T_12476; // @[Mux.scala 46:19:@11703.4]
  wire [7:0] _T_12477; // @[Mux.scala 46:16:@11704.4]
  wire  _T_12478; // @[Mux.scala 46:19:@11705.4]
  wire [7:0] _T_12479; // @[Mux.scala 46:16:@11706.4]
  wire  _T_12480; // @[Mux.scala 46:19:@11707.4]
  wire [7:0] _T_12481; // @[Mux.scala 46:16:@11708.4]
  wire  _T_12482; // @[Mux.scala 46:19:@11709.4]
  wire [7:0] _T_12483; // @[Mux.scala 46:16:@11710.4]
  wire  _T_12484; // @[Mux.scala 46:19:@11711.4]
  wire [7:0] _T_12485; // @[Mux.scala 46:16:@11712.4]
  wire  _T_12486; // @[Mux.scala 46:19:@11713.4]
  wire [7:0] _T_12487; // @[Mux.scala 46:16:@11714.4]
  wire  _T_12488; // @[Mux.scala 46:19:@11715.4]
  wire [7:0] _T_12489; // @[Mux.scala 46:16:@11716.4]
  wire  _T_12490; // @[Mux.scala 46:19:@11717.4]
  wire [7:0] _T_12491; // @[Mux.scala 46:16:@11718.4]
  wire  _T_12492; // @[Mux.scala 46:19:@11719.4]
  wire [7:0] _T_12493; // @[Mux.scala 46:16:@11720.4]
  wire  _T_12494; // @[Mux.scala 46:19:@11721.4]
  wire [7:0] _T_12495; // @[Mux.scala 46:16:@11722.4]
  wire  _T_12496; // @[Mux.scala 46:19:@11723.4]
  wire [7:0] _T_12497; // @[Mux.scala 46:16:@11724.4]
  wire  _T_12498; // @[Mux.scala 46:19:@11725.4]
  wire [7:0] _T_12499; // @[Mux.scala 46:16:@11726.4]
  wire  _T_12500; // @[Mux.scala 46:19:@11727.4]
  wire [7:0] _T_12501; // @[Mux.scala 46:16:@11728.4]
  wire  _T_12502; // @[Mux.scala 46:19:@11729.4]
  wire [7:0] _T_12503; // @[Mux.scala 46:16:@11730.4]
  wire  _T_12504; // @[Mux.scala 46:19:@11731.4]
  wire [7:0] _T_12505; // @[Mux.scala 46:16:@11732.4]
  wire  _T_12506; // @[Mux.scala 46:19:@11733.4]
  wire [7:0] _T_12507; // @[Mux.scala 46:16:@11734.4]
  wire  _T_12508; // @[Mux.scala 46:19:@11735.4]
  wire [7:0] _T_12509; // @[Mux.scala 46:16:@11736.4]
  wire  _T_12510; // @[Mux.scala 46:19:@11737.4]
  wire [7:0] _T_12511; // @[Mux.scala 46:16:@11738.4]
  wire  _T_12512; // @[Mux.scala 46:19:@11739.4]
  wire [7:0] _T_12513; // @[Mux.scala 46:16:@11740.4]
  wire  _T_12514; // @[Mux.scala 46:19:@11741.4]
  wire [7:0] _T_12515; // @[Mux.scala 46:16:@11742.4]
  wire  _T_12543; // @[Mux.scala 46:19:@11744.4]
  wire [7:0] _T_12544; // @[Mux.scala 46:16:@11745.4]
  wire  _T_12545; // @[Mux.scala 46:19:@11746.4]
  wire [7:0] _T_12546; // @[Mux.scala 46:16:@11747.4]
  wire  _T_12547; // @[Mux.scala 46:19:@11748.4]
  wire [7:0] _T_12548; // @[Mux.scala 46:16:@11749.4]
  wire  _T_12549; // @[Mux.scala 46:19:@11750.4]
  wire [7:0] _T_12550; // @[Mux.scala 46:16:@11751.4]
  wire  _T_12551; // @[Mux.scala 46:19:@11752.4]
  wire [7:0] _T_12552; // @[Mux.scala 46:16:@11753.4]
  wire  _T_12553; // @[Mux.scala 46:19:@11754.4]
  wire [7:0] _T_12554; // @[Mux.scala 46:16:@11755.4]
  wire  _T_12555; // @[Mux.scala 46:19:@11756.4]
  wire [7:0] _T_12556; // @[Mux.scala 46:16:@11757.4]
  wire  _T_12557; // @[Mux.scala 46:19:@11758.4]
  wire [7:0] _T_12558; // @[Mux.scala 46:16:@11759.4]
  wire  _T_12559; // @[Mux.scala 46:19:@11760.4]
  wire [7:0] _T_12560; // @[Mux.scala 46:16:@11761.4]
  wire  _T_12561; // @[Mux.scala 46:19:@11762.4]
  wire [7:0] _T_12562; // @[Mux.scala 46:16:@11763.4]
  wire  _T_12563; // @[Mux.scala 46:19:@11764.4]
  wire [7:0] _T_12564; // @[Mux.scala 46:16:@11765.4]
  wire  _T_12565; // @[Mux.scala 46:19:@11766.4]
  wire [7:0] _T_12566; // @[Mux.scala 46:16:@11767.4]
  wire  _T_12567; // @[Mux.scala 46:19:@11768.4]
  wire [7:0] _T_12568; // @[Mux.scala 46:16:@11769.4]
  wire  _T_12569; // @[Mux.scala 46:19:@11770.4]
  wire [7:0] _T_12570; // @[Mux.scala 46:16:@11771.4]
  wire  _T_12571; // @[Mux.scala 46:19:@11772.4]
  wire [7:0] _T_12572; // @[Mux.scala 46:16:@11773.4]
  wire  _T_12573; // @[Mux.scala 46:19:@11774.4]
  wire [7:0] _T_12574; // @[Mux.scala 46:16:@11775.4]
  wire  _T_12575; // @[Mux.scala 46:19:@11776.4]
  wire [7:0] _T_12576; // @[Mux.scala 46:16:@11777.4]
  wire  _T_12577; // @[Mux.scala 46:19:@11778.4]
  wire [7:0] _T_12578; // @[Mux.scala 46:16:@11779.4]
  wire  _T_12579; // @[Mux.scala 46:19:@11780.4]
  wire [7:0] _T_12580; // @[Mux.scala 46:16:@11781.4]
  wire  _T_12581; // @[Mux.scala 46:19:@11782.4]
  wire [7:0] _T_12582; // @[Mux.scala 46:16:@11783.4]
  wire  _T_12583; // @[Mux.scala 46:19:@11784.4]
  wire [7:0] _T_12584; // @[Mux.scala 46:16:@11785.4]
  wire  _T_12585; // @[Mux.scala 46:19:@11786.4]
  wire [7:0] _T_12586; // @[Mux.scala 46:16:@11787.4]
  wire  _T_12587; // @[Mux.scala 46:19:@11788.4]
  wire [7:0] _T_12588; // @[Mux.scala 46:16:@11789.4]
  wire  _T_12589; // @[Mux.scala 46:19:@11790.4]
  wire [7:0] _T_12590; // @[Mux.scala 46:16:@11791.4]
  wire  _T_12591; // @[Mux.scala 46:19:@11792.4]
  wire [7:0] _T_12592; // @[Mux.scala 46:16:@11793.4]
  wire  _T_12593; // @[Mux.scala 46:19:@11794.4]
  wire [7:0] _T_12594; // @[Mux.scala 46:16:@11795.4]
  wire  _T_12623; // @[Mux.scala 46:19:@11797.4]
  wire [7:0] _T_12624; // @[Mux.scala 46:16:@11798.4]
  wire  _T_12625; // @[Mux.scala 46:19:@11799.4]
  wire [7:0] _T_12626; // @[Mux.scala 46:16:@11800.4]
  wire  _T_12627; // @[Mux.scala 46:19:@11801.4]
  wire [7:0] _T_12628; // @[Mux.scala 46:16:@11802.4]
  wire  _T_12629; // @[Mux.scala 46:19:@11803.4]
  wire [7:0] _T_12630; // @[Mux.scala 46:16:@11804.4]
  wire  _T_12631; // @[Mux.scala 46:19:@11805.4]
  wire [7:0] _T_12632; // @[Mux.scala 46:16:@11806.4]
  wire  _T_12633; // @[Mux.scala 46:19:@11807.4]
  wire [7:0] _T_12634; // @[Mux.scala 46:16:@11808.4]
  wire  _T_12635; // @[Mux.scala 46:19:@11809.4]
  wire [7:0] _T_12636; // @[Mux.scala 46:16:@11810.4]
  wire  _T_12637; // @[Mux.scala 46:19:@11811.4]
  wire [7:0] _T_12638; // @[Mux.scala 46:16:@11812.4]
  wire  _T_12639; // @[Mux.scala 46:19:@11813.4]
  wire [7:0] _T_12640; // @[Mux.scala 46:16:@11814.4]
  wire  _T_12641; // @[Mux.scala 46:19:@11815.4]
  wire [7:0] _T_12642; // @[Mux.scala 46:16:@11816.4]
  wire  _T_12643; // @[Mux.scala 46:19:@11817.4]
  wire [7:0] _T_12644; // @[Mux.scala 46:16:@11818.4]
  wire  _T_12645; // @[Mux.scala 46:19:@11819.4]
  wire [7:0] _T_12646; // @[Mux.scala 46:16:@11820.4]
  wire  _T_12647; // @[Mux.scala 46:19:@11821.4]
  wire [7:0] _T_12648; // @[Mux.scala 46:16:@11822.4]
  wire  _T_12649; // @[Mux.scala 46:19:@11823.4]
  wire [7:0] _T_12650; // @[Mux.scala 46:16:@11824.4]
  wire  _T_12651; // @[Mux.scala 46:19:@11825.4]
  wire [7:0] _T_12652; // @[Mux.scala 46:16:@11826.4]
  wire  _T_12653; // @[Mux.scala 46:19:@11827.4]
  wire [7:0] _T_12654; // @[Mux.scala 46:16:@11828.4]
  wire  _T_12655; // @[Mux.scala 46:19:@11829.4]
  wire [7:0] _T_12656; // @[Mux.scala 46:16:@11830.4]
  wire  _T_12657; // @[Mux.scala 46:19:@11831.4]
  wire [7:0] _T_12658; // @[Mux.scala 46:16:@11832.4]
  wire  _T_12659; // @[Mux.scala 46:19:@11833.4]
  wire [7:0] _T_12660; // @[Mux.scala 46:16:@11834.4]
  wire  _T_12661; // @[Mux.scala 46:19:@11835.4]
  wire [7:0] _T_12662; // @[Mux.scala 46:16:@11836.4]
  wire  _T_12663; // @[Mux.scala 46:19:@11837.4]
  wire [7:0] _T_12664; // @[Mux.scala 46:16:@11838.4]
  wire  _T_12665; // @[Mux.scala 46:19:@11839.4]
  wire [7:0] _T_12666; // @[Mux.scala 46:16:@11840.4]
  wire  _T_12667; // @[Mux.scala 46:19:@11841.4]
  wire [7:0] _T_12668; // @[Mux.scala 46:16:@11842.4]
  wire  _T_12669; // @[Mux.scala 46:19:@11843.4]
  wire [7:0] _T_12670; // @[Mux.scala 46:16:@11844.4]
  wire  _T_12671; // @[Mux.scala 46:19:@11845.4]
  wire [7:0] _T_12672; // @[Mux.scala 46:16:@11846.4]
  wire  _T_12673; // @[Mux.scala 46:19:@11847.4]
  wire [7:0] _T_12674; // @[Mux.scala 46:16:@11848.4]
  wire  _T_12675; // @[Mux.scala 46:19:@11849.4]
  wire [7:0] _T_12676; // @[Mux.scala 46:16:@11850.4]
  wire  _T_12706; // @[Mux.scala 46:19:@11852.4]
  wire [7:0] _T_12707; // @[Mux.scala 46:16:@11853.4]
  wire  _T_12708; // @[Mux.scala 46:19:@11854.4]
  wire [7:0] _T_12709; // @[Mux.scala 46:16:@11855.4]
  wire  _T_12710; // @[Mux.scala 46:19:@11856.4]
  wire [7:0] _T_12711; // @[Mux.scala 46:16:@11857.4]
  wire  _T_12712; // @[Mux.scala 46:19:@11858.4]
  wire [7:0] _T_12713; // @[Mux.scala 46:16:@11859.4]
  wire  _T_12714; // @[Mux.scala 46:19:@11860.4]
  wire [7:0] _T_12715; // @[Mux.scala 46:16:@11861.4]
  wire  _T_12716; // @[Mux.scala 46:19:@11862.4]
  wire [7:0] _T_12717; // @[Mux.scala 46:16:@11863.4]
  wire  _T_12718; // @[Mux.scala 46:19:@11864.4]
  wire [7:0] _T_12719; // @[Mux.scala 46:16:@11865.4]
  wire  _T_12720; // @[Mux.scala 46:19:@11866.4]
  wire [7:0] _T_12721; // @[Mux.scala 46:16:@11867.4]
  wire  _T_12722; // @[Mux.scala 46:19:@11868.4]
  wire [7:0] _T_12723; // @[Mux.scala 46:16:@11869.4]
  wire  _T_12724; // @[Mux.scala 46:19:@11870.4]
  wire [7:0] _T_12725; // @[Mux.scala 46:16:@11871.4]
  wire  _T_12726; // @[Mux.scala 46:19:@11872.4]
  wire [7:0] _T_12727; // @[Mux.scala 46:16:@11873.4]
  wire  _T_12728; // @[Mux.scala 46:19:@11874.4]
  wire [7:0] _T_12729; // @[Mux.scala 46:16:@11875.4]
  wire  _T_12730; // @[Mux.scala 46:19:@11876.4]
  wire [7:0] _T_12731; // @[Mux.scala 46:16:@11877.4]
  wire  _T_12732; // @[Mux.scala 46:19:@11878.4]
  wire [7:0] _T_12733; // @[Mux.scala 46:16:@11879.4]
  wire  _T_12734; // @[Mux.scala 46:19:@11880.4]
  wire [7:0] _T_12735; // @[Mux.scala 46:16:@11881.4]
  wire  _T_12736; // @[Mux.scala 46:19:@11882.4]
  wire [7:0] _T_12737; // @[Mux.scala 46:16:@11883.4]
  wire  _T_12738; // @[Mux.scala 46:19:@11884.4]
  wire [7:0] _T_12739; // @[Mux.scala 46:16:@11885.4]
  wire  _T_12740; // @[Mux.scala 46:19:@11886.4]
  wire [7:0] _T_12741; // @[Mux.scala 46:16:@11887.4]
  wire  _T_12742; // @[Mux.scala 46:19:@11888.4]
  wire [7:0] _T_12743; // @[Mux.scala 46:16:@11889.4]
  wire  _T_12744; // @[Mux.scala 46:19:@11890.4]
  wire [7:0] _T_12745; // @[Mux.scala 46:16:@11891.4]
  wire  _T_12746; // @[Mux.scala 46:19:@11892.4]
  wire [7:0] _T_12747; // @[Mux.scala 46:16:@11893.4]
  wire  _T_12748; // @[Mux.scala 46:19:@11894.4]
  wire [7:0] _T_12749; // @[Mux.scala 46:16:@11895.4]
  wire  _T_12750; // @[Mux.scala 46:19:@11896.4]
  wire [7:0] _T_12751; // @[Mux.scala 46:16:@11897.4]
  wire  _T_12752; // @[Mux.scala 46:19:@11898.4]
  wire [7:0] _T_12753; // @[Mux.scala 46:16:@11899.4]
  wire  _T_12754; // @[Mux.scala 46:19:@11900.4]
  wire [7:0] _T_12755; // @[Mux.scala 46:16:@11901.4]
  wire  _T_12756; // @[Mux.scala 46:19:@11902.4]
  wire [7:0] _T_12757; // @[Mux.scala 46:16:@11903.4]
  wire  _T_12758; // @[Mux.scala 46:19:@11904.4]
  wire [7:0] _T_12759; // @[Mux.scala 46:16:@11905.4]
  wire  _T_12760; // @[Mux.scala 46:19:@11906.4]
  wire [7:0] _T_12761; // @[Mux.scala 46:16:@11907.4]
  wire  _T_12792; // @[Mux.scala 46:19:@11909.4]
  wire [7:0] _T_12793; // @[Mux.scala 46:16:@11910.4]
  wire  _T_12794; // @[Mux.scala 46:19:@11911.4]
  wire [7:0] _T_12795; // @[Mux.scala 46:16:@11912.4]
  wire  _T_12796; // @[Mux.scala 46:19:@11913.4]
  wire [7:0] _T_12797; // @[Mux.scala 46:16:@11914.4]
  wire  _T_12798; // @[Mux.scala 46:19:@11915.4]
  wire [7:0] _T_12799; // @[Mux.scala 46:16:@11916.4]
  wire  _T_12800; // @[Mux.scala 46:19:@11917.4]
  wire [7:0] _T_12801; // @[Mux.scala 46:16:@11918.4]
  wire  _T_12802; // @[Mux.scala 46:19:@11919.4]
  wire [7:0] _T_12803; // @[Mux.scala 46:16:@11920.4]
  wire  _T_12804; // @[Mux.scala 46:19:@11921.4]
  wire [7:0] _T_12805; // @[Mux.scala 46:16:@11922.4]
  wire  _T_12806; // @[Mux.scala 46:19:@11923.4]
  wire [7:0] _T_12807; // @[Mux.scala 46:16:@11924.4]
  wire  _T_12808; // @[Mux.scala 46:19:@11925.4]
  wire [7:0] _T_12809; // @[Mux.scala 46:16:@11926.4]
  wire  _T_12810; // @[Mux.scala 46:19:@11927.4]
  wire [7:0] _T_12811; // @[Mux.scala 46:16:@11928.4]
  wire  _T_12812; // @[Mux.scala 46:19:@11929.4]
  wire [7:0] _T_12813; // @[Mux.scala 46:16:@11930.4]
  wire  _T_12814; // @[Mux.scala 46:19:@11931.4]
  wire [7:0] _T_12815; // @[Mux.scala 46:16:@11932.4]
  wire  _T_12816; // @[Mux.scala 46:19:@11933.4]
  wire [7:0] _T_12817; // @[Mux.scala 46:16:@11934.4]
  wire  _T_12818; // @[Mux.scala 46:19:@11935.4]
  wire [7:0] _T_12819; // @[Mux.scala 46:16:@11936.4]
  wire  _T_12820; // @[Mux.scala 46:19:@11937.4]
  wire [7:0] _T_12821; // @[Mux.scala 46:16:@11938.4]
  wire  _T_12822; // @[Mux.scala 46:19:@11939.4]
  wire [7:0] _T_12823; // @[Mux.scala 46:16:@11940.4]
  wire  _T_12824; // @[Mux.scala 46:19:@11941.4]
  wire [7:0] _T_12825; // @[Mux.scala 46:16:@11942.4]
  wire  _T_12826; // @[Mux.scala 46:19:@11943.4]
  wire [7:0] _T_12827; // @[Mux.scala 46:16:@11944.4]
  wire  _T_12828; // @[Mux.scala 46:19:@11945.4]
  wire [7:0] _T_12829; // @[Mux.scala 46:16:@11946.4]
  wire  _T_12830; // @[Mux.scala 46:19:@11947.4]
  wire [7:0] _T_12831; // @[Mux.scala 46:16:@11948.4]
  wire  _T_12832; // @[Mux.scala 46:19:@11949.4]
  wire [7:0] _T_12833; // @[Mux.scala 46:16:@11950.4]
  wire  _T_12834; // @[Mux.scala 46:19:@11951.4]
  wire [7:0] _T_12835; // @[Mux.scala 46:16:@11952.4]
  wire  _T_12836; // @[Mux.scala 46:19:@11953.4]
  wire [7:0] _T_12837; // @[Mux.scala 46:16:@11954.4]
  wire  _T_12838; // @[Mux.scala 46:19:@11955.4]
  wire [7:0] _T_12839; // @[Mux.scala 46:16:@11956.4]
  wire  _T_12840; // @[Mux.scala 46:19:@11957.4]
  wire [7:0] _T_12841; // @[Mux.scala 46:16:@11958.4]
  wire  _T_12842; // @[Mux.scala 46:19:@11959.4]
  wire [7:0] _T_12843; // @[Mux.scala 46:16:@11960.4]
  wire  _T_12844; // @[Mux.scala 46:19:@11961.4]
  wire [7:0] _T_12845; // @[Mux.scala 46:16:@11962.4]
  wire  _T_12846; // @[Mux.scala 46:19:@11963.4]
  wire [7:0] _T_12847; // @[Mux.scala 46:16:@11964.4]
  wire  _T_12848; // @[Mux.scala 46:19:@11965.4]
  wire [7:0] _T_12849; // @[Mux.scala 46:16:@11966.4]
  wire  _T_12881; // @[Mux.scala 46:19:@11968.4]
  wire [7:0] _T_12882; // @[Mux.scala 46:16:@11969.4]
  wire  _T_12883; // @[Mux.scala 46:19:@11970.4]
  wire [7:0] _T_12884; // @[Mux.scala 46:16:@11971.4]
  wire  _T_12885; // @[Mux.scala 46:19:@11972.4]
  wire [7:0] _T_12886; // @[Mux.scala 46:16:@11973.4]
  wire  _T_12887; // @[Mux.scala 46:19:@11974.4]
  wire [7:0] _T_12888; // @[Mux.scala 46:16:@11975.4]
  wire  _T_12889; // @[Mux.scala 46:19:@11976.4]
  wire [7:0] _T_12890; // @[Mux.scala 46:16:@11977.4]
  wire  _T_12891; // @[Mux.scala 46:19:@11978.4]
  wire [7:0] _T_12892; // @[Mux.scala 46:16:@11979.4]
  wire  _T_12893; // @[Mux.scala 46:19:@11980.4]
  wire [7:0] _T_12894; // @[Mux.scala 46:16:@11981.4]
  wire  _T_12895; // @[Mux.scala 46:19:@11982.4]
  wire [7:0] _T_12896; // @[Mux.scala 46:16:@11983.4]
  wire  _T_12897; // @[Mux.scala 46:19:@11984.4]
  wire [7:0] _T_12898; // @[Mux.scala 46:16:@11985.4]
  wire  _T_12899; // @[Mux.scala 46:19:@11986.4]
  wire [7:0] _T_12900; // @[Mux.scala 46:16:@11987.4]
  wire  _T_12901; // @[Mux.scala 46:19:@11988.4]
  wire [7:0] _T_12902; // @[Mux.scala 46:16:@11989.4]
  wire  _T_12903; // @[Mux.scala 46:19:@11990.4]
  wire [7:0] _T_12904; // @[Mux.scala 46:16:@11991.4]
  wire  _T_12905; // @[Mux.scala 46:19:@11992.4]
  wire [7:0] _T_12906; // @[Mux.scala 46:16:@11993.4]
  wire  _T_12907; // @[Mux.scala 46:19:@11994.4]
  wire [7:0] _T_12908; // @[Mux.scala 46:16:@11995.4]
  wire  _T_12909; // @[Mux.scala 46:19:@11996.4]
  wire [7:0] _T_12910; // @[Mux.scala 46:16:@11997.4]
  wire  _T_12911; // @[Mux.scala 46:19:@11998.4]
  wire [7:0] _T_12912; // @[Mux.scala 46:16:@11999.4]
  wire  _T_12913; // @[Mux.scala 46:19:@12000.4]
  wire [7:0] _T_12914; // @[Mux.scala 46:16:@12001.4]
  wire  _T_12915; // @[Mux.scala 46:19:@12002.4]
  wire [7:0] _T_12916; // @[Mux.scala 46:16:@12003.4]
  wire  _T_12917; // @[Mux.scala 46:19:@12004.4]
  wire [7:0] _T_12918; // @[Mux.scala 46:16:@12005.4]
  wire  _T_12919; // @[Mux.scala 46:19:@12006.4]
  wire [7:0] _T_12920; // @[Mux.scala 46:16:@12007.4]
  wire  _T_12921; // @[Mux.scala 46:19:@12008.4]
  wire [7:0] _T_12922; // @[Mux.scala 46:16:@12009.4]
  wire  _T_12923; // @[Mux.scala 46:19:@12010.4]
  wire [7:0] _T_12924; // @[Mux.scala 46:16:@12011.4]
  wire  _T_12925; // @[Mux.scala 46:19:@12012.4]
  wire [7:0] _T_12926; // @[Mux.scala 46:16:@12013.4]
  wire  _T_12927; // @[Mux.scala 46:19:@12014.4]
  wire [7:0] _T_12928; // @[Mux.scala 46:16:@12015.4]
  wire  _T_12929; // @[Mux.scala 46:19:@12016.4]
  wire [7:0] _T_12930; // @[Mux.scala 46:16:@12017.4]
  wire  _T_12931; // @[Mux.scala 46:19:@12018.4]
  wire [7:0] _T_12932; // @[Mux.scala 46:16:@12019.4]
  wire  _T_12933; // @[Mux.scala 46:19:@12020.4]
  wire [7:0] _T_12934; // @[Mux.scala 46:16:@12021.4]
  wire  _T_12935; // @[Mux.scala 46:19:@12022.4]
  wire [7:0] _T_12936; // @[Mux.scala 46:16:@12023.4]
  wire  _T_12937; // @[Mux.scala 46:19:@12024.4]
  wire [7:0] _T_12938; // @[Mux.scala 46:16:@12025.4]
  wire  _T_12939; // @[Mux.scala 46:19:@12026.4]
  wire [7:0] _T_12940; // @[Mux.scala 46:16:@12027.4]
  wire  _T_12973; // @[Mux.scala 46:19:@12029.4]
  wire [7:0] _T_12974; // @[Mux.scala 46:16:@12030.4]
  wire  _T_12975; // @[Mux.scala 46:19:@12031.4]
  wire [7:0] _T_12976; // @[Mux.scala 46:16:@12032.4]
  wire  _T_12977; // @[Mux.scala 46:19:@12033.4]
  wire [7:0] _T_12978; // @[Mux.scala 46:16:@12034.4]
  wire  _T_12979; // @[Mux.scala 46:19:@12035.4]
  wire [7:0] _T_12980; // @[Mux.scala 46:16:@12036.4]
  wire  _T_12981; // @[Mux.scala 46:19:@12037.4]
  wire [7:0] _T_12982; // @[Mux.scala 46:16:@12038.4]
  wire  _T_12983; // @[Mux.scala 46:19:@12039.4]
  wire [7:0] _T_12984; // @[Mux.scala 46:16:@12040.4]
  wire  _T_12985; // @[Mux.scala 46:19:@12041.4]
  wire [7:0] _T_12986; // @[Mux.scala 46:16:@12042.4]
  wire  _T_12987; // @[Mux.scala 46:19:@12043.4]
  wire [7:0] _T_12988; // @[Mux.scala 46:16:@12044.4]
  wire  _T_12989; // @[Mux.scala 46:19:@12045.4]
  wire [7:0] _T_12990; // @[Mux.scala 46:16:@12046.4]
  wire  _T_12991; // @[Mux.scala 46:19:@12047.4]
  wire [7:0] _T_12992; // @[Mux.scala 46:16:@12048.4]
  wire  _T_12993; // @[Mux.scala 46:19:@12049.4]
  wire [7:0] _T_12994; // @[Mux.scala 46:16:@12050.4]
  wire  _T_12995; // @[Mux.scala 46:19:@12051.4]
  wire [7:0] _T_12996; // @[Mux.scala 46:16:@12052.4]
  wire  _T_12997; // @[Mux.scala 46:19:@12053.4]
  wire [7:0] _T_12998; // @[Mux.scala 46:16:@12054.4]
  wire  _T_12999; // @[Mux.scala 46:19:@12055.4]
  wire [7:0] _T_13000; // @[Mux.scala 46:16:@12056.4]
  wire  _T_13001; // @[Mux.scala 46:19:@12057.4]
  wire [7:0] _T_13002; // @[Mux.scala 46:16:@12058.4]
  wire  _T_13003; // @[Mux.scala 46:19:@12059.4]
  wire [7:0] _T_13004; // @[Mux.scala 46:16:@12060.4]
  wire  _T_13005; // @[Mux.scala 46:19:@12061.4]
  wire [7:0] _T_13006; // @[Mux.scala 46:16:@12062.4]
  wire  _T_13007; // @[Mux.scala 46:19:@12063.4]
  wire [7:0] _T_13008; // @[Mux.scala 46:16:@12064.4]
  wire  _T_13009; // @[Mux.scala 46:19:@12065.4]
  wire [7:0] _T_13010; // @[Mux.scala 46:16:@12066.4]
  wire  _T_13011; // @[Mux.scala 46:19:@12067.4]
  wire [7:0] _T_13012; // @[Mux.scala 46:16:@12068.4]
  wire  _T_13013; // @[Mux.scala 46:19:@12069.4]
  wire [7:0] _T_13014; // @[Mux.scala 46:16:@12070.4]
  wire  _T_13015; // @[Mux.scala 46:19:@12071.4]
  wire [7:0] _T_13016; // @[Mux.scala 46:16:@12072.4]
  wire  _T_13017; // @[Mux.scala 46:19:@12073.4]
  wire [7:0] _T_13018; // @[Mux.scala 46:16:@12074.4]
  wire  _T_13019; // @[Mux.scala 46:19:@12075.4]
  wire [7:0] _T_13020; // @[Mux.scala 46:16:@12076.4]
  wire  _T_13021; // @[Mux.scala 46:19:@12077.4]
  wire [7:0] _T_13022; // @[Mux.scala 46:16:@12078.4]
  wire  _T_13023; // @[Mux.scala 46:19:@12079.4]
  wire [7:0] _T_13024; // @[Mux.scala 46:16:@12080.4]
  wire  _T_13025; // @[Mux.scala 46:19:@12081.4]
  wire [7:0] _T_13026; // @[Mux.scala 46:16:@12082.4]
  wire  _T_13027; // @[Mux.scala 46:19:@12083.4]
  wire [7:0] _T_13028; // @[Mux.scala 46:16:@12084.4]
  wire  _T_13029; // @[Mux.scala 46:19:@12085.4]
  wire [7:0] _T_13030; // @[Mux.scala 46:16:@12086.4]
  wire  _T_13031; // @[Mux.scala 46:19:@12087.4]
  wire [7:0] _T_13032; // @[Mux.scala 46:16:@12088.4]
  wire  _T_13033; // @[Mux.scala 46:19:@12089.4]
  wire [7:0] _T_13034; // @[Mux.scala 46:16:@12090.4]
  wire  _T_13068; // @[Mux.scala 46:19:@12092.4]
  wire [7:0] _T_13069; // @[Mux.scala 46:16:@12093.4]
  wire  _T_13070; // @[Mux.scala 46:19:@12094.4]
  wire [7:0] _T_13071; // @[Mux.scala 46:16:@12095.4]
  wire  _T_13072; // @[Mux.scala 46:19:@12096.4]
  wire [7:0] _T_13073; // @[Mux.scala 46:16:@12097.4]
  wire  _T_13074; // @[Mux.scala 46:19:@12098.4]
  wire [7:0] _T_13075; // @[Mux.scala 46:16:@12099.4]
  wire  _T_13076; // @[Mux.scala 46:19:@12100.4]
  wire [7:0] _T_13077; // @[Mux.scala 46:16:@12101.4]
  wire  _T_13078; // @[Mux.scala 46:19:@12102.4]
  wire [7:0] _T_13079; // @[Mux.scala 46:16:@12103.4]
  wire  _T_13080; // @[Mux.scala 46:19:@12104.4]
  wire [7:0] _T_13081; // @[Mux.scala 46:16:@12105.4]
  wire  _T_13082; // @[Mux.scala 46:19:@12106.4]
  wire [7:0] _T_13083; // @[Mux.scala 46:16:@12107.4]
  wire  _T_13084; // @[Mux.scala 46:19:@12108.4]
  wire [7:0] _T_13085; // @[Mux.scala 46:16:@12109.4]
  wire  _T_13086; // @[Mux.scala 46:19:@12110.4]
  wire [7:0] _T_13087; // @[Mux.scala 46:16:@12111.4]
  wire  _T_13088; // @[Mux.scala 46:19:@12112.4]
  wire [7:0] _T_13089; // @[Mux.scala 46:16:@12113.4]
  wire  _T_13090; // @[Mux.scala 46:19:@12114.4]
  wire [7:0] _T_13091; // @[Mux.scala 46:16:@12115.4]
  wire  _T_13092; // @[Mux.scala 46:19:@12116.4]
  wire [7:0] _T_13093; // @[Mux.scala 46:16:@12117.4]
  wire  _T_13094; // @[Mux.scala 46:19:@12118.4]
  wire [7:0] _T_13095; // @[Mux.scala 46:16:@12119.4]
  wire  _T_13096; // @[Mux.scala 46:19:@12120.4]
  wire [7:0] _T_13097; // @[Mux.scala 46:16:@12121.4]
  wire  _T_13098; // @[Mux.scala 46:19:@12122.4]
  wire [7:0] _T_13099; // @[Mux.scala 46:16:@12123.4]
  wire  _T_13100; // @[Mux.scala 46:19:@12124.4]
  wire [7:0] _T_13101; // @[Mux.scala 46:16:@12125.4]
  wire  _T_13102; // @[Mux.scala 46:19:@12126.4]
  wire [7:0] _T_13103; // @[Mux.scala 46:16:@12127.4]
  wire  _T_13104; // @[Mux.scala 46:19:@12128.4]
  wire [7:0] _T_13105; // @[Mux.scala 46:16:@12129.4]
  wire  _T_13106; // @[Mux.scala 46:19:@12130.4]
  wire [7:0] _T_13107; // @[Mux.scala 46:16:@12131.4]
  wire  _T_13108; // @[Mux.scala 46:19:@12132.4]
  wire [7:0] _T_13109; // @[Mux.scala 46:16:@12133.4]
  wire  _T_13110; // @[Mux.scala 46:19:@12134.4]
  wire [7:0] _T_13111; // @[Mux.scala 46:16:@12135.4]
  wire  _T_13112; // @[Mux.scala 46:19:@12136.4]
  wire [7:0] _T_13113; // @[Mux.scala 46:16:@12137.4]
  wire  _T_13114; // @[Mux.scala 46:19:@12138.4]
  wire [7:0] _T_13115; // @[Mux.scala 46:16:@12139.4]
  wire  _T_13116; // @[Mux.scala 46:19:@12140.4]
  wire [7:0] _T_13117; // @[Mux.scala 46:16:@12141.4]
  wire  _T_13118; // @[Mux.scala 46:19:@12142.4]
  wire [7:0] _T_13119; // @[Mux.scala 46:16:@12143.4]
  wire  _T_13120; // @[Mux.scala 46:19:@12144.4]
  wire [7:0] _T_13121; // @[Mux.scala 46:16:@12145.4]
  wire  _T_13122; // @[Mux.scala 46:19:@12146.4]
  wire [7:0] _T_13123; // @[Mux.scala 46:16:@12147.4]
  wire  _T_13124; // @[Mux.scala 46:19:@12148.4]
  wire [7:0] _T_13125; // @[Mux.scala 46:16:@12149.4]
  wire  _T_13126; // @[Mux.scala 46:19:@12150.4]
  wire [7:0] _T_13127; // @[Mux.scala 46:16:@12151.4]
  wire  _T_13128; // @[Mux.scala 46:19:@12152.4]
  wire [7:0] _T_13129; // @[Mux.scala 46:16:@12153.4]
  wire  _T_13130; // @[Mux.scala 46:19:@12154.4]
  wire [7:0] _T_13131; // @[Mux.scala 46:16:@12155.4]
  wire  _T_13166; // @[Mux.scala 46:19:@12157.4]
  wire [7:0] _T_13167; // @[Mux.scala 46:16:@12158.4]
  wire  _T_13168; // @[Mux.scala 46:19:@12159.4]
  wire [7:0] _T_13169; // @[Mux.scala 46:16:@12160.4]
  wire  _T_13170; // @[Mux.scala 46:19:@12161.4]
  wire [7:0] _T_13171; // @[Mux.scala 46:16:@12162.4]
  wire  _T_13172; // @[Mux.scala 46:19:@12163.4]
  wire [7:0] _T_13173; // @[Mux.scala 46:16:@12164.4]
  wire  _T_13174; // @[Mux.scala 46:19:@12165.4]
  wire [7:0] _T_13175; // @[Mux.scala 46:16:@12166.4]
  wire  _T_13176; // @[Mux.scala 46:19:@12167.4]
  wire [7:0] _T_13177; // @[Mux.scala 46:16:@12168.4]
  wire  _T_13178; // @[Mux.scala 46:19:@12169.4]
  wire [7:0] _T_13179; // @[Mux.scala 46:16:@12170.4]
  wire  _T_13180; // @[Mux.scala 46:19:@12171.4]
  wire [7:0] _T_13181; // @[Mux.scala 46:16:@12172.4]
  wire  _T_13182; // @[Mux.scala 46:19:@12173.4]
  wire [7:0] _T_13183; // @[Mux.scala 46:16:@12174.4]
  wire  _T_13184; // @[Mux.scala 46:19:@12175.4]
  wire [7:0] _T_13185; // @[Mux.scala 46:16:@12176.4]
  wire  _T_13186; // @[Mux.scala 46:19:@12177.4]
  wire [7:0] _T_13187; // @[Mux.scala 46:16:@12178.4]
  wire  _T_13188; // @[Mux.scala 46:19:@12179.4]
  wire [7:0] _T_13189; // @[Mux.scala 46:16:@12180.4]
  wire  _T_13190; // @[Mux.scala 46:19:@12181.4]
  wire [7:0] _T_13191; // @[Mux.scala 46:16:@12182.4]
  wire  _T_13192; // @[Mux.scala 46:19:@12183.4]
  wire [7:0] _T_13193; // @[Mux.scala 46:16:@12184.4]
  wire  _T_13194; // @[Mux.scala 46:19:@12185.4]
  wire [7:0] _T_13195; // @[Mux.scala 46:16:@12186.4]
  wire  _T_13196; // @[Mux.scala 46:19:@12187.4]
  wire [7:0] _T_13197; // @[Mux.scala 46:16:@12188.4]
  wire  _T_13198; // @[Mux.scala 46:19:@12189.4]
  wire [7:0] _T_13199; // @[Mux.scala 46:16:@12190.4]
  wire  _T_13200; // @[Mux.scala 46:19:@12191.4]
  wire [7:0] _T_13201; // @[Mux.scala 46:16:@12192.4]
  wire  _T_13202; // @[Mux.scala 46:19:@12193.4]
  wire [7:0] _T_13203; // @[Mux.scala 46:16:@12194.4]
  wire  _T_13204; // @[Mux.scala 46:19:@12195.4]
  wire [7:0] _T_13205; // @[Mux.scala 46:16:@12196.4]
  wire  _T_13206; // @[Mux.scala 46:19:@12197.4]
  wire [7:0] _T_13207; // @[Mux.scala 46:16:@12198.4]
  wire  _T_13208; // @[Mux.scala 46:19:@12199.4]
  wire [7:0] _T_13209; // @[Mux.scala 46:16:@12200.4]
  wire  _T_13210; // @[Mux.scala 46:19:@12201.4]
  wire [7:0] _T_13211; // @[Mux.scala 46:16:@12202.4]
  wire  _T_13212; // @[Mux.scala 46:19:@12203.4]
  wire [7:0] _T_13213; // @[Mux.scala 46:16:@12204.4]
  wire  _T_13214; // @[Mux.scala 46:19:@12205.4]
  wire [7:0] _T_13215; // @[Mux.scala 46:16:@12206.4]
  wire  _T_13216; // @[Mux.scala 46:19:@12207.4]
  wire [7:0] _T_13217; // @[Mux.scala 46:16:@12208.4]
  wire  _T_13218; // @[Mux.scala 46:19:@12209.4]
  wire [7:0] _T_13219; // @[Mux.scala 46:16:@12210.4]
  wire  _T_13220; // @[Mux.scala 46:19:@12211.4]
  wire [7:0] _T_13221; // @[Mux.scala 46:16:@12212.4]
  wire  _T_13222; // @[Mux.scala 46:19:@12213.4]
  wire [7:0] _T_13223; // @[Mux.scala 46:16:@12214.4]
  wire  _T_13224; // @[Mux.scala 46:19:@12215.4]
  wire [7:0] _T_13225; // @[Mux.scala 46:16:@12216.4]
  wire  _T_13226; // @[Mux.scala 46:19:@12217.4]
  wire [7:0] _T_13227; // @[Mux.scala 46:16:@12218.4]
  wire  _T_13228; // @[Mux.scala 46:19:@12219.4]
  wire [7:0] _T_13229; // @[Mux.scala 46:16:@12220.4]
  wire  _T_13230; // @[Mux.scala 46:19:@12221.4]
  wire [7:0] _T_13231; // @[Mux.scala 46:16:@12222.4]
  wire  _T_13267; // @[Mux.scala 46:19:@12224.4]
  wire [7:0] _T_13268; // @[Mux.scala 46:16:@12225.4]
  wire  _T_13269; // @[Mux.scala 46:19:@12226.4]
  wire [7:0] _T_13270; // @[Mux.scala 46:16:@12227.4]
  wire  _T_13271; // @[Mux.scala 46:19:@12228.4]
  wire [7:0] _T_13272; // @[Mux.scala 46:16:@12229.4]
  wire  _T_13273; // @[Mux.scala 46:19:@12230.4]
  wire [7:0] _T_13274; // @[Mux.scala 46:16:@12231.4]
  wire  _T_13275; // @[Mux.scala 46:19:@12232.4]
  wire [7:0] _T_13276; // @[Mux.scala 46:16:@12233.4]
  wire  _T_13277; // @[Mux.scala 46:19:@12234.4]
  wire [7:0] _T_13278; // @[Mux.scala 46:16:@12235.4]
  wire  _T_13279; // @[Mux.scala 46:19:@12236.4]
  wire [7:0] _T_13280; // @[Mux.scala 46:16:@12237.4]
  wire  _T_13281; // @[Mux.scala 46:19:@12238.4]
  wire [7:0] _T_13282; // @[Mux.scala 46:16:@12239.4]
  wire  _T_13283; // @[Mux.scala 46:19:@12240.4]
  wire [7:0] _T_13284; // @[Mux.scala 46:16:@12241.4]
  wire  _T_13285; // @[Mux.scala 46:19:@12242.4]
  wire [7:0] _T_13286; // @[Mux.scala 46:16:@12243.4]
  wire  _T_13287; // @[Mux.scala 46:19:@12244.4]
  wire [7:0] _T_13288; // @[Mux.scala 46:16:@12245.4]
  wire  _T_13289; // @[Mux.scala 46:19:@12246.4]
  wire [7:0] _T_13290; // @[Mux.scala 46:16:@12247.4]
  wire  _T_13291; // @[Mux.scala 46:19:@12248.4]
  wire [7:0] _T_13292; // @[Mux.scala 46:16:@12249.4]
  wire  _T_13293; // @[Mux.scala 46:19:@12250.4]
  wire [7:0] _T_13294; // @[Mux.scala 46:16:@12251.4]
  wire  _T_13295; // @[Mux.scala 46:19:@12252.4]
  wire [7:0] _T_13296; // @[Mux.scala 46:16:@12253.4]
  wire  _T_13297; // @[Mux.scala 46:19:@12254.4]
  wire [7:0] _T_13298; // @[Mux.scala 46:16:@12255.4]
  wire  _T_13299; // @[Mux.scala 46:19:@12256.4]
  wire [7:0] _T_13300; // @[Mux.scala 46:16:@12257.4]
  wire  _T_13301; // @[Mux.scala 46:19:@12258.4]
  wire [7:0] _T_13302; // @[Mux.scala 46:16:@12259.4]
  wire  _T_13303; // @[Mux.scala 46:19:@12260.4]
  wire [7:0] _T_13304; // @[Mux.scala 46:16:@12261.4]
  wire  _T_13305; // @[Mux.scala 46:19:@12262.4]
  wire [7:0] _T_13306; // @[Mux.scala 46:16:@12263.4]
  wire  _T_13307; // @[Mux.scala 46:19:@12264.4]
  wire [7:0] _T_13308; // @[Mux.scala 46:16:@12265.4]
  wire  _T_13309; // @[Mux.scala 46:19:@12266.4]
  wire [7:0] _T_13310; // @[Mux.scala 46:16:@12267.4]
  wire  _T_13311; // @[Mux.scala 46:19:@12268.4]
  wire [7:0] _T_13312; // @[Mux.scala 46:16:@12269.4]
  wire  _T_13313; // @[Mux.scala 46:19:@12270.4]
  wire [7:0] _T_13314; // @[Mux.scala 46:16:@12271.4]
  wire  _T_13315; // @[Mux.scala 46:19:@12272.4]
  wire [7:0] _T_13316; // @[Mux.scala 46:16:@12273.4]
  wire  _T_13317; // @[Mux.scala 46:19:@12274.4]
  wire [7:0] _T_13318; // @[Mux.scala 46:16:@12275.4]
  wire  _T_13319; // @[Mux.scala 46:19:@12276.4]
  wire [7:0] _T_13320; // @[Mux.scala 46:16:@12277.4]
  wire  _T_13321; // @[Mux.scala 46:19:@12278.4]
  wire [7:0] _T_13322; // @[Mux.scala 46:16:@12279.4]
  wire  _T_13323; // @[Mux.scala 46:19:@12280.4]
  wire [7:0] _T_13324; // @[Mux.scala 46:16:@12281.4]
  wire  _T_13325; // @[Mux.scala 46:19:@12282.4]
  wire [7:0] _T_13326; // @[Mux.scala 46:16:@12283.4]
  wire  _T_13327; // @[Mux.scala 46:19:@12284.4]
  wire [7:0] _T_13328; // @[Mux.scala 46:16:@12285.4]
  wire  _T_13329; // @[Mux.scala 46:19:@12286.4]
  wire [7:0] _T_13330; // @[Mux.scala 46:16:@12287.4]
  wire  _T_13331; // @[Mux.scala 46:19:@12288.4]
  wire [7:0] _T_13332; // @[Mux.scala 46:16:@12289.4]
  wire  _T_13333; // @[Mux.scala 46:19:@12290.4]
  wire [7:0] _T_13334; // @[Mux.scala 46:16:@12291.4]
  wire  _T_13371; // @[Mux.scala 46:19:@12293.4]
  wire [7:0] _T_13372; // @[Mux.scala 46:16:@12294.4]
  wire  _T_13373; // @[Mux.scala 46:19:@12295.4]
  wire [7:0] _T_13374; // @[Mux.scala 46:16:@12296.4]
  wire  _T_13375; // @[Mux.scala 46:19:@12297.4]
  wire [7:0] _T_13376; // @[Mux.scala 46:16:@12298.4]
  wire  _T_13377; // @[Mux.scala 46:19:@12299.4]
  wire [7:0] _T_13378; // @[Mux.scala 46:16:@12300.4]
  wire  _T_13379; // @[Mux.scala 46:19:@12301.4]
  wire [7:0] _T_13380; // @[Mux.scala 46:16:@12302.4]
  wire  _T_13381; // @[Mux.scala 46:19:@12303.4]
  wire [7:0] _T_13382; // @[Mux.scala 46:16:@12304.4]
  wire  _T_13383; // @[Mux.scala 46:19:@12305.4]
  wire [7:0] _T_13384; // @[Mux.scala 46:16:@12306.4]
  wire  _T_13385; // @[Mux.scala 46:19:@12307.4]
  wire [7:0] _T_13386; // @[Mux.scala 46:16:@12308.4]
  wire  _T_13387; // @[Mux.scala 46:19:@12309.4]
  wire [7:0] _T_13388; // @[Mux.scala 46:16:@12310.4]
  wire  _T_13389; // @[Mux.scala 46:19:@12311.4]
  wire [7:0] _T_13390; // @[Mux.scala 46:16:@12312.4]
  wire  _T_13391; // @[Mux.scala 46:19:@12313.4]
  wire [7:0] _T_13392; // @[Mux.scala 46:16:@12314.4]
  wire  _T_13393; // @[Mux.scala 46:19:@12315.4]
  wire [7:0] _T_13394; // @[Mux.scala 46:16:@12316.4]
  wire  _T_13395; // @[Mux.scala 46:19:@12317.4]
  wire [7:0] _T_13396; // @[Mux.scala 46:16:@12318.4]
  wire  _T_13397; // @[Mux.scala 46:19:@12319.4]
  wire [7:0] _T_13398; // @[Mux.scala 46:16:@12320.4]
  wire  _T_13399; // @[Mux.scala 46:19:@12321.4]
  wire [7:0] _T_13400; // @[Mux.scala 46:16:@12322.4]
  wire  _T_13401; // @[Mux.scala 46:19:@12323.4]
  wire [7:0] _T_13402; // @[Mux.scala 46:16:@12324.4]
  wire  _T_13403; // @[Mux.scala 46:19:@12325.4]
  wire [7:0] _T_13404; // @[Mux.scala 46:16:@12326.4]
  wire  _T_13405; // @[Mux.scala 46:19:@12327.4]
  wire [7:0] _T_13406; // @[Mux.scala 46:16:@12328.4]
  wire  _T_13407; // @[Mux.scala 46:19:@12329.4]
  wire [7:0] _T_13408; // @[Mux.scala 46:16:@12330.4]
  wire  _T_13409; // @[Mux.scala 46:19:@12331.4]
  wire [7:0] _T_13410; // @[Mux.scala 46:16:@12332.4]
  wire  _T_13411; // @[Mux.scala 46:19:@12333.4]
  wire [7:0] _T_13412; // @[Mux.scala 46:16:@12334.4]
  wire  _T_13413; // @[Mux.scala 46:19:@12335.4]
  wire [7:0] _T_13414; // @[Mux.scala 46:16:@12336.4]
  wire  _T_13415; // @[Mux.scala 46:19:@12337.4]
  wire [7:0] _T_13416; // @[Mux.scala 46:16:@12338.4]
  wire  _T_13417; // @[Mux.scala 46:19:@12339.4]
  wire [7:0] _T_13418; // @[Mux.scala 46:16:@12340.4]
  wire  _T_13419; // @[Mux.scala 46:19:@12341.4]
  wire [7:0] _T_13420; // @[Mux.scala 46:16:@12342.4]
  wire  _T_13421; // @[Mux.scala 46:19:@12343.4]
  wire [7:0] _T_13422; // @[Mux.scala 46:16:@12344.4]
  wire  _T_13423; // @[Mux.scala 46:19:@12345.4]
  wire [7:0] _T_13424; // @[Mux.scala 46:16:@12346.4]
  wire  _T_13425; // @[Mux.scala 46:19:@12347.4]
  wire [7:0] _T_13426; // @[Mux.scala 46:16:@12348.4]
  wire  _T_13427; // @[Mux.scala 46:19:@12349.4]
  wire [7:0] _T_13428; // @[Mux.scala 46:16:@12350.4]
  wire  _T_13429; // @[Mux.scala 46:19:@12351.4]
  wire [7:0] _T_13430; // @[Mux.scala 46:16:@12352.4]
  wire  _T_13431; // @[Mux.scala 46:19:@12353.4]
  wire [7:0] _T_13432; // @[Mux.scala 46:16:@12354.4]
  wire  _T_13433; // @[Mux.scala 46:19:@12355.4]
  wire [7:0] _T_13434; // @[Mux.scala 46:16:@12356.4]
  wire  _T_13435; // @[Mux.scala 46:19:@12357.4]
  wire [7:0] _T_13436; // @[Mux.scala 46:16:@12358.4]
  wire  _T_13437; // @[Mux.scala 46:19:@12359.4]
  wire [7:0] _T_13438; // @[Mux.scala 46:16:@12360.4]
  wire  _T_13439; // @[Mux.scala 46:19:@12361.4]
  wire [7:0] _T_13440; // @[Mux.scala 46:16:@12362.4]
  wire  _T_13478; // @[Mux.scala 46:19:@12364.4]
  wire [7:0] _T_13479; // @[Mux.scala 46:16:@12365.4]
  wire  _T_13480; // @[Mux.scala 46:19:@12366.4]
  wire [7:0] _T_13481; // @[Mux.scala 46:16:@12367.4]
  wire  _T_13482; // @[Mux.scala 46:19:@12368.4]
  wire [7:0] _T_13483; // @[Mux.scala 46:16:@12369.4]
  wire  _T_13484; // @[Mux.scala 46:19:@12370.4]
  wire [7:0] _T_13485; // @[Mux.scala 46:16:@12371.4]
  wire  _T_13486; // @[Mux.scala 46:19:@12372.4]
  wire [7:0] _T_13487; // @[Mux.scala 46:16:@12373.4]
  wire  _T_13488; // @[Mux.scala 46:19:@12374.4]
  wire [7:0] _T_13489; // @[Mux.scala 46:16:@12375.4]
  wire  _T_13490; // @[Mux.scala 46:19:@12376.4]
  wire [7:0] _T_13491; // @[Mux.scala 46:16:@12377.4]
  wire  _T_13492; // @[Mux.scala 46:19:@12378.4]
  wire [7:0] _T_13493; // @[Mux.scala 46:16:@12379.4]
  wire  _T_13494; // @[Mux.scala 46:19:@12380.4]
  wire [7:0] _T_13495; // @[Mux.scala 46:16:@12381.4]
  wire  _T_13496; // @[Mux.scala 46:19:@12382.4]
  wire [7:0] _T_13497; // @[Mux.scala 46:16:@12383.4]
  wire  _T_13498; // @[Mux.scala 46:19:@12384.4]
  wire [7:0] _T_13499; // @[Mux.scala 46:16:@12385.4]
  wire  _T_13500; // @[Mux.scala 46:19:@12386.4]
  wire [7:0] _T_13501; // @[Mux.scala 46:16:@12387.4]
  wire  _T_13502; // @[Mux.scala 46:19:@12388.4]
  wire [7:0] _T_13503; // @[Mux.scala 46:16:@12389.4]
  wire  _T_13504; // @[Mux.scala 46:19:@12390.4]
  wire [7:0] _T_13505; // @[Mux.scala 46:16:@12391.4]
  wire  _T_13506; // @[Mux.scala 46:19:@12392.4]
  wire [7:0] _T_13507; // @[Mux.scala 46:16:@12393.4]
  wire  _T_13508; // @[Mux.scala 46:19:@12394.4]
  wire [7:0] _T_13509; // @[Mux.scala 46:16:@12395.4]
  wire  _T_13510; // @[Mux.scala 46:19:@12396.4]
  wire [7:0] _T_13511; // @[Mux.scala 46:16:@12397.4]
  wire  _T_13512; // @[Mux.scala 46:19:@12398.4]
  wire [7:0] _T_13513; // @[Mux.scala 46:16:@12399.4]
  wire  _T_13514; // @[Mux.scala 46:19:@12400.4]
  wire [7:0] _T_13515; // @[Mux.scala 46:16:@12401.4]
  wire  _T_13516; // @[Mux.scala 46:19:@12402.4]
  wire [7:0] _T_13517; // @[Mux.scala 46:16:@12403.4]
  wire  _T_13518; // @[Mux.scala 46:19:@12404.4]
  wire [7:0] _T_13519; // @[Mux.scala 46:16:@12405.4]
  wire  _T_13520; // @[Mux.scala 46:19:@12406.4]
  wire [7:0] _T_13521; // @[Mux.scala 46:16:@12407.4]
  wire  _T_13522; // @[Mux.scala 46:19:@12408.4]
  wire [7:0] _T_13523; // @[Mux.scala 46:16:@12409.4]
  wire  _T_13524; // @[Mux.scala 46:19:@12410.4]
  wire [7:0] _T_13525; // @[Mux.scala 46:16:@12411.4]
  wire  _T_13526; // @[Mux.scala 46:19:@12412.4]
  wire [7:0] _T_13527; // @[Mux.scala 46:16:@12413.4]
  wire  _T_13528; // @[Mux.scala 46:19:@12414.4]
  wire [7:0] _T_13529; // @[Mux.scala 46:16:@12415.4]
  wire  _T_13530; // @[Mux.scala 46:19:@12416.4]
  wire [7:0] _T_13531; // @[Mux.scala 46:16:@12417.4]
  wire  _T_13532; // @[Mux.scala 46:19:@12418.4]
  wire [7:0] _T_13533; // @[Mux.scala 46:16:@12419.4]
  wire  _T_13534; // @[Mux.scala 46:19:@12420.4]
  wire [7:0] _T_13535; // @[Mux.scala 46:16:@12421.4]
  wire  _T_13536; // @[Mux.scala 46:19:@12422.4]
  wire [7:0] _T_13537; // @[Mux.scala 46:16:@12423.4]
  wire  _T_13538; // @[Mux.scala 46:19:@12424.4]
  wire [7:0] _T_13539; // @[Mux.scala 46:16:@12425.4]
  wire  _T_13540; // @[Mux.scala 46:19:@12426.4]
  wire [7:0] _T_13541; // @[Mux.scala 46:16:@12427.4]
  wire  _T_13542; // @[Mux.scala 46:19:@12428.4]
  wire [7:0] _T_13543; // @[Mux.scala 46:16:@12429.4]
  wire  _T_13544; // @[Mux.scala 46:19:@12430.4]
  wire [7:0] _T_13545; // @[Mux.scala 46:16:@12431.4]
  wire  _T_13546; // @[Mux.scala 46:19:@12432.4]
  wire [7:0] _T_13547; // @[Mux.scala 46:16:@12433.4]
  wire  _T_13548; // @[Mux.scala 46:19:@12434.4]
  wire [7:0] _T_13549; // @[Mux.scala 46:16:@12435.4]
  wire  _T_13588; // @[Mux.scala 46:19:@12437.4]
  wire [7:0] _T_13589; // @[Mux.scala 46:16:@12438.4]
  wire  _T_13590; // @[Mux.scala 46:19:@12439.4]
  wire [7:0] _T_13591; // @[Mux.scala 46:16:@12440.4]
  wire  _T_13592; // @[Mux.scala 46:19:@12441.4]
  wire [7:0] _T_13593; // @[Mux.scala 46:16:@12442.4]
  wire  _T_13594; // @[Mux.scala 46:19:@12443.4]
  wire [7:0] _T_13595; // @[Mux.scala 46:16:@12444.4]
  wire  _T_13596; // @[Mux.scala 46:19:@12445.4]
  wire [7:0] _T_13597; // @[Mux.scala 46:16:@12446.4]
  wire  _T_13598; // @[Mux.scala 46:19:@12447.4]
  wire [7:0] _T_13599; // @[Mux.scala 46:16:@12448.4]
  wire  _T_13600; // @[Mux.scala 46:19:@12449.4]
  wire [7:0] _T_13601; // @[Mux.scala 46:16:@12450.4]
  wire  _T_13602; // @[Mux.scala 46:19:@12451.4]
  wire [7:0] _T_13603; // @[Mux.scala 46:16:@12452.4]
  wire  _T_13604; // @[Mux.scala 46:19:@12453.4]
  wire [7:0] _T_13605; // @[Mux.scala 46:16:@12454.4]
  wire  _T_13606; // @[Mux.scala 46:19:@12455.4]
  wire [7:0] _T_13607; // @[Mux.scala 46:16:@12456.4]
  wire  _T_13608; // @[Mux.scala 46:19:@12457.4]
  wire [7:0] _T_13609; // @[Mux.scala 46:16:@12458.4]
  wire  _T_13610; // @[Mux.scala 46:19:@12459.4]
  wire [7:0] _T_13611; // @[Mux.scala 46:16:@12460.4]
  wire  _T_13612; // @[Mux.scala 46:19:@12461.4]
  wire [7:0] _T_13613; // @[Mux.scala 46:16:@12462.4]
  wire  _T_13614; // @[Mux.scala 46:19:@12463.4]
  wire [7:0] _T_13615; // @[Mux.scala 46:16:@12464.4]
  wire  _T_13616; // @[Mux.scala 46:19:@12465.4]
  wire [7:0] _T_13617; // @[Mux.scala 46:16:@12466.4]
  wire  _T_13618; // @[Mux.scala 46:19:@12467.4]
  wire [7:0] _T_13619; // @[Mux.scala 46:16:@12468.4]
  wire  _T_13620; // @[Mux.scala 46:19:@12469.4]
  wire [7:0] _T_13621; // @[Mux.scala 46:16:@12470.4]
  wire  _T_13622; // @[Mux.scala 46:19:@12471.4]
  wire [7:0] _T_13623; // @[Mux.scala 46:16:@12472.4]
  wire  _T_13624; // @[Mux.scala 46:19:@12473.4]
  wire [7:0] _T_13625; // @[Mux.scala 46:16:@12474.4]
  wire  _T_13626; // @[Mux.scala 46:19:@12475.4]
  wire [7:0] _T_13627; // @[Mux.scala 46:16:@12476.4]
  wire  _T_13628; // @[Mux.scala 46:19:@12477.4]
  wire [7:0] _T_13629; // @[Mux.scala 46:16:@12478.4]
  wire  _T_13630; // @[Mux.scala 46:19:@12479.4]
  wire [7:0] _T_13631; // @[Mux.scala 46:16:@12480.4]
  wire  _T_13632; // @[Mux.scala 46:19:@12481.4]
  wire [7:0] _T_13633; // @[Mux.scala 46:16:@12482.4]
  wire  _T_13634; // @[Mux.scala 46:19:@12483.4]
  wire [7:0] _T_13635; // @[Mux.scala 46:16:@12484.4]
  wire  _T_13636; // @[Mux.scala 46:19:@12485.4]
  wire [7:0] _T_13637; // @[Mux.scala 46:16:@12486.4]
  wire  _T_13638; // @[Mux.scala 46:19:@12487.4]
  wire [7:0] _T_13639; // @[Mux.scala 46:16:@12488.4]
  wire  _T_13640; // @[Mux.scala 46:19:@12489.4]
  wire [7:0] _T_13641; // @[Mux.scala 46:16:@12490.4]
  wire  _T_13642; // @[Mux.scala 46:19:@12491.4]
  wire [7:0] _T_13643; // @[Mux.scala 46:16:@12492.4]
  wire  _T_13644; // @[Mux.scala 46:19:@12493.4]
  wire [7:0] _T_13645; // @[Mux.scala 46:16:@12494.4]
  wire  _T_13646; // @[Mux.scala 46:19:@12495.4]
  wire [7:0] _T_13647; // @[Mux.scala 46:16:@12496.4]
  wire  _T_13648; // @[Mux.scala 46:19:@12497.4]
  wire [7:0] _T_13649; // @[Mux.scala 46:16:@12498.4]
  wire  _T_13650; // @[Mux.scala 46:19:@12499.4]
  wire [7:0] _T_13651; // @[Mux.scala 46:16:@12500.4]
  wire  _T_13652; // @[Mux.scala 46:19:@12501.4]
  wire [7:0] _T_13653; // @[Mux.scala 46:16:@12502.4]
  wire  _T_13654; // @[Mux.scala 46:19:@12503.4]
  wire [7:0] _T_13655; // @[Mux.scala 46:16:@12504.4]
  wire  _T_13656; // @[Mux.scala 46:19:@12505.4]
  wire [7:0] _T_13657; // @[Mux.scala 46:16:@12506.4]
  wire  _T_13658; // @[Mux.scala 46:19:@12507.4]
  wire [7:0] _T_13659; // @[Mux.scala 46:16:@12508.4]
  wire  _T_13660; // @[Mux.scala 46:19:@12509.4]
  wire [7:0] _T_13661; // @[Mux.scala 46:16:@12510.4]
  wire  _T_13701; // @[Mux.scala 46:19:@12512.4]
  wire [7:0] _T_13702; // @[Mux.scala 46:16:@12513.4]
  wire  _T_13703; // @[Mux.scala 46:19:@12514.4]
  wire [7:0] _T_13704; // @[Mux.scala 46:16:@12515.4]
  wire  _T_13705; // @[Mux.scala 46:19:@12516.4]
  wire [7:0] _T_13706; // @[Mux.scala 46:16:@12517.4]
  wire  _T_13707; // @[Mux.scala 46:19:@12518.4]
  wire [7:0] _T_13708; // @[Mux.scala 46:16:@12519.4]
  wire  _T_13709; // @[Mux.scala 46:19:@12520.4]
  wire [7:0] _T_13710; // @[Mux.scala 46:16:@12521.4]
  wire  _T_13711; // @[Mux.scala 46:19:@12522.4]
  wire [7:0] _T_13712; // @[Mux.scala 46:16:@12523.4]
  wire  _T_13713; // @[Mux.scala 46:19:@12524.4]
  wire [7:0] _T_13714; // @[Mux.scala 46:16:@12525.4]
  wire  _T_13715; // @[Mux.scala 46:19:@12526.4]
  wire [7:0] _T_13716; // @[Mux.scala 46:16:@12527.4]
  wire  _T_13717; // @[Mux.scala 46:19:@12528.4]
  wire [7:0] _T_13718; // @[Mux.scala 46:16:@12529.4]
  wire  _T_13719; // @[Mux.scala 46:19:@12530.4]
  wire [7:0] _T_13720; // @[Mux.scala 46:16:@12531.4]
  wire  _T_13721; // @[Mux.scala 46:19:@12532.4]
  wire [7:0] _T_13722; // @[Mux.scala 46:16:@12533.4]
  wire  _T_13723; // @[Mux.scala 46:19:@12534.4]
  wire [7:0] _T_13724; // @[Mux.scala 46:16:@12535.4]
  wire  _T_13725; // @[Mux.scala 46:19:@12536.4]
  wire [7:0] _T_13726; // @[Mux.scala 46:16:@12537.4]
  wire  _T_13727; // @[Mux.scala 46:19:@12538.4]
  wire [7:0] _T_13728; // @[Mux.scala 46:16:@12539.4]
  wire  _T_13729; // @[Mux.scala 46:19:@12540.4]
  wire [7:0] _T_13730; // @[Mux.scala 46:16:@12541.4]
  wire  _T_13731; // @[Mux.scala 46:19:@12542.4]
  wire [7:0] _T_13732; // @[Mux.scala 46:16:@12543.4]
  wire  _T_13733; // @[Mux.scala 46:19:@12544.4]
  wire [7:0] _T_13734; // @[Mux.scala 46:16:@12545.4]
  wire  _T_13735; // @[Mux.scala 46:19:@12546.4]
  wire [7:0] _T_13736; // @[Mux.scala 46:16:@12547.4]
  wire  _T_13737; // @[Mux.scala 46:19:@12548.4]
  wire [7:0] _T_13738; // @[Mux.scala 46:16:@12549.4]
  wire  _T_13739; // @[Mux.scala 46:19:@12550.4]
  wire [7:0] _T_13740; // @[Mux.scala 46:16:@12551.4]
  wire  _T_13741; // @[Mux.scala 46:19:@12552.4]
  wire [7:0] _T_13742; // @[Mux.scala 46:16:@12553.4]
  wire  _T_13743; // @[Mux.scala 46:19:@12554.4]
  wire [7:0] _T_13744; // @[Mux.scala 46:16:@12555.4]
  wire  _T_13745; // @[Mux.scala 46:19:@12556.4]
  wire [7:0] _T_13746; // @[Mux.scala 46:16:@12557.4]
  wire  _T_13747; // @[Mux.scala 46:19:@12558.4]
  wire [7:0] _T_13748; // @[Mux.scala 46:16:@12559.4]
  wire  _T_13749; // @[Mux.scala 46:19:@12560.4]
  wire [7:0] _T_13750; // @[Mux.scala 46:16:@12561.4]
  wire  _T_13751; // @[Mux.scala 46:19:@12562.4]
  wire [7:0] _T_13752; // @[Mux.scala 46:16:@12563.4]
  wire  _T_13753; // @[Mux.scala 46:19:@12564.4]
  wire [7:0] _T_13754; // @[Mux.scala 46:16:@12565.4]
  wire  _T_13755; // @[Mux.scala 46:19:@12566.4]
  wire [7:0] _T_13756; // @[Mux.scala 46:16:@12567.4]
  wire  _T_13757; // @[Mux.scala 46:19:@12568.4]
  wire [7:0] _T_13758; // @[Mux.scala 46:16:@12569.4]
  wire  _T_13759; // @[Mux.scala 46:19:@12570.4]
  wire [7:0] _T_13760; // @[Mux.scala 46:16:@12571.4]
  wire  _T_13761; // @[Mux.scala 46:19:@12572.4]
  wire [7:0] _T_13762; // @[Mux.scala 46:16:@12573.4]
  wire  _T_13763; // @[Mux.scala 46:19:@12574.4]
  wire [7:0] _T_13764; // @[Mux.scala 46:16:@12575.4]
  wire  _T_13765; // @[Mux.scala 46:19:@12576.4]
  wire [7:0] _T_13766; // @[Mux.scala 46:16:@12577.4]
  wire  _T_13767; // @[Mux.scala 46:19:@12578.4]
  wire [7:0] _T_13768; // @[Mux.scala 46:16:@12579.4]
  wire  _T_13769; // @[Mux.scala 46:19:@12580.4]
  wire [7:0] _T_13770; // @[Mux.scala 46:16:@12581.4]
  wire  _T_13771; // @[Mux.scala 46:19:@12582.4]
  wire [7:0] _T_13772; // @[Mux.scala 46:16:@12583.4]
  wire  _T_13773; // @[Mux.scala 46:19:@12584.4]
  wire [7:0] _T_13774; // @[Mux.scala 46:16:@12585.4]
  wire  _T_13775; // @[Mux.scala 46:19:@12586.4]
  wire [7:0] _T_13776; // @[Mux.scala 46:16:@12587.4]
  wire  _T_13817; // @[Mux.scala 46:19:@12589.4]
  wire [7:0] _T_13818; // @[Mux.scala 46:16:@12590.4]
  wire  _T_13819; // @[Mux.scala 46:19:@12591.4]
  wire [7:0] _T_13820; // @[Mux.scala 46:16:@12592.4]
  wire  _T_13821; // @[Mux.scala 46:19:@12593.4]
  wire [7:0] _T_13822; // @[Mux.scala 46:16:@12594.4]
  wire  _T_13823; // @[Mux.scala 46:19:@12595.4]
  wire [7:0] _T_13824; // @[Mux.scala 46:16:@12596.4]
  wire  _T_13825; // @[Mux.scala 46:19:@12597.4]
  wire [7:0] _T_13826; // @[Mux.scala 46:16:@12598.4]
  wire  _T_13827; // @[Mux.scala 46:19:@12599.4]
  wire [7:0] _T_13828; // @[Mux.scala 46:16:@12600.4]
  wire  _T_13829; // @[Mux.scala 46:19:@12601.4]
  wire [7:0] _T_13830; // @[Mux.scala 46:16:@12602.4]
  wire  _T_13831; // @[Mux.scala 46:19:@12603.4]
  wire [7:0] _T_13832; // @[Mux.scala 46:16:@12604.4]
  wire  _T_13833; // @[Mux.scala 46:19:@12605.4]
  wire [7:0] _T_13834; // @[Mux.scala 46:16:@12606.4]
  wire  _T_13835; // @[Mux.scala 46:19:@12607.4]
  wire [7:0] _T_13836; // @[Mux.scala 46:16:@12608.4]
  wire  _T_13837; // @[Mux.scala 46:19:@12609.4]
  wire [7:0] _T_13838; // @[Mux.scala 46:16:@12610.4]
  wire  _T_13839; // @[Mux.scala 46:19:@12611.4]
  wire [7:0] _T_13840; // @[Mux.scala 46:16:@12612.4]
  wire  _T_13841; // @[Mux.scala 46:19:@12613.4]
  wire [7:0] _T_13842; // @[Mux.scala 46:16:@12614.4]
  wire  _T_13843; // @[Mux.scala 46:19:@12615.4]
  wire [7:0] _T_13844; // @[Mux.scala 46:16:@12616.4]
  wire  _T_13845; // @[Mux.scala 46:19:@12617.4]
  wire [7:0] _T_13846; // @[Mux.scala 46:16:@12618.4]
  wire  _T_13847; // @[Mux.scala 46:19:@12619.4]
  wire [7:0] _T_13848; // @[Mux.scala 46:16:@12620.4]
  wire  _T_13849; // @[Mux.scala 46:19:@12621.4]
  wire [7:0] _T_13850; // @[Mux.scala 46:16:@12622.4]
  wire  _T_13851; // @[Mux.scala 46:19:@12623.4]
  wire [7:0] _T_13852; // @[Mux.scala 46:16:@12624.4]
  wire  _T_13853; // @[Mux.scala 46:19:@12625.4]
  wire [7:0] _T_13854; // @[Mux.scala 46:16:@12626.4]
  wire  _T_13855; // @[Mux.scala 46:19:@12627.4]
  wire [7:0] _T_13856; // @[Mux.scala 46:16:@12628.4]
  wire  _T_13857; // @[Mux.scala 46:19:@12629.4]
  wire [7:0] _T_13858; // @[Mux.scala 46:16:@12630.4]
  wire  _T_13859; // @[Mux.scala 46:19:@12631.4]
  wire [7:0] _T_13860; // @[Mux.scala 46:16:@12632.4]
  wire  _T_13861; // @[Mux.scala 46:19:@12633.4]
  wire [7:0] _T_13862; // @[Mux.scala 46:16:@12634.4]
  wire  _T_13863; // @[Mux.scala 46:19:@12635.4]
  wire [7:0] _T_13864; // @[Mux.scala 46:16:@12636.4]
  wire  _T_13865; // @[Mux.scala 46:19:@12637.4]
  wire [7:0] _T_13866; // @[Mux.scala 46:16:@12638.4]
  wire  _T_13867; // @[Mux.scala 46:19:@12639.4]
  wire [7:0] _T_13868; // @[Mux.scala 46:16:@12640.4]
  wire  _T_13869; // @[Mux.scala 46:19:@12641.4]
  wire [7:0] _T_13870; // @[Mux.scala 46:16:@12642.4]
  wire  _T_13871; // @[Mux.scala 46:19:@12643.4]
  wire [7:0] _T_13872; // @[Mux.scala 46:16:@12644.4]
  wire  _T_13873; // @[Mux.scala 46:19:@12645.4]
  wire [7:0] _T_13874; // @[Mux.scala 46:16:@12646.4]
  wire  _T_13875; // @[Mux.scala 46:19:@12647.4]
  wire [7:0] _T_13876; // @[Mux.scala 46:16:@12648.4]
  wire  _T_13877; // @[Mux.scala 46:19:@12649.4]
  wire [7:0] _T_13878; // @[Mux.scala 46:16:@12650.4]
  wire  _T_13879; // @[Mux.scala 46:19:@12651.4]
  wire [7:0] _T_13880; // @[Mux.scala 46:16:@12652.4]
  wire  _T_13881; // @[Mux.scala 46:19:@12653.4]
  wire [7:0] _T_13882; // @[Mux.scala 46:16:@12654.4]
  wire  _T_13883; // @[Mux.scala 46:19:@12655.4]
  wire [7:0] _T_13884; // @[Mux.scala 46:16:@12656.4]
  wire  _T_13885; // @[Mux.scala 46:19:@12657.4]
  wire [7:0] _T_13886; // @[Mux.scala 46:16:@12658.4]
  wire  _T_13887; // @[Mux.scala 46:19:@12659.4]
  wire [7:0] _T_13888; // @[Mux.scala 46:16:@12660.4]
  wire  _T_13889; // @[Mux.scala 46:19:@12661.4]
  wire [7:0] _T_13890; // @[Mux.scala 46:16:@12662.4]
  wire  _T_13891; // @[Mux.scala 46:19:@12663.4]
  wire [7:0] _T_13892; // @[Mux.scala 46:16:@12664.4]
  wire  _T_13893; // @[Mux.scala 46:19:@12665.4]
  wire [7:0] _T_13894; // @[Mux.scala 46:16:@12666.4]
  wire  _T_13936; // @[Mux.scala 46:19:@12668.4]
  wire [7:0] _T_13937; // @[Mux.scala 46:16:@12669.4]
  wire  _T_13938; // @[Mux.scala 46:19:@12670.4]
  wire [7:0] _T_13939; // @[Mux.scala 46:16:@12671.4]
  wire  _T_13940; // @[Mux.scala 46:19:@12672.4]
  wire [7:0] _T_13941; // @[Mux.scala 46:16:@12673.4]
  wire  _T_13942; // @[Mux.scala 46:19:@12674.4]
  wire [7:0] _T_13943; // @[Mux.scala 46:16:@12675.4]
  wire  _T_13944; // @[Mux.scala 46:19:@12676.4]
  wire [7:0] _T_13945; // @[Mux.scala 46:16:@12677.4]
  wire  _T_13946; // @[Mux.scala 46:19:@12678.4]
  wire [7:0] _T_13947; // @[Mux.scala 46:16:@12679.4]
  wire  _T_13948; // @[Mux.scala 46:19:@12680.4]
  wire [7:0] _T_13949; // @[Mux.scala 46:16:@12681.4]
  wire  _T_13950; // @[Mux.scala 46:19:@12682.4]
  wire [7:0] _T_13951; // @[Mux.scala 46:16:@12683.4]
  wire  _T_13952; // @[Mux.scala 46:19:@12684.4]
  wire [7:0] _T_13953; // @[Mux.scala 46:16:@12685.4]
  wire  _T_13954; // @[Mux.scala 46:19:@12686.4]
  wire [7:0] _T_13955; // @[Mux.scala 46:16:@12687.4]
  wire  _T_13956; // @[Mux.scala 46:19:@12688.4]
  wire [7:0] _T_13957; // @[Mux.scala 46:16:@12689.4]
  wire  _T_13958; // @[Mux.scala 46:19:@12690.4]
  wire [7:0] _T_13959; // @[Mux.scala 46:16:@12691.4]
  wire  _T_13960; // @[Mux.scala 46:19:@12692.4]
  wire [7:0] _T_13961; // @[Mux.scala 46:16:@12693.4]
  wire  _T_13962; // @[Mux.scala 46:19:@12694.4]
  wire [7:0] _T_13963; // @[Mux.scala 46:16:@12695.4]
  wire  _T_13964; // @[Mux.scala 46:19:@12696.4]
  wire [7:0] _T_13965; // @[Mux.scala 46:16:@12697.4]
  wire  _T_13966; // @[Mux.scala 46:19:@12698.4]
  wire [7:0] _T_13967; // @[Mux.scala 46:16:@12699.4]
  wire  _T_13968; // @[Mux.scala 46:19:@12700.4]
  wire [7:0] _T_13969; // @[Mux.scala 46:16:@12701.4]
  wire  _T_13970; // @[Mux.scala 46:19:@12702.4]
  wire [7:0] _T_13971; // @[Mux.scala 46:16:@12703.4]
  wire  _T_13972; // @[Mux.scala 46:19:@12704.4]
  wire [7:0] _T_13973; // @[Mux.scala 46:16:@12705.4]
  wire  _T_13974; // @[Mux.scala 46:19:@12706.4]
  wire [7:0] _T_13975; // @[Mux.scala 46:16:@12707.4]
  wire  _T_13976; // @[Mux.scala 46:19:@12708.4]
  wire [7:0] _T_13977; // @[Mux.scala 46:16:@12709.4]
  wire  _T_13978; // @[Mux.scala 46:19:@12710.4]
  wire [7:0] _T_13979; // @[Mux.scala 46:16:@12711.4]
  wire  _T_13980; // @[Mux.scala 46:19:@12712.4]
  wire [7:0] _T_13981; // @[Mux.scala 46:16:@12713.4]
  wire  _T_13982; // @[Mux.scala 46:19:@12714.4]
  wire [7:0] _T_13983; // @[Mux.scala 46:16:@12715.4]
  wire  _T_13984; // @[Mux.scala 46:19:@12716.4]
  wire [7:0] _T_13985; // @[Mux.scala 46:16:@12717.4]
  wire  _T_13986; // @[Mux.scala 46:19:@12718.4]
  wire [7:0] _T_13987; // @[Mux.scala 46:16:@12719.4]
  wire  _T_13988; // @[Mux.scala 46:19:@12720.4]
  wire [7:0] _T_13989; // @[Mux.scala 46:16:@12721.4]
  wire  _T_13990; // @[Mux.scala 46:19:@12722.4]
  wire [7:0] _T_13991; // @[Mux.scala 46:16:@12723.4]
  wire  _T_13992; // @[Mux.scala 46:19:@12724.4]
  wire [7:0] _T_13993; // @[Mux.scala 46:16:@12725.4]
  wire  _T_13994; // @[Mux.scala 46:19:@12726.4]
  wire [7:0] _T_13995; // @[Mux.scala 46:16:@12727.4]
  wire  _T_13996; // @[Mux.scala 46:19:@12728.4]
  wire [7:0] _T_13997; // @[Mux.scala 46:16:@12729.4]
  wire  _T_13998; // @[Mux.scala 46:19:@12730.4]
  wire [7:0] _T_13999; // @[Mux.scala 46:16:@12731.4]
  wire  _T_14000; // @[Mux.scala 46:19:@12732.4]
  wire [7:0] _T_14001; // @[Mux.scala 46:16:@12733.4]
  wire  _T_14002; // @[Mux.scala 46:19:@12734.4]
  wire [7:0] _T_14003; // @[Mux.scala 46:16:@12735.4]
  wire  _T_14004; // @[Mux.scala 46:19:@12736.4]
  wire [7:0] _T_14005; // @[Mux.scala 46:16:@12737.4]
  wire  _T_14006; // @[Mux.scala 46:19:@12738.4]
  wire [7:0] _T_14007; // @[Mux.scala 46:16:@12739.4]
  wire  _T_14008; // @[Mux.scala 46:19:@12740.4]
  wire [7:0] _T_14009; // @[Mux.scala 46:16:@12741.4]
  wire  _T_14010; // @[Mux.scala 46:19:@12742.4]
  wire [7:0] _T_14011; // @[Mux.scala 46:16:@12743.4]
  wire  _T_14012; // @[Mux.scala 46:19:@12744.4]
  wire [7:0] _T_14013; // @[Mux.scala 46:16:@12745.4]
  wire  _T_14014; // @[Mux.scala 46:19:@12746.4]
  wire [7:0] _T_14015; // @[Mux.scala 46:16:@12747.4]
  wire  _T_14058; // @[Mux.scala 46:19:@12749.4]
  wire [7:0] _T_14059; // @[Mux.scala 46:16:@12750.4]
  wire  _T_14060; // @[Mux.scala 46:19:@12751.4]
  wire [7:0] _T_14061; // @[Mux.scala 46:16:@12752.4]
  wire  _T_14062; // @[Mux.scala 46:19:@12753.4]
  wire [7:0] _T_14063; // @[Mux.scala 46:16:@12754.4]
  wire  _T_14064; // @[Mux.scala 46:19:@12755.4]
  wire [7:0] _T_14065; // @[Mux.scala 46:16:@12756.4]
  wire  _T_14066; // @[Mux.scala 46:19:@12757.4]
  wire [7:0] _T_14067; // @[Mux.scala 46:16:@12758.4]
  wire  _T_14068; // @[Mux.scala 46:19:@12759.4]
  wire [7:0] _T_14069; // @[Mux.scala 46:16:@12760.4]
  wire  _T_14070; // @[Mux.scala 46:19:@12761.4]
  wire [7:0] _T_14071; // @[Mux.scala 46:16:@12762.4]
  wire  _T_14072; // @[Mux.scala 46:19:@12763.4]
  wire [7:0] _T_14073; // @[Mux.scala 46:16:@12764.4]
  wire  _T_14074; // @[Mux.scala 46:19:@12765.4]
  wire [7:0] _T_14075; // @[Mux.scala 46:16:@12766.4]
  wire  _T_14076; // @[Mux.scala 46:19:@12767.4]
  wire [7:0] _T_14077; // @[Mux.scala 46:16:@12768.4]
  wire  _T_14078; // @[Mux.scala 46:19:@12769.4]
  wire [7:0] _T_14079; // @[Mux.scala 46:16:@12770.4]
  wire  _T_14080; // @[Mux.scala 46:19:@12771.4]
  wire [7:0] _T_14081; // @[Mux.scala 46:16:@12772.4]
  wire  _T_14082; // @[Mux.scala 46:19:@12773.4]
  wire [7:0] _T_14083; // @[Mux.scala 46:16:@12774.4]
  wire  _T_14084; // @[Mux.scala 46:19:@12775.4]
  wire [7:0] _T_14085; // @[Mux.scala 46:16:@12776.4]
  wire  _T_14086; // @[Mux.scala 46:19:@12777.4]
  wire [7:0] _T_14087; // @[Mux.scala 46:16:@12778.4]
  wire  _T_14088; // @[Mux.scala 46:19:@12779.4]
  wire [7:0] _T_14089; // @[Mux.scala 46:16:@12780.4]
  wire  _T_14090; // @[Mux.scala 46:19:@12781.4]
  wire [7:0] _T_14091; // @[Mux.scala 46:16:@12782.4]
  wire  _T_14092; // @[Mux.scala 46:19:@12783.4]
  wire [7:0] _T_14093; // @[Mux.scala 46:16:@12784.4]
  wire  _T_14094; // @[Mux.scala 46:19:@12785.4]
  wire [7:0] _T_14095; // @[Mux.scala 46:16:@12786.4]
  wire  _T_14096; // @[Mux.scala 46:19:@12787.4]
  wire [7:0] _T_14097; // @[Mux.scala 46:16:@12788.4]
  wire  _T_14098; // @[Mux.scala 46:19:@12789.4]
  wire [7:0] _T_14099; // @[Mux.scala 46:16:@12790.4]
  wire  _T_14100; // @[Mux.scala 46:19:@12791.4]
  wire [7:0] _T_14101; // @[Mux.scala 46:16:@12792.4]
  wire  _T_14102; // @[Mux.scala 46:19:@12793.4]
  wire [7:0] _T_14103; // @[Mux.scala 46:16:@12794.4]
  wire  _T_14104; // @[Mux.scala 46:19:@12795.4]
  wire [7:0] _T_14105; // @[Mux.scala 46:16:@12796.4]
  wire  _T_14106; // @[Mux.scala 46:19:@12797.4]
  wire [7:0] _T_14107; // @[Mux.scala 46:16:@12798.4]
  wire  _T_14108; // @[Mux.scala 46:19:@12799.4]
  wire [7:0] _T_14109; // @[Mux.scala 46:16:@12800.4]
  wire  _T_14110; // @[Mux.scala 46:19:@12801.4]
  wire [7:0] _T_14111; // @[Mux.scala 46:16:@12802.4]
  wire  _T_14112; // @[Mux.scala 46:19:@12803.4]
  wire [7:0] _T_14113; // @[Mux.scala 46:16:@12804.4]
  wire  _T_14114; // @[Mux.scala 46:19:@12805.4]
  wire [7:0] _T_14115; // @[Mux.scala 46:16:@12806.4]
  wire  _T_14116; // @[Mux.scala 46:19:@12807.4]
  wire [7:0] _T_14117; // @[Mux.scala 46:16:@12808.4]
  wire  _T_14118; // @[Mux.scala 46:19:@12809.4]
  wire [7:0] _T_14119; // @[Mux.scala 46:16:@12810.4]
  wire  _T_14120; // @[Mux.scala 46:19:@12811.4]
  wire [7:0] _T_14121; // @[Mux.scala 46:16:@12812.4]
  wire  _T_14122; // @[Mux.scala 46:19:@12813.4]
  wire [7:0] _T_14123; // @[Mux.scala 46:16:@12814.4]
  wire  _T_14124; // @[Mux.scala 46:19:@12815.4]
  wire [7:0] _T_14125; // @[Mux.scala 46:16:@12816.4]
  wire  _T_14126; // @[Mux.scala 46:19:@12817.4]
  wire [7:0] _T_14127; // @[Mux.scala 46:16:@12818.4]
  wire  _T_14128; // @[Mux.scala 46:19:@12819.4]
  wire [7:0] _T_14129; // @[Mux.scala 46:16:@12820.4]
  wire  _T_14130; // @[Mux.scala 46:19:@12821.4]
  wire [7:0] _T_14131; // @[Mux.scala 46:16:@12822.4]
  wire  _T_14132; // @[Mux.scala 46:19:@12823.4]
  wire [7:0] _T_14133; // @[Mux.scala 46:16:@12824.4]
  wire  _T_14134; // @[Mux.scala 46:19:@12825.4]
  wire [7:0] _T_14135; // @[Mux.scala 46:16:@12826.4]
  wire  _T_14136; // @[Mux.scala 46:19:@12827.4]
  wire [7:0] _T_14137; // @[Mux.scala 46:16:@12828.4]
  wire  _T_14138; // @[Mux.scala 46:19:@12829.4]
  wire [7:0] _T_14139; // @[Mux.scala 46:16:@12830.4]
  wire  _T_14183; // @[Mux.scala 46:19:@12832.4]
  wire [7:0] _T_14184; // @[Mux.scala 46:16:@12833.4]
  wire  _T_14185; // @[Mux.scala 46:19:@12834.4]
  wire [7:0] _T_14186; // @[Mux.scala 46:16:@12835.4]
  wire  _T_14187; // @[Mux.scala 46:19:@12836.4]
  wire [7:0] _T_14188; // @[Mux.scala 46:16:@12837.4]
  wire  _T_14189; // @[Mux.scala 46:19:@12838.4]
  wire [7:0] _T_14190; // @[Mux.scala 46:16:@12839.4]
  wire  _T_14191; // @[Mux.scala 46:19:@12840.4]
  wire [7:0] _T_14192; // @[Mux.scala 46:16:@12841.4]
  wire  _T_14193; // @[Mux.scala 46:19:@12842.4]
  wire [7:0] _T_14194; // @[Mux.scala 46:16:@12843.4]
  wire  _T_14195; // @[Mux.scala 46:19:@12844.4]
  wire [7:0] _T_14196; // @[Mux.scala 46:16:@12845.4]
  wire  _T_14197; // @[Mux.scala 46:19:@12846.4]
  wire [7:0] _T_14198; // @[Mux.scala 46:16:@12847.4]
  wire  _T_14199; // @[Mux.scala 46:19:@12848.4]
  wire [7:0] _T_14200; // @[Mux.scala 46:16:@12849.4]
  wire  _T_14201; // @[Mux.scala 46:19:@12850.4]
  wire [7:0] _T_14202; // @[Mux.scala 46:16:@12851.4]
  wire  _T_14203; // @[Mux.scala 46:19:@12852.4]
  wire [7:0] _T_14204; // @[Mux.scala 46:16:@12853.4]
  wire  _T_14205; // @[Mux.scala 46:19:@12854.4]
  wire [7:0] _T_14206; // @[Mux.scala 46:16:@12855.4]
  wire  _T_14207; // @[Mux.scala 46:19:@12856.4]
  wire [7:0] _T_14208; // @[Mux.scala 46:16:@12857.4]
  wire  _T_14209; // @[Mux.scala 46:19:@12858.4]
  wire [7:0] _T_14210; // @[Mux.scala 46:16:@12859.4]
  wire  _T_14211; // @[Mux.scala 46:19:@12860.4]
  wire [7:0] _T_14212; // @[Mux.scala 46:16:@12861.4]
  wire  _T_14213; // @[Mux.scala 46:19:@12862.4]
  wire [7:0] _T_14214; // @[Mux.scala 46:16:@12863.4]
  wire  _T_14215; // @[Mux.scala 46:19:@12864.4]
  wire [7:0] _T_14216; // @[Mux.scala 46:16:@12865.4]
  wire  _T_14217; // @[Mux.scala 46:19:@12866.4]
  wire [7:0] _T_14218; // @[Mux.scala 46:16:@12867.4]
  wire  _T_14219; // @[Mux.scala 46:19:@12868.4]
  wire [7:0] _T_14220; // @[Mux.scala 46:16:@12869.4]
  wire  _T_14221; // @[Mux.scala 46:19:@12870.4]
  wire [7:0] _T_14222; // @[Mux.scala 46:16:@12871.4]
  wire  _T_14223; // @[Mux.scala 46:19:@12872.4]
  wire [7:0] _T_14224; // @[Mux.scala 46:16:@12873.4]
  wire  _T_14225; // @[Mux.scala 46:19:@12874.4]
  wire [7:0] _T_14226; // @[Mux.scala 46:16:@12875.4]
  wire  _T_14227; // @[Mux.scala 46:19:@12876.4]
  wire [7:0] _T_14228; // @[Mux.scala 46:16:@12877.4]
  wire  _T_14229; // @[Mux.scala 46:19:@12878.4]
  wire [7:0] _T_14230; // @[Mux.scala 46:16:@12879.4]
  wire  _T_14231; // @[Mux.scala 46:19:@12880.4]
  wire [7:0] _T_14232; // @[Mux.scala 46:16:@12881.4]
  wire  _T_14233; // @[Mux.scala 46:19:@12882.4]
  wire [7:0] _T_14234; // @[Mux.scala 46:16:@12883.4]
  wire  _T_14235; // @[Mux.scala 46:19:@12884.4]
  wire [7:0] _T_14236; // @[Mux.scala 46:16:@12885.4]
  wire  _T_14237; // @[Mux.scala 46:19:@12886.4]
  wire [7:0] _T_14238; // @[Mux.scala 46:16:@12887.4]
  wire  _T_14239; // @[Mux.scala 46:19:@12888.4]
  wire [7:0] _T_14240; // @[Mux.scala 46:16:@12889.4]
  wire  _T_14241; // @[Mux.scala 46:19:@12890.4]
  wire [7:0] _T_14242; // @[Mux.scala 46:16:@12891.4]
  wire  _T_14243; // @[Mux.scala 46:19:@12892.4]
  wire [7:0] _T_14244; // @[Mux.scala 46:16:@12893.4]
  wire  _T_14245; // @[Mux.scala 46:19:@12894.4]
  wire [7:0] _T_14246; // @[Mux.scala 46:16:@12895.4]
  wire  _T_14247; // @[Mux.scala 46:19:@12896.4]
  wire [7:0] _T_14248; // @[Mux.scala 46:16:@12897.4]
  wire  _T_14249; // @[Mux.scala 46:19:@12898.4]
  wire [7:0] _T_14250; // @[Mux.scala 46:16:@12899.4]
  wire  _T_14251; // @[Mux.scala 46:19:@12900.4]
  wire [7:0] _T_14252; // @[Mux.scala 46:16:@12901.4]
  wire  _T_14253; // @[Mux.scala 46:19:@12902.4]
  wire [7:0] _T_14254; // @[Mux.scala 46:16:@12903.4]
  wire  _T_14255; // @[Mux.scala 46:19:@12904.4]
  wire [7:0] _T_14256; // @[Mux.scala 46:16:@12905.4]
  wire  _T_14257; // @[Mux.scala 46:19:@12906.4]
  wire [7:0] _T_14258; // @[Mux.scala 46:16:@12907.4]
  wire  _T_14259; // @[Mux.scala 46:19:@12908.4]
  wire [7:0] _T_14260; // @[Mux.scala 46:16:@12909.4]
  wire  _T_14261; // @[Mux.scala 46:19:@12910.4]
  wire [7:0] _T_14262; // @[Mux.scala 46:16:@12911.4]
  wire  _T_14263; // @[Mux.scala 46:19:@12912.4]
  wire [7:0] _T_14264; // @[Mux.scala 46:16:@12913.4]
  wire  _T_14265; // @[Mux.scala 46:19:@12914.4]
  wire [7:0] _T_14266; // @[Mux.scala 46:16:@12915.4]
  wire  _T_14311; // @[Mux.scala 46:19:@12917.4]
  wire [7:0] _T_14312; // @[Mux.scala 46:16:@12918.4]
  wire  _T_14313; // @[Mux.scala 46:19:@12919.4]
  wire [7:0] _T_14314; // @[Mux.scala 46:16:@12920.4]
  wire  _T_14315; // @[Mux.scala 46:19:@12921.4]
  wire [7:0] _T_14316; // @[Mux.scala 46:16:@12922.4]
  wire  _T_14317; // @[Mux.scala 46:19:@12923.4]
  wire [7:0] _T_14318; // @[Mux.scala 46:16:@12924.4]
  wire  _T_14319; // @[Mux.scala 46:19:@12925.4]
  wire [7:0] _T_14320; // @[Mux.scala 46:16:@12926.4]
  wire  _T_14321; // @[Mux.scala 46:19:@12927.4]
  wire [7:0] _T_14322; // @[Mux.scala 46:16:@12928.4]
  wire  _T_14323; // @[Mux.scala 46:19:@12929.4]
  wire [7:0] _T_14324; // @[Mux.scala 46:16:@12930.4]
  wire  _T_14325; // @[Mux.scala 46:19:@12931.4]
  wire [7:0] _T_14326; // @[Mux.scala 46:16:@12932.4]
  wire  _T_14327; // @[Mux.scala 46:19:@12933.4]
  wire [7:0] _T_14328; // @[Mux.scala 46:16:@12934.4]
  wire  _T_14329; // @[Mux.scala 46:19:@12935.4]
  wire [7:0] _T_14330; // @[Mux.scala 46:16:@12936.4]
  wire  _T_14331; // @[Mux.scala 46:19:@12937.4]
  wire [7:0] _T_14332; // @[Mux.scala 46:16:@12938.4]
  wire  _T_14333; // @[Mux.scala 46:19:@12939.4]
  wire [7:0] _T_14334; // @[Mux.scala 46:16:@12940.4]
  wire  _T_14335; // @[Mux.scala 46:19:@12941.4]
  wire [7:0] _T_14336; // @[Mux.scala 46:16:@12942.4]
  wire  _T_14337; // @[Mux.scala 46:19:@12943.4]
  wire [7:0] _T_14338; // @[Mux.scala 46:16:@12944.4]
  wire  _T_14339; // @[Mux.scala 46:19:@12945.4]
  wire [7:0] _T_14340; // @[Mux.scala 46:16:@12946.4]
  wire  _T_14341; // @[Mux.scala 46:19:@12947.4]
  wire [7:0] _T_14342; // @[Mux.scala 46:16:@12948.4]
  wire  _T_14343; // @[Mux.scala 46:19:@12949.4]
  wire [7:0] _T_14344; // @[Mux.scala 46:16:@12950.4]
  wire  _T_14345; // @[Mux.scala 46:19:@12951.4]
  wire [7:0] _T_14346; // @[Mux.scala 46:16:@12952.4]
  wire  _T_14347; // @[Mux.scala 46:19:@12953.4]
  wire [7:0] _T_14348; // @[Mux.scala 46:16:@12954.4]
  wire  _T_14349; // @[Mux.scala 46:19:@12955.4]
  wire [7:0] _T_14350; // @[Mux.scala 46:16:@12956.4]
  wire  _T_14351; // @[Mux.scala 46:19:@12957.4]
  wire [7:0] _T_14352; // @[Mux.scala 46:16:@12958.4]
  wire  _T_14353; // @[Mux.scala 46:19:@12959.4]
  wire [7:0] _T_14354; // @[Mux.scala 46:16:@12960.4]
  wire  _T_14355; // @[Mux.scala 46:19:@12961.4]
  wire [7:0] _T_14356; // @[Mux.scala 46:16:@12962.4]
  wire  _T_14357; // @[Mux.scala 46:19:@12963.4]
  wire [7:0] _T_14358; // @[Mux.scala 46:16:@12964.4]
  wire  _T_14359; // @[Mux.scala 46:19:@12965.4]
  wire [7:0] _T_14360; // @[Mux.scala 46:16:@12966.4]
  wire  _T_14361; // @[Mux.scala 46:19:@12967.4]
  wire [7:0] _T_14362; // @[Mux.scala 46:16:@12968.4]
  wire  _T_14363; // @[Mux.scala 46:19:@12969.4]
  wire [7:0] _T_14364; // @[Mux.scala 46:16:@12970.4]
  wire  _T_14365; // @[Mux.scala 46:19:@12971.4]
  wire [7:0] _T_14366; // @[Mux.scala 46:16:@12972.4]
  wire  _T_14367; // @[Mux.scala 46:19:@12973.4]
  wire [7:0] _T_14368; // @[Mux.scala 46:16:@12974.4]
  wire  _T_14369; // @[Mux.scala 46:19:@12975.4]
  wire [7:0] _T_14370; // @[Mux.scala 46:16:@12976.4]
  wire  _T_14371; // @[Mux.scala 46:19:@12977.4]
  wire [7:0] _T_14372; // @[Mux.scala 46:16:@12978.4]
  wire  _T_14373; // @[Mux.scala 46:19:@12979.4]
  wire [7:0] _T_14374; // @[Mux.scala 46:16:@12980.4]
  wire  _T_14375; // @[Mux.scala 46:19:@12981.4]
  wire [7:0] _T_14376; // @[Mux.scala 46:16:@12982.4]
  wire  _T_14377; // @[Mux.scala 46:19:@12983.4]
  wire [7:0] _T_14378; // @[Mux.scala 46:16:@12984.4]
  wire  _T_14379; // @[Mux.scala 46:19:@12985.4]
  wire [7:0] _T_14380; // @[Mux.scala 46:16:@12986.4]
  wire  _T_14381; // @[Mux.scala 46:19:@12987.4]
  wire [7:0] _T_14382; // @[Mux.scala 46:16:@12988.4]
  wire  _T_14383; // @[Mux.scala 46:19:@12989.4]
  wire [7:0] _T_14384; // @[Mux.scala 46:16:@12990.4]
  wire  _T_14385; // @[Mux.scala 46:19:@12991.4]
  wire [7:0] _T_14386; // @[Mux.scala 46:16:@12992.4]
  wire  _T_14387; // @[Mux.scala 46:19:@12993.4]
  wire [7:0] _T_14388; // @[Mux.scala 46:16:@12994.4]
  wire  _T_14389; // @[Mux.scala 46:19:@12995.4]
  wire [7:0] _T_14390; // @[Mux.scala 46:16:@12996.4]
  wire  _T_14391; // @[Mux.scala 46:19:@12997.4]
  wire [7:0] _T_14392; // @[Mux.scala 46:16:@12998.4]
  wire  _T_14393; // @[Mux.scala 46:19:@12999.4]
  wire [7:0] _T_14394; // @[Mux.scala 46:16:@13000.4]
  wire  _T_14395; // @[Mux.scala 46:19:@13001.4]
  wire [7:0] _T_14396; // @[Mux.scala 46:16:@13002.4]
  wire  _T_14442; // @[Mux.scala 46:19:@13004.4]
  wire [7:0] _T_14443; // @[Mux.scala 46:16:@13005.4]
  wire  _T_14444; // @[Mux.scala 46:19:@13006.4]
  wire [7:0] _T_14445; // @[Mux.scala 46:16:@13007.4]
  wire  _T_14446; // @[Mux.scala 46:19:@13008.4]
  wire [7:0] _T_14447; // @[Mux.scala 46:16:@13009.4]
  wire  _T_14448; // @[Mux.scala 46:19:@13010.4]
  wire [7:0] _T_14449; // @[Mux.scala 46:16:@13011.4]
  wire  _T_14450; // @[Mux.scala 46:19:@13012.4]
  wire [7:0] _T_14451; // @[Mux.scala 46:16:@13013.4]
  wire  _T_14452; // @[Mux.scala 46:19:@13014.4]
  wire [7:0] _T_14453; // @[Mux.scala 46:16:@13015.4]
  wire  _T_14454; // @[Mux.scala 46:19:@13016.4]
  wire [7:0] _T_14455; // @[Mux.scala 46:16:@13017.4]
  wire  _T_14456; // @[Mux.scala 46:19:@13018.4]
  wire [7:0] _T_14457; // @[Mux.scala 46:16:@13019.4]
  wire  _T_14458; // @[Mux.scala 46:19:@13020.4]
  wire [7:0] _T_14459; // @[Mux.scala 46:16:@13021.4]
  wire  _T_14460; // @[Mux.scala 46:19:@13022.4]
  wire [7:0] _T_14461; // @[Mux.scala 46:16:@13023.4]
  wire  _T_14462; // @[Mux.scala 46:19:@13024.4]
  wire [7:0] _T_14463; // @[Mux.scala 46:16:@13025.4]
  wire  _T_14464; // @[Mux.scala 46:19:@13026.4]
  wire [7:0] _T_14465; // @[Mux.scala 46:16:@13027.4]
  wire  _T_14466; // @[Mux.scala 46:19:@13028.4]
  wire [7:0] _T_14467; // @[Mux.scala 46:16:@13029.4]
  wire  _T_14468; // @[Mux.scala 46:19:@13030.4]
  wire [7:0] _T_14469; // @[Mux.scala 46:16:@13031.4]
  wire  _T_14470; // @[Mux.scala 46:19:@13032.4]
  wire [7:0] _T_14471; // @[Mux.scala 46:16:@13033.4]
  wire  _T_14472; // @[Mux.scala 46:19:@13034.4]
  wire [7:0] _T_14473; // @[Mux.scala 46:16:@13035.4]
  wire  _T_14474; // @[Mux.scala 46:19:@13036.4]
  wire [7:0] _T_14475; // @[Mux.scala 46:16:@13037.4]
  wire  _T_14476; // @[Mux.scala 46:19:@13038.4]
  wire [7:0] _T_14477; // @[Mux.scala 46:16:@13039.4]
  wire  _T_14478; // @[Mux.scala 46:19:@13040.4]
  wire [7:0] _T_14479; // @[Mux.scala 46:16:@13041.4]
  wire  _T_14480; // @[Mux.scala 46:19:@13042.4]
  wire [7:0] _T_14481; // @[Mux.scala 46:16:@13043.4]
  wire  _T_14482; // @[Mux.scala 46:19:@13044.4]
  wire [7:0] _T_14483; // @[Mux.scala 46:16:@13045.4]
  wire  _T_14484; // @[Mux.scala 46:19:@13046.4]
  wire [7:0] _T_14485; // @[Mux.scala 46:16:@13047.4]
  wire  _T_14486; // @[Mux.scala 46:19:@13048.4]
  wire [7:0] _T_14487; // @[Mux.scala 46:16:@13049.4]
  wire  _T_14488; // @[Mux.scala 46:19:@13050.4]
  wire [7:0] _T_14489; // @[Mux.scala 46:16:@13051.4]
  wire  _T_14490; // @[Mux.scala 46:19:@13052.4]
  wire [7:0] _T_14491; // @[Mux.scala 46:16:@13053.4]
  wire  _T_14492; // @[Mux.scala 46:19:@13054.4]
  wire [7:0] _T_14493; // @[Mux.scala 46:16:@13055.4]
  wire  _T_14494; // @[Mux.scala 46:19:@13056.4]
  wire [7:0] _T_14495; // @[Mux.scala 46:16:@13057.4]
  wire  _T_14496; // @[Mux.scala 46:19:@13058.4]
  wire [7:0] _T_14497; // @[Mux.scala 46:16:@13059.4]
  wire  _T_14498; // @[Mux.scala 46:19:@13060.4]
  wire [7:0] _T_14499; // @[Mux.scala 46:16:@13061.4]
  wire  _T_14500; // @[Mux.scala 46:19:@13062.4]
  wire [7:0] _T_14501; // @[Mux.scala 46:16:@13063.4]
  wire  _T_14502; // @[Mux.scala 46:19:@13064.4]
  wire [7:0] _T_14503; // @[Mux.scala 46:16:@13065.4]
  wire  _T_14504; // @[Mux.scala 46:19:@13066.4]
  wire [7:0] _T_14505; // @[Mux.scala 46:16:@13067.4]
  wire  _T_14506; // @[Mux.scala 46:19:@13068.4]
  wire [7:0] _T_14507; // @[Mux.scala 46:16:@13069.4]
  wire  _T_14508; // @[Mux.scala 46:19:@13070.4]
  wire [7:0] _T_14509; // @[Mux.scala 46:16:@13071.4]
  wire  _T_14510; // @[Mux.scala 46:19:@13072.4]
  wire [7:0] _T_14511; // @[Mux.scala 46:16:@13073.4]
  wire  _T_14512; // @[Mux.scala 46:19:@13074.4]
  wire [7:0] _T_14513; // @[Mux.scala 46:16:@13075.4]
  wire  _T_14514; // @[Mux.scala 46:19:@13076.4]
  wire [7:0] _T_14515; // @[Mux.scala 46:16:@13077.4]
  wire  _T_14516; // @[Mux.scala 46:19:@13078.4]
  wire [7:0] _T_14517; // @[Mux.scala 46:16:@13079.4]
  wire  _T_14518; // @[Mux.scala 46:19:@13080.4]
  wire [7:0] _T_14519; // @[Mux.scala 46:16:@13081.4]
  wire  _T_14520; // @[Mux.scala 46:19:@13082.4]
  wire [7:0] _T_14521; // @[Mux.scala 46:16:@13083.4]
  wire  _T_14522; // @[Mux.scala 46:19:@13084.4]
  wire [7:0] _T_14523; // @[Mux.scala 46:16:@13085.4]
  wire  _T_14524; // @[Mux.scala 46:19:@13086.4]
  wire [7:0] _T_14525; // @[Mux.scala 46:16:@13087.4]
  wire  _T_14526; // @[Mux.scala 46:19:@13088.4]
  wire [7:0] _T_14527; // @[Mux.scala 46:16:@13089.4]
  wire  _T_14528; // @[Mux.scala 46:19:@13090.4]
  wire [7:0] _T_14529; // @[Mux.scala 46:16:@13091.4]
  wire  _T_14576; // @[Mux.scala 46:19:@13093.4]
  wire [7:0] _T_14577; // @[Mux.scala 46:16:@13094.4]
  wire  _T_14578; // @[Mux.scala 46:19:@13095.4]
  wire [7:0] _T_14579; // @[Mux.scala 46:16:@13096.4]
  wire  _T_14580; // @[Mux.scala 46:19:@13097.4]
  wire [7:0] _T_14581; // @[Mux.scala 46:16:@13098.4]
  wire  _T_14582; // @[Mux.scala 46:19:@13099.4]
  wire [7:0] _T_14583; // @[Mux.scala 46:16:@13100.4]
  wire  _T_14584; // @[Mux.scala 46:19:@13101.4]
  wire [7:0] _T_14585; // @[Mux.scala 46:16:@13102.4]
  wire  _T_14586; // @[Mux.scala 46:19:@13103.4]
  wire [7:0] _T_14587; // @[Mux.scala 46:16:@13104.4]
  wire  _T_14588; // @[Mux.scala 46:19:@13105.4]
  wire [7:0] _T_14589; // @[Mux.scala 46:16:@13106.4]
  wire  _T_14590; // @[Mux.scala 46:19:@13107.4]
  wire [7:0] _T_14591; // @[Mux.scala 46:16:@13108.4]
  wire  _T_14592; // @[Mux.scala 46:19:@13109.4]
  wire [7:0] _T_14593; // @[Mux.scala 46:16:@13110.4]
  wire  _T_14594; // @[Mux.scala 46:19:@13111.4]
  wire [7:0] _T_14595; // @[Mux.scala 46:16:@13112.4]
  wire  _T_14596; // @[Mux.scala 46:19:@13113.4]
  wire [7:0] _T_14597; // @[Mux.scala 46:16:@13114.4]
  wire  _T_14598; // @[Mux.scala 46:19:@13115.4]
  wire [7:0] _T_14599; // @[Mux.scala 46:16:@13116.4]
  wire  _T_14600; // @[Mux.scala 46:19:@13117.4]
  wire [7:0] _T_14601; // @[Mux.scala 46:16:@13118.4]
  wire  _T_14602; // @[Mux.scala 46:19:@13119.4]
  wire [7:0] _T_14603; // @[Mux.scala 46:16:@13120.4]
  wire  _T_14604; // @[Mux.scala 46:19:@13121.4]
  wire [7:0] _T_14605; // @[Mux.scala 46:16:@13122.4]
  wire  _T_14606; // @[Mux.scala 46:19:@13123.4]
  wire [7:0] _T_14607; // @[Mux.scala 46:16:@13124.4]
  wire  _T_14608; // @[Mux.scala 46:19:@13125.4]
  wire [7:0] _T_14609; // @[Mux.scala 46:16:@13126.4]
  wire  _T_14610; // @[Mux.scala 46:19:@13127.4]
  wire [7:0] _T_14611; // @[Mux.scala 46:16:@13128.4]
  wire  _T_14612; // @[Mux.scala 46:19:@13129.4]
  wire [7:0] _T_14613; // @[Mux.scala 46:16:@13130.4]
  wire  _T_14614; // @[Mux.scala 46:19:@13131.4]
  wire [7:0] _T_14615; // @[Mux.scala 46:16:@13132.4]
  wire  _T_14616; // @[Mux.scala 46:19:@13133.4]
  wire [7:0] _T_14617; // @[Mux.scala 46:16:@13134.4]
  wire  _T_14618; // @[Mux.scala 46:19:@13135.4]
  wire [7:0] _T_14619; // @[Mux.scala 46:16:@13136.4]
  wire  _T_14620; // @[Mux.scala 46:19:@13137.4]
  wire [7:0] _T_14621; // @[Mux.scala 46:16:@13138.4]
  wire  _T_14622; // @[Mux.scala 46:19:@13139.4]
  wire [7:0] _T_14623; // @[Mux.scala 46:16:@13140.4]
  wire  _T_14624; // @[Mux.scala 46:19:@13141.4]
  wire [7:0] _T_14625; // @[Mux.scala 46:16:@13142.4]
  wire  _T_14626; // @[Mux.scala 46:19:@13143.4]
  wire [7:0] _T_14627; // @[Mux.scala 46:16:@13144.4]
  wire  _T_14628; // @[Mux.scala 46:19:@13145.4]
  wire [7:0] _T_14629; // @[Mux.scala 46:16:@13146.4]
  wire  _T_14630; // @[Mux.scala 46:19:@13147.4]
  wire [7:0] _T_14631; // @[Mux.scala 46:16:@13148.4]
  wire  _T_14632; // @[Mux.scala 46:19:@13149.4]
  wire [7:0] _T_14633; // @[Mux.scala 46:16:@13150.4]
  wire  _T_14634; // @[Mux.scala 46:19:@13151.4]
  wire [7:0] _T_14635; // @[Mux.scala 46:16:@13152.4]
  wire  _T_14636; // @[Mux.scala 46:19:@13153.4]
  wire [7:0] _T_14637; // @[Mux.scala 46:16:@13154.4]
  wire  _T_14638; // @[Mux.scala 46:19:@13155.4]
  wire [7:0] _T_14639; // @[Mux.scala 46:16:@13156.4]
  wire  _T_14640; // @[Mux.scala 46:19:@13157.4]
  wire [7:0] _T_14641; // @[Mux.scala 46:16:@13158.4]
  wire  _T_14642; // @[Mux.scala 46:19:@13159.4]
  wire [7:0] _T_14643; // @[Mux.scala 46:16:@13160.4]
  wire  _T_14644; // @[Mux.scala 46:19:@13161.4]
  wire [7:0] _T_14645; // @[Mux.scala 46:16:@13162.4]
  wire  _T_14646; // @[Mux.scala 46:19:@13163.4]
  wire [7:0] _T_14647; // @[Mux.scala 46:16:@13164.4]
  wire  _T_14648; // @[Mux.scala 46:19:@13165.4]
  wire [7:0] _T_14649; // @[Mux.scala 46:16:@13166.4]
  wire  _T_14650; // @[Mux.scala 46:19:@13167.4]
  wire [7:0] _T_14651; // @[Mux.scala 46:16:@13168.4]
  wire  _T_14652; // @[Mux.scala 46:19:@13169.4]
  wire [7:0] _T_14653; // @[Mux.scala 46:16:@13170.4]
  wire  _T_14654; // @[Mux.scala 46:19:@13171.4]
  wire [7:0] _T_14655; // @[Mux.scala 46:16:@13172.4]
  wire  _T_14656; // @[Mux.scala 46:19:@13173.4]
  wire [7:0] _T_14657; // @[Mux.scala 46:16:@13174.4]
  wire  _T_14658; // @[Mux.scala 46:19:@13175.4]
  wire [7:0] _T_14659; // @[Mux.scala 46:16:@13176.4]
  wire  _T_14660; // @[Mux.scala 46:19:@13177.4]
  wire [7:0] _T_14661; // @[Mux.scala 46:16:@13178.4]
  wire  _T_14662; // @[Mux.scala 46:19:@13179.4]
  wire [7:0] _T_14663; // @[Mux.scala 46:16:@13180.4]
  wire  _T_14664; // @[Mux.scala 46:19:@13181.4]
  wire [7:0] _T_14665; // @[Mux.scala 46:16:@13182.4]
  wire  _T_14713; // @[Mux.scala 46:19:@13184.4]
  wire [7:0] _T_14714; // @[Mux.scala 46:16:@13185.4]
  wire  _T_14715; // @[Mux.scala 46:19:@13186.4]
  wire [7:0] _T_14716; // @[Mux.scala 46:16:@13187.4]
  wire  _T_14717; // @[Mux.scala 46:19:@13188.4]
  wire [7:0] _T_14718; // @[Mux.scala 46:16:@13189.4]
  wire  _T_14719; // @[Mux.scala 46:19:@13190.4]
  wire [7:0] _T_14720; // @[Mux.scala 46:16:@13191.4]
  wire  _T_14721; // @[Mux.scala 46:19:@13192.4]
  wire [7:0] _T_14722; // @[Mux.scala 46:16:@13193.4]
  wire  _T_14723; // @[Mux.scala 46:19:@13194.4]
  wire [7:0] _T_14724; // @[Mux.scala 46:16:@13195.4]
  wire  _T_14725; // @[Mux.scala 46:19:@13196.4]
  wire [7:0] _T_14726; // @[Mux.scala 46:16:@13197.4]
  wire  _T_14727; // @[Mux.scala 46:19:@13198.4]
  wire [7:0] _T_14728; // @[Mux.scala 46:16:@13199.4]
  wire  _T_14729; // @[Mux.scala 46:19:@13200.4]
  wire [7:0] _T_14730; // @[Mux.scala 46:16:@13201.4]
  wire  _T_14731; // @[Mux.scala 46:19:@13202.4]
  wire [7:0] _T_14732; // @[Mux.scala 46:16:@13203.4]
  wire  _T_14733; // @[Mux.scala 46:19:@13204.4]
  wire [7:0] _T_14734; // @[Mux.scala 46:16:@13205.4]
  wire  _T_14735; // @[Mux.scala 46:19:@13206.4]
  wire [7:0] _T_14736; // @[Mux.scala 46:16:@13207.4]
  wire  _T_14737; // @[Mux.scala 46:19:@13208.4]
  wire [7:0] _T_14738; // @[Mux.scala 46:16:@13209.4]
  wire  _T_14739; // @[Mux.scala 46:19:@13210.4]
  wire [7:0] _T_14740; // @[Mux.scala 46:16:@13211.4]
  wire  _T_14741; // @[Mux.scala 46:19:@13212.4]
  wire [7:0] _T_14742; // @[Mux.scala 46:16:@13213.4]
  wire  _T_14743; // @[Mux.scala 46:19:@13214.4]
  wire [7:0] _T_14744; // @[Mux.scala 46:16:@13215.4]
  wire  _T_14745; // @[Mux.scala 46:19:@13216.4]
  wire [7:0] _T_14746; // @[Mux.scala 46:16:@13217.4]
  wire  _T_14747; // @[Mux.scala 46:19:@13218.4]
  wire [7:0] _T_14748; // @[Mux.scala 46:16:@13219.4]
  wire  _T_14749; // @[Mux.scala 46:19:@13220.4]
  wire [7:0] _T_14750; // @[Mux.scala 46:16:@13221.4]
  wire  _T_14751; // @[Mux.scala 46:19:@13222.4]
  wire [7:0] _T_14752; // @[Mux.scala 46:16:@13223.4]
  wire  _T_14753; // @[Mux.scala 46:19:@13224.4]
  wire [7:0] _T_14754; // @[Mux.scala 46:16:@13225.4]
  wire  _T_14755; // @[Mux.scala 46:19:@13226.4]
  wire [7:0] _T_14756; // @[Mux.scala 46:16:@13227.4]
  wire  _T_14757; // @[Mux.scala 46:19:@13228.4]
  wire [7:0] _T_14758; // @[Mux.scala 46:16:@13229.4]
  wire  _T_14759; // @[Mux.scala 46:19:@13230.4]
  wire [7:0] _T_14760; // @[Mux.scala 46:16:@13231.4]
  wire  _T_14761; // @[Mux.scala 46:19:@13232.4]
  wire [7:0] _T_14762; // @[Mux.scala 46:16:@13233.4]
  wire  _T_14763; // @[Mux.scala 46:19:@13234.4]
  wire [7:0] _T_14764; // @[Mux.scala 46:16:@13235.4]
  wire  _T_14765; // @[Mux.scala 46:19:@13236.4]
  wire [7:0] _T_14766; // @[Mux.scala 46:16:@13237.4]
  wire  _T_14767; // @[Mux.scala 46:19:@13238.4]
  wire [7:0] _T_14768; // @[Mux.scala 46:16:@13239.4]
  wire  _T_14769; // @[Mux.scala 46:19:@13240.4]
  wire [7:0] _T_14770; // @[Mux.scala 46:16:@13241.4]
  wire  _T_14771; // @[Mux.scala 46:19:@13242.4]
  wire [7:0] _T_14772; // @[Mux.scala 46:16:@13243.4]
  wire  _T_14773; // @[Mux.scala 46:19:@13244.4]
  wire [7:0] _T_14774; // @[Mux.scala 46:16:@13245.4]
  wire  _T_14775; // @[Mux.scala 46:19:@13246.4]
  wire [7:0] _T_14776; // @[Mux.scala 46:16:@13247.4]
  wire  _T_14777; // @[Mux.scala 46:19:@13248.4]
  wire [7:0] _T_14778; // @[Mux.scala 46:16:@13249.4]
  wire  _T_14779; // @[Mux.scala 46:19:@13250.4]
  wire [7:0] _T_14780; // @[Mux.scala 46:16:@13251.4]
  wire  _T_14781; // @[Mux.scala 46:19:@13252.4]
  wire [7:0] _T_14782; // @[Mux.scala 46:16:@13253.4]
  wire  _T_14783; // @[Mux.scala 46:19:@13254.4]
  wire [7:0] _T_14784; // @[Mux.scala 46:16:@13255.4]
  wire  _T_14785; // @[Mux.scala 46:19:@13256.4]
  wire [7:0] _T_14786; // @[Mux.scala 46:16:@13257.4]
  wire  _T_14787; // @[Mux.scala 46:19:@13258.4]
  wire [7:0] _T_14788; // @[Mux.scala 46:16:@13259.4]
  wire  _T_14789; // @[Mux.scala 46:19:@13260.4]
  wire [7:0] _T_14790; // @[Mux.scala 46:16:@13261.4]
  wire  _T_14791; // @[Mux.scala 46:19:@13262.4]
  wire [7:0] _T_14792; // @[Mux.scala 46:16:@13263.4]
  wire  _T_14793; // @[Mux.scala 46:19:@13264.4]
  wire [7:0] _T_14794; // @[Mux.scala 46:16:@13265.4]
  wire  _T_14795; // @[Mux.scala 46:19:@13266.4]
  wire [7:0] _T_14796; // @[Mux.scala 46:16:@13267.4]
  wire  _T_14797; // @[Mux.scala 46:19:@13268.4]
  wire [7:0] _T_14798; // @[Mux.scala 46:16:@13269.4]
  wire  _T_14799; // @[Mux.scala 46:19:@13270.4]
  wire [7:0] _T_14800; // @[Mux.scala 46:16:@13271.4]
  wire  _T_14801; // @[Mux.scala 46:19:@13272.4]
  wire [7:0] _T_14802; // @[Mux.scala 46:16:@13273.4]
  wire  _T_14803; // @[Mux.scala 46:19:@13274.4]
  wire [7:0] _T_14804; // @[Mux.scala 46:16:@13275.4]
  wire  _T_14853; // @[Mux.scala 46:19:@13277.4]
  wire [7:0] _T_14854; // @[Mux.scala 46:16:@13278.4]
  wire  _T_14855; // @[Mux.scala 46:19:@13279.4]
  wire [7:0] _T_14856; // @[Mux.scala 46:16:@13280.4]
  wire  _T_14857; // @[Mux.scala 46:19:@13281.4]
  wire [7:0] _T_14858; // @[Mux.scala 46:16:@13282.4]
  wire  _T_14859; // @[Mux.scala 46:19:@13283.4]
  wire [7:0] _T_14860; // @[Mux.scala 46:16:@13284.4]
  wire  _T_14861; // @[Mux.scala 46:19:@13285.4]
  wire [7:0] _T_14862; // @[Mux.scala 46:16:@13286.4]
  wire  _T_14863; // @[Mux.scala 46:19:@13287.4]
  wire [7:0] _T_14864; // @[Mux.scala 46:16:@13288.4]
  wire  _T_14865; // @[Mux.scala 46:19:@13289.4]
  wire [7:0] _T_14866; // @[Mux.scala 46:16:@13290.4]
  wire  _T_14867; // @[Mux.scala 46:19:@13291.4]
  wire [7:0] _T_14868; // @[Mux.scala 46:16:@13292.4]
  wire  _T_14869; // @[Mux.scala 46:19:@13293.4]
  wire [7:0] _T_14870; // @[Mux.scala 46:16:@13294.4]
  wire  _T_14871; // @[Mux.scala 46:19:@13295.4]
  wire [7:0] _T_14872; // @[Mux.scala 46:16:@13296.4]
  wire  _T_14873; // @[Mux.scala 46:19:@13297.4]
  wire [7:0] _T_14874; // @[Mux.scala 46:16:@13298.4]
  wire  _T_14875; // @[Mux.scala 46:19:@13299.4]
  wire [7:0] _T_14876; // @[Mux.scala 46:16:@13300.4]
  wire  _T_14877; // @[Mux.scala 46:19:@13301.4]
  wire [7:0] _T_14878; // @[Mux.scala 46:16:@13302.4]
  wire  _T_14879; // @[Mux.scala 46:19:@13303.4]
  wire [7:0] _T_14880; // @[Mux.scala 46:16:@13304.4]
  wire  _T_14881; // @[Mux.scala 46:19:@13305.4]
  wire [7:0] _T_14882; // @[Mux.scala 46:16:@13306.4]
  wire  _T_14883; // @[Mux.scala 46:19:@13307.4]
  wire [7:0] _T_14884; // @[Mux.scala 46:16:@13308.4]
  wire  _T_14885; // @[Mux.scala 46:19:@13309.4]
  wire [7:0] _T_14886; // @[Mux.scala 46:16:@13310.4]
  wire  _T_14887; // @[Mux.scala 46:19:@13311.4]
  wire [7:0] _T_14888; // @[Mux.scala 46:16:@13312.4]
  wire  _T_14889; // @[Mux.scala 46:19:@13313.4]
  wire [7:0] _T_14890; // @[Mux.scala 46:16:@13314.4]
  wire  _T_14891; // @[Mux.scala 46:19:@13315.4]
  wire [7:0] _T_14892; // @[Mux.scala 46:16:@13316.4]
  wire  _T_14893; // @[Mux.scala 46:19:@13317.4]
  wire [7:0] _T_14894; // @[Mux.scala 46:16:@13318.4]
  wire  _T_14895; // @[Mux.scala 46:19:@13319.4]
  wire [7:0] _T_14896; // @[Mux.scala 46:16:@13320.4]
  wire  _T_14897; // @[Mux.scala 46:19:@13321.4]
  wire [7:0] _T_14898; // @[Mux.scala 46:16:@13322.4]
  wire  _T_14899; // @[Mux.scala 46:19:@13323.4]
  wire [7:0] _T_14900; // @[Mux.scala 46:16:@13324.4]
  wire  _T_14901; // @[Mux.scala 46:19:@13325.4]
  wire [7:0] _T_14902; // @[Mux.scala 46:16:@13326.4]
  wire  _T_14903; // @[Mux.scala 46:19:@13327.4]
  wire [7:0] _T_14904; // @[Mux.scala 46:16:@13328.4]
  wire  _T_14905; // @[Mux.scala 46:19:@13329.4]
  wire [7:0] _T_14906; // @[Mux.scala 46:16:@13330.4]
  wire  _T_14907; // @[Mux.scala 46:19:@13331.4]
  wire [7:0] _T_14908; // @[Mux.scala 46:16:@13332.4]
  wire  _T_14909; // @[Mux.scala 46:19:@13333.4]
  wire [7:0] _T_14910; // @[Mux.scala 46:16:@13334.4]
  wire  _T_14911; // @[Mux.scala 46:19:@13335.4]
  wire [7:0] _T_14912; // @[Mux.scala 46:16:@13336.4]
  wire  _T_14913; // @[Mux.scala 46:19:@13337.4]
  wire [7:0] _T_14914; // @[Mux.scala 46:16:@13338.4]
  wire  _T_14915; // @[Mux.scala 46:19:@13339.4]
  wire [7:0] _T_14916; // @[Mux.scala 46:16:@13340.4]
  wire  _T_14917; // @[Mux.scala 46:19:@13341.4]
  wire [7:0] _T_14918; // @[Mux.scala 46:16:@13342.4]
  wire  _T_14919; // @[Mux.scala 46:19:@13343.4]
  wire [7:0] _T_14920; // @[Mux.scala 46:16:@13344.4]
  wire  _T_14921; // @[Mux.scala 46:19:@13345.4]
  wire [7:0] _T_14922; // @[Mux.scala 46:16:@13346.4]
  wire  _T_14923; // @[Mux.scala 46:19:@13347.4]
  wire [7:0] _T_14924; // @[Mux.scala 46:16:@13348.4]
  wire  _T_14925; // @[Mux.scala 46:19:@13349.4]
  wire [7:0] _T_14926; // @[Mux.scala 46:16:@13350.4]
  wire  _T_14927; // @[Mux.scala 46:19:@13351.4]
  wire [7:0] _T_14928; // @[Mux.scala 46:16:@13352.4]
  wire  _T_14929; // @[Mux.scala 46:19:@13353.4]
  wire [7:0] _T_14930; // @[Mux.scala 46:16:@13354.4]
  wire  _T_14931; // @[Mux.scala 46:19:@13355.4]
  wire [7:0] _T_14932; // @[Mux.scala 46:16:@13356.4]
  wire  _T_14933; // @[Mux.scala 46:19:@13357.4]
  wire [7:0] _T_14934; // @[Mux.scala 46:16:@13358.4]
  wire  _T_14935; // @[Mux.scala 46:19:@13359.4]
  wire [7:0] _T_14936; // @[Mux.scala 46:16:@13360.4]
  wire  _T_14937; // @[Mux.scala 46:19:@13361.4]
  wire [7:0] _T_14938; // @[Mux.scala 46:16:@13362.4]
  wire  _T_14939; // @[Mux.scala 46:19:@13363.4]
  wire [7:0] _T_14940; // @[Mux.scala 46:16:@13364.4]
  wire  _T_14941; // @[Mux.scala 46:19:@13365.4]
  wire [7:0] _T_14942; // @[Mux.scala 46:16:@13366.4]
  wire  _T_14943; // @[Mux.scala 46:19:@13367.4]
  wire [7:0] _T_14944; // @[Mux.scala 46:16:@13368.4]
  wire  _T_14945; // @[Mux.scala 46:19:@13369.4]
  wire [7:0] _T_14946; // @[Mux.scala 46:16:@13370.4]
  wire  _T_14996; // @[Mux.scala 46:19:@13372.4]
  wire [7:0] _T_14997; // @[Mux.scala 46:16:@13373.4]
  wire  _T_14998; // @[Mux.scala 46:19:@13374.4]
  wire [7:0] _T_14999; // @[Mux.scala 46:16:@13375.4]
  wire  _T_15000; // @[Mux.scala 46:19:@13376.4]
  wire [7:0] _T_15001; // @[Mux.scala 46:16:@13377.4]
  wire  _T_15002; // @[Mux.scala 46:19:@13378.4]
  wire [7:0] _T_15003; // @[Mux.scala 46:16:@13379.4]
  wire  _T_15004; // @[Mux.scala 46:19:@13380.4]
  wire [7:0] _T_15005; // @[Mux.scala 46:16:@13381.4]
  wire  _T_15006; // @[Mux.scala 46:19:@13382.4]
  wire [7:0] _T_15007; // @[Mux.scala 46:16:@13383.4]
  wire  _T_15008; // @[Mux.scala 46:19:@13384.4]
  wire [7:0] _T_15009; // @[Mux.scala 46:16:@13385.4]
  wire  _T_15010; // @[Mux.scala 46:19:@13386.4]
  wire [7:0] _T_15011; // @[Mux.scala 46:16:@13387.4]
  wire  _T_15012; // @[Mux.scala 46:19:@13388.4]
  wire [7:0] _T_15013; // @[Mux.scala 46:16:@13389.4]
  wire  _T_15014; // @[Mux.scala 46:19:@13390.4]
  wire [7:0] _T_15015; // @[Mux.scala 46:16:@13391.4]
  wire  _T_15016; // @[Mux.scala 46:19:@13392.4]
  wire [7:0] _T_15017; // @[Mux.scala 46:16:@13393.4]
  wire  _T_15018; // @[Mux.scala 46:19:@13394.4]
  wire [7:0] _T_15019; // @[Mux.scala 46:16:@13395.4]
  wire  _T_15020; // @[Mux.scala 46:19:@13396.4]
  wire [7:0] _T_15021; // @[Mux.scala 46:16:@13397.4]
  wire  _T_15022; // @[Mux.scala 46:19:@13398.4]
  wire [7:0] _T_15023; // @[Mux.scala 46:16:@13399.4]
  wire  _T_15024; // @[Mux.scala 46:19:@13400.4]
  wire [7:0] _T_15025; // @[Mux.scala 46:16:@13401.4]
  wire  _T_15026; // @[Mux.scala 46:19:@13402.4]
  wire [7:0] _T_15027; // @[Mux.scala 46:16:@13403.4]
  wire  _T_15028; // @[Mux.scala 46:19:@13404.4]
  wire [7:0] _T_15029; // @[Mux.scala 46:16:@13405.4]
  wire  _T_15030; // @[Mux.scala 46:19:@13406.4]
  wire [7:0] _T_15031; // @[Mux.scala 46:16:@13407.4]
  wire  _T_15032; // @[Mux.scala 46:19:@13408.4]
  wire [7:0] _T_15033; // @[Mux.scala 46:16:@13409.4]
  wire  _T_15034; // @[Mux.scala 46:19:@13410.4]
  wire [7:0] _T_15035; // @[Mux.scala 46:16:@13411.4]
  wire  _T_15036; // @[Mux.scala 46:19:@13412.4]
  wire [7:0] _T_15037; // @[Mux.scala 46:16:@13413.4]
  wire  _T_15038; // @[Mux.scala 46:19:@13414.4]
  wire [7:0] _T_15039; // @[Mux.scala 46:16:@13415.4]
  wire  _T_15040; // @[Mux.scala 46:19:@13416.4]
  wire [7:0] _T_15041; // @[Mux.scala 46:16:@13417.4]
  wire  _T_15042; // @[Mux.scala 46:19:@13418.4]
  wire [7:0] _T_15043; // @[Mux.scala 46:16:@13419.4]
  wire  _T_15044; // @[Mux.scala 46:19:@13420.4]
  wire [7:0] _T_15045; // @[Mux.scala 46:16:@13421.4]
  wire  _T_15046; // @[Mux.scala 46:19:@13422.4]
  wire [7:0] _T_15047; // @[Mux.scala 46:16:@13423.4]
  wire  _T_15048; // @[Mux.scala 46:19:@13424.4]
  wire [7:0] _T_15049; // @[Mux.scala 46:16:@13425.4]
  wire  _T_15050; // @[Mux.scala 46:19:@13426.4]
  wire [7:0] _T_15051; // @[Mux.scala 46:16:@13427.4]
  wire  _T_15052; // @[Mux.scala 46:19:@13428.4]
  wire [7:0] _T_15053; // @[Mux.scala 46:16:@13429.4]
  wire  _T_15054; // @[Mux.scala 46:19:@13430.4]
  wire [7:0] _T_15055; // @[Mux.scala 46:16:@13431.4]
  wire  _T_15056; // @[Mux.scala 46:19:@13432.4]
  wire [7:0] _T_15057; // @[Mux.scala 46:16:@13433.4]
  wire  _T_15058; // @[Mux.scala 46:19:@13434.4]
  wire [7:0] _T_15059; // @[Mux.scala 46:16:@13435.4]
  wire  _T_15060; // @[Mux.scala 46:19:@13436.4]
  wire [7:0] _T_15061; // @[Mux.scala 46:16:@13437.4]
  wire  _T_15062; // @[Mux.scala 46:19:@13438.4]
  wire [7:0] _T_15063; // @[Mux.scala 46:16:@13439.4]
  wire  _T_15064; // @[Mux.scala 46:19:@13440.4]
  wire [7:0] _T_15065; // @[Mux.scala 46:16:@13441.4]
  wire  _T_15066; // @[Mux.scala 46:19:@13442.4]
  wire [7:0] _T_15067; // @[Mux.scala 46:16:@13443.4]
  wire  _T_15068; // @[Mux.scala 46:19:@13444.4]
  wire [7:0] _T_15069; // @[Mux.scala 46:16:@13445.4]
  wire  _T_15070; // @[Mux.scala 46:19:@13446.4]
  wire [7:0] _T_15071; // @[Mux.scala 46:16:@13447.4]
  wire  _T_15072; // @[Mux.scala 46:19:@13448.4]
  wire [7:0] _T_15073; // @[Mux.scala 46:16:@13449.4]
  wire  _T_15074; // @[Mux.scala 46:19:@13450.4]
  wire [7:0] _T_15075; // @[Mux.scala 46:16:@13451.4]
  wire  _T_15076; // @[Mux.scala 46:19:@13452.4]
  wire [7:0] _T_15077; // @[Mux.scala 46:16:@13453.4]
  wire  _T_15078; // @[Mux.scala 46:19:@13454.4]
  wire [7:0] _T_15079; // @[Mux.scala 46:16:@13455.4]
  wire  _T_15080; // @[Mux.scala 46:19:@13456.4]
  wire [7:0] _T_15081; // @[Mux.scala 46:16:@13457.4]
  wire  _T_15082; // @[Mux.scala 46:19:@13458.4]
  wire [7:0] _T_15083; // @[Mux.scala 46:16:@13459.4]
  wire  _T_15084; // @[Mux.scala 46:19:@13460.4]
  wire [7:0] _T_15085; // @[Mux.scala 46:16:@13461.4]
  wire  _T_15086; // @[Mux.scala 46:19:@13462.4]
  wire [7:0] _T_15087; // @[Mux.scala 46:16:@13463.4]
  wire  _T_15088; // @[Mux.scala 46:19:@13464.4]
  wire [7:0] _T_15089; // @[Mux.scala 46:16:@13465.4]
  wire  _T_15090; // @[Mux.scala 46:19:@13466.4]
  wire [7:0] _T_15091; // @[Mux.scala 46:16:@13467.4]
  wire  _T_15142; // @[Mux.scala 46:19:@13469.4]
  wire [7:0] _T_15143; // @[Mux.scala 46:16:@13470.4]
  wire  _T_15144; // @[Mux.scala 46:19:@13471.4]
  wire [7:0] _T_15145; // @[Mux.scala 46:16:@13472.4]
  wire  _T_15146; // @[Mux.scala 46:19:@13473.4]
  wire [7:0] _T_15147; // @[Mux.scala 46:16:@13474.4]
  wire  _T_15148; // @[Mux.scala 46:19:@13475.4]
  wire [7:0] _T_15149; // @[Mux.scala 46:16:@13476.4]
  wire  _T_15150; // @[Mux.scala 46:19:@13477.4]
  wire [7:0] _T_15151; // @[Mux.scala 46:16:@13478.4]
  wire  _T_15152; // @[Mux.scala 46:19:@13479.4]
  wire [7:0] _T_15153; // @[Mux.scala 46:16:@13480.4]
  wire  _T_15154; // @[Mux.scala 46:19:@13481.4]
  wire [7:0] _T_15155; // @[Mux.scala 46:16:@13482.4]
  wire  _T_15156; // @[Mux.scala 46:19:@13483.4]
  wire [7:0] _T_15157; // @[Mux.scala 46:16:@13484.4]
  wire  _T_15158; // @[Mux.scala 46:19:@13485.4]
  wire [7:0] _T_15159; // @[Mux.scala 46:16:@13486.4]
  wire  _T_15160; // @[Mux.scala 46:19:@13487.4]
  wire [7:0] _T_15161; // @[Mux.scala 46:16:@13488.4]
  wire  _T_15162; // @[Mux.scala 46:19:@13489.4]
  wire [7:0] _T_15163; // @[Mux.scala 46:16:@13490.4]
  wire  _T_15164; // @[Mux.scala 46:19:@13491.4]
  wire [7:0] _T_15165; // @[Mux.scala 46:16:@13492.4]
  wire  _T_15166; // @[Mux.scala 46:19:@13493.4]
  wire [7:0] _T_15167; // @[Mux.scala 46:16:@13494.4]
  wire  _T_15168; // @[Mux.scala 46:19:@13495.4]
  wire [7:0] _T_15169; // @[Mux.scala 46:16:@13496.4]
  wire  _T_15170; // @[Mux.scala 46:19:@13497.4]
  wire [7:0] _T_15171; // @[Mux.scala 46:16:@13498.4]
  wire  _T_15172; // @[Mux.scala 46:19:@13499.4]
  wire [7:0] _T_15173; // @[Mux.scala 46:16:@13500.4]
  wire  _T_15174; // @[Mux.scala 46:19:@13501.4]
  wire [7:0] _T_15175; // @[Mux.scala 46:16:@13502.4]
  wire  _T_15176; // @[Mux.scala 46:19:@13503.4]
  wire [7:0] _T_15177; // @[Mux.scala 46:16:@13504.4]
  wire  _T_15178; // @[Mux.scala 46:19:@13505.4]
  wire [7:0] _T_15179; // @[Mux.scala 46:16:@13506.4]
  wire  _T_15180; // @[Mux.scala 46:19:@13507.4]
  wire [7:0] _T_15181; // @[Mux.scala 46:16:@13508.4]
  wire  _T_15182; // @[Mux.scala 46:19:@13509.4]
  wire [7:0] _T_15183; // @[Mux.scala 46:16:@13510.4]
  wire  _T_15184; // @[Mux.scala 46:19:@13511.4]
  wire [7:0] _T_15185; // @[Mux.scala 46:16:@13512.4]
  wire  _T_15186; // @[Mux.scala 46:19:@13513.4]
  wire [7:0] _T_15187; // @[Mux.scala 46:16:@13514.4]
  wire  _T_15188; // @[Mux.scala 46:19:@13515.4]
  wire [7:0] _T_15189; // @[Mux.scala 46:16:@13516.4]
  wire  _T_15190; // @[Mux.scala 46:19:@13517.4]
  wire [7:0] _T_15191; // @[Mux.scala 46:16:@13518.4]
  wire  _T_15192; // @[Mux.scala 46:19:@13519.4]
  wire [7:0] _T_15193; // @[Mux.scala 46:16:@13520.4]
  wire  _T_15194; // @[Mux.scala 46:19:@13521.4]
  wire [7:0] _T_15195; // @[Mux.scala 46:16:@13522.4]
  wire  _T_15196; // @[Mux.scala 46:19:@13523.4]
  wire [7:0] _T_15197; // @[Mux.scala 46:16:@13524.4]
  wire  _T_15198; // @[Mux.scala 46:19:@13525.4]
  wire [7:0] _T_15199; // @[Mux.scala 46:16:@13526.4]
  wire  _T_15200; // @[Mux.scala 46:19:@13527.4]
  wire [7:0] _T_15201; // @[Mux.scala 46:16:@13528.4]
  wire  _T_15202; // @[Mux.scala 46:19:@13529.4]
  wire [7:0] _T_15203; // @[Mux.scala 46:16:@13530.4]
  wire  _T_15204; // @[Mux.scala 46:19:@13531.4]
  wire [7:0] _T_15205; // @[Mux.scala 46:16:@13532.4]
  wire  _T_15206; // @[Mux.scala 46:19:@13533.4]
  wire [7:0] _T_15207; // @[Mux.scala 46:16:@13534.4]
  wire  _T_15208; // @[Mux.scala 46:19:@13535.4]
  wire [7:0] _T_15209; // @[Mux.scala 46:16:@13536.4]
  wire  _T_15210; // @[Mux.scala 46:19:@13537.4]
  wire [7:0] _T_15211; // @[Mux.scala 46:16:@13538.4]
  wire  _T_15212; // @[Mux.scala 46:19:@13539.4]
  wire [7:0] _T_15213; // @[Mux.scala 46:16:@13540.4]
  wire  _T_15214; // @[Mux.scala 46:19:@13541.4]
  wire [7:0] _T_15215; // @[Mux.scala 46:16:@13542.4]
  wire  _T_15216; // @[Mux.scala 46:19:@13543.4]
  wire [7:0] _T_15217; // @[Mux.scala 46:16:@13544.4]
  wire  _T_15218; // @[Mux.scala 46:19:@13545.4]
  wire [7:0] _T_15219; // @[Mux.scala 46:16:@13546.4]
  wire  _T_15220; // @[Mux.scala 46:19:@13547.4]
  wire [7:0] _T_15221; // @[Mux.scala 46:16:@13548.4]
  wire  _T_15222; // @[Mux.scala 46:19:@13549.4]
  wire [7:0] _T_15223; // @[Mux.scala 46:16:@13550.4]
  wire  _T_15224; // @[Mux.scala 46:19:@13551.4]
  wire [7:0] _T_15225; // @[Mux.scala 46:16:@13552.4]
  wire  _T_15226; // @[Mux.scala 46:19:@13553.4]
  wire [7:0] _T_15227; // @[Mux.scala 46:16:@13554.4]
  wire  _T_15228; // @[Mux.scala 46:19:@13555.4]
  wire [7:0] _T_15229; // @[Mux.scala 46:16:@13556.4]
  wire  _T_15230; // @[Mux.scala 46:19:@13557.4]
  wire [7:0] _T_15231; // @[Mux.scala 46:16:@13558.4]
  wire  _T_15232; // @[Mux.scala 46:19:@13559.4]
  wire [7:0] _T_15233; // @[Mux.scala 46:16:@13560.4]
  wire  _T_15234; // @[Mux.scala 46:19:@13561.4]
  wire [7:0] _T_15235; // @[Mux.scala 46:16:@13562.4]
  wire  _T_15236; // @[Mux.scala 46:19:@13563.4]
  wire [7:0] _T_15237; // @[Mux.scala 46:16:@13564.4]
  wire  _T_15238; // @[Mux.scala 46:19:@13565.4]
  wire [7:0] _T_15239; // @[Mux.scala 46:16:@13566.4]
  wire  _T_15291; // @[Mux.scala 46:19:@13568.4]
  wire [7:0] _T_15292; // @[Mux.scala 46:16:@13569.4]
  wire  _T_15293; // @[Mux.scala 46:19:@13570.4]
  wire [7:0] _T_15294; // @[Mux.scala 46:16:@13571.4]
  wire  _T_15295; // @[Mux.scala 46:19:@13572.4]
  wire [7:0] _T_15296; // @[Mux.scala 46:16:@13573.4]
  wire  _T_15297; // @[Mux.scala 46:19:@13574.4]
  wire [7:0] _T_15298; // @[Mux.scala 46:16:@13575.4]
  wire  _T_15299; // @[Mux.scala 46:19:@13576.4]
  wire [7:0] _T_15300; // @[Mux.scala 46:16:@13577.4]
  wire  _T_15301; // @[Mux.scala 46:19:@13578.4]
  wire [7:0] _T_15302; // @[Mux.scala 46:16:@13579.4]
  wire  _T_15303; // @[Mux.scala 46:19:@13580.4]
  wire [7:0] _T_15304; // @[Mux.scala 46:16:@13581.4]
  wire  _T_15305; // @[Mux.scala 46:19:@13582.4]
  wire [7:0] _T_15306; // @[Mux.scala 46:16:@13583.4]
  wire  _T_15307; // @[Mux.scala 46:19:@13584.4]
  wire [7:0] _T_15308; // @[Mux.scala 46:16:@13585.4]
  wire  _T_15309; // @[Mux.scala 46:19:@13586.4]
  wire [7:0] _T_15310; // @[Mux.scala 46:16:@13587.4]
  wire  _T_15311; // @[Mux.scala 46:19:@13588.4]
  wire [7:0] _T_15312; // @[Mux.scala 46:16:@13589.4]
  wire  _T_15313; // @[Mux.scala 46:19:@13590.4]
  wire [7:0] _T_15314; // @[Mux.scala 46:16:@13591.4]
  wire  _T_15315; // @[Mux.scala 46:19:@13592.4]
  wire [7:0] _T_15316; // @[Mux.scala 46:16:@13593.4]
  wire  _T_15317; // @[Mux.scala 46:19:@13594.4]
  wire [7:0] _T_15318; // @[Mux.scala 46:16:@13595.4]
  wire  _T_15319; // @[Mux.scala 46:19:@13596.4]
  wire [7:0] _T_15320; // @[Mux.scala 46:16:@13597.4]
  wire  _T_15321; // @[Mux.scala 46:19:@13598.4]
  wire [7:0] _T_15322; // @[Mux.scala 46:16:@13599.4]
  wire  _T_15323; // @[Mux.scala 46:19:@13600.4]
  wire [7:0] _T_15324; // @[Mux.scala 46:16:@13601.4]
  wire  _T_15325; // @[Mux.scala 46:19:@13602.4]
  wire [7:0] _T_15326; // @[Mux.scala 46:16:@13603.4]
  wire  _T_15327; // @[Mux.scala 46:19:@13604.4]
  wire [7:0] _T_15328; // @[Mux.scala 46:16:@13605.4]
  wire  _T_15329; // @[Mux.scala 46:19:@13606.4]
  wire [7:0] _T_15330; // @[Mux.scala 46:16:@13607.4]
  wire  _T_15331; // @[Mux.scala 46:19:@13608.4]
  wire [7:0] _T_15332; // @[Mux.scala 46:16:@13609.4]
  wire  _T_15333; // @[Mux.scala 46:19:@13610.4]
  wire [7:0] _T_15334; // @[Mux.scala 46:16:@13611.4]
  wire  _T_15335; // @[Mux.scala 46:19:@13612.4]
  wire [7:0] _T_15336; // @[Mux.scala 46:16:@13613.4]
  wire  _T_15337; // @[Mux.scala 46:19:@13614.4]
  wire [7:0] _T_15338; // @[Mux.scala 46:16:@13615.4]
  wire  _T_15339; // @[Mux.scala 46:19:@13616.4]
  wire [7:0] _T_15340; // @[Mux.scala 46:16:@13617.4]
  wire  _T_15341; // @[Mux.scala 46:19:@13618.4]
  wire [7:0] _T_15342; // @[Mux.scala 46:16:@13619.4]
  wire  _T_15343; // @[Mux.scala 46:19:@13620.4]
  wire [7:0] _T_15344; // @[Mux.scala 46:16:@13621.4]
  wire  _T_15345; // @[Mux.scala 46:19:@13622.4]
  wire [7:0] _T_15346; // @[Mux.scala 46:16:@13623.4]
  wire  _T_15347; // @[Mux.scala 46:19:@13624.4]
  wire [7:0] _T_15348; // @[Mux.scala 46:16:@13625.4]
  wire  _T_15349; // @[Mux.scala 46:19:@13626.4]
  wire [7:0] _T_15350; // @[Mux.scala 46:16:@13627.4]
  wire  _T_15351; // @[Mux.scala 46:19:@13628.4]
  wire [7:0] _T_15352; // @[Mux.scala 46:16:@13629.4]
  wire  _T_15353; // @[Mux.scala 46:19:@13630.4]
  wire [7:0] _T_15354; // @[Mux.scala 46:16:@13631.4]
  wire  _T_15355; // @[Mux.scala 46:19:@13632.4]
  wire [7:0] _T_15356; // @[Mux.scala 46:16:@13633.4]
  wire  _T_15357; // @[Mux.scala 46:19:@13634.4]
  wire [7:0] _T_15358; // @[Mux.scala 46:16:@13635.4]
  wire  _T_15359; // @[Mux.scala 46:19:@13636.4]
  wire [7:0] _T_15360; // @[Mux.scala 46:16:@13637.4]
  wire  _T_15361; // @[Mux.scala 46:19:@13638.4]
  wire [7:0] _T_15362; // @[Mux.scala 46:16:@13639.4]
  wire  _T_15363; // @[Mux.scala 46:19:@13640.4]
  wire [7:0] _T_15364; // @[Mux.scala 46:16:@13641.4]
  wire  _T_15365; // @[Mux.scala 46:19:@13642.4]
  wire [7:0] _T_15366; // @[Mux.scala 46:16:@13643.4]
  wire  _T_15367; // @[Mux.scala 46:19:@13644.4]
  wire [7:0] _T_15368; // @[Mux.scala 46:16:@13645.4]
  wire  _T_15369; // @[Mux.scala 46:19:@13646.4]
  wire [7:0] _T_15370; // @[Mux.scala 46:16:@13647.4]
  wire  _T_15371; // @[Mux.scala 46:19:@13648.4]
  wire [7:0] _T_15372; // @[Mux.scala 46:16:@13649.4]
  wire  _T_15373; // @[Mux.scala 46:19:@13650.4]
  wire [7:0] _T_15374; // @[Mux.scala 46:16:@13651.4]
  wire  _T_15375; // @[Mux.scala 46:19:@13652.4]
  wire [7:0] _T_15376; // @[Mux.scala 46:16:@13653.4]
  wire  _T_15377; // @[Mux.scala 46:19:@13654.4]
  wire [7:0] _T_15378; // @[Mux.scala 46:16:@13655.4]
  wire  _T_15379; // @[Mux.scala 46:19:@13656.4]
  wire [7:0] _T_15380; // @[Mux.scala 46:16:@13657.4]
  wire  _T_15381; // @[Mux.scala 46:19:@13658.4]
  wire [7:0] _T_15382; // @[Mux.scala 46:16:@13659.4]
  wire  _T_15383; // @[Mux.scala 46:19:@13660.4]
  wire [7:0] _T_15384; // @[Mux.scala 46:16:@13661.4]
  wire  _T_15385; // @[Mux.scala 46:19:@13662.4]
  wire [7:0] _T_15386; // @[Mux.scala 46:16:@13663.4]
  wire  _T_15387; // @[Mux.scala 46:19:@13664.4]
  wire [7:0] _T_15388; // @[Mux.scala 46:16:@13665.4]
  wire  _T_15389; // @[Mux.scala 46:19:@13666.4]
  wire [7:0] _T_15390; // @[Mux.scala 46:16:@13667.4]
  wire  _T_15443; // @[Mux.scala 46:19:@13669.4]
  wire [7:0] _T_15444; // @[Mux.scala 46:16:@13670.4]
  wire  _T_15445; // @[Mux.scala 46:19:@13671.4]
  wire [7:0] _T_15446; // @[Mux.scala 46:16:@13672.4]
  wire  _T_15447; // @[Mux.scala 46:19:@13673.4]
  wire [7:0] _T_15448; // @[Mux.scala 46:16:@13674.4]
  wire  _T_15449; // @[Mux.scala 46:19:@13675.4]
  wire [7:0] _T_15450; // @[Mux.scala 46:16:@13676.4]
  wire  _T_15451; // @[Mux.scala 46:19:@13677.4]
  wire [7:0] _T_15452; // @[Mux.scala 46:16:@13678.4]
  wire  _T_15453; // @[Mux.scala 46:19:@13679.4]
  wire [7:0] _T_15454; // @[Mux.scala 46:16:@13680.4]
  wire  _T_15455; // @[Mux.scala 46:19:@13681.4]
  wire [7:0] _T_15456; // @[Mux.scala 46:16:@13682.4]
  wire  _T_15457; // @[Mux.scala 46:19:@13683.4]
  wire [7:0] _T_15458; // @[Mux.scala 46:16:@13684.4]
  wire  _T_15459; // @[Mux.scala 46:19:@13685.4]
  wire [7:0] _T_15460; // @[Mux.scala 46:16:@13686.4]
  wire  _T_15461; // @[Mux.scala 46:19:@13687.4]
  wire [7:0] _T_15462; // @[Mux.scala 46:16:@13688.4]
  wire  _T_15463; // @[Mux.scala 46:19:@13689.4]
  wire [7:0] _T_15464; // @[Mux.scala 46:16:@13690.4]
  wire  _T_15465; // @[Mux.scala 46:19:@13691.4]
  wire [7:0] _T_15466; // @[Mux.scala 46:16:@13692.4]
  wire  _T_15467; // @[Mux.scala 46:19:@13693.4]
  wire [7:0] _T_15468; // @[Mux.scala 46:16:@13694.4]
  wire  _T_15469; // @[Mux.scala 46:19:@13695.4]
  wire [7:0] _T_15470; // @[Mux.scala 46:16:@13696.4]
  wire  _T_15471; // @[Mux.scala 46:19:@13697.4]
  wire [7:0] _T_15472; // @[Mux.scala 46:16:@13698.4]
  wire  _T_15473; // @[Mux.scala 46:19:@13699.4]
  wire [7:0] _T_15474; // @[Mux.scala 46:16:@13700.4]
  wire  _T_15475; // @[Mux.scala 46:19:@13701.4]
  wire [7:0] _T_15476; // @[Mux.scala 46:16:@13702.4]
  wire  _T_15477; // @[Mux.scala 46:19:@13703.4]
  wire [7:0] _T_15478; // @[Mux.scala 46:16:@13704.4]
  wire  _T_15479; // @[Mux.scala 46:19:@13705.4]
  wire [7:0] _T_15480; // @[Mux.scala 46:16:@13706.4]
  wire  _T_15481; // @[Mux.scala 46:19:@13707.4]
  wire [7:0] _T_15482; // @[Mux.scala 46:16:@13708.4]
  wire  _T_15483; // @[Mux.scala 46:19:@13709.4]
  wire [7:0] _T_15484; // @[Mux.scala 46:16:@13710.4]
  wire  _T_15485; // @[Mux.scala 46:19:@13711.4]
  wire [7:0] _T_15486; // @[Mux.scala 46:16:@13712.4]
  wire  _T_15487; // @[Mux.scala 46:19:@13713.4]
  wire [7:0] _T_15488; // @[Mux.scala 46:16:@13714.4]
  wire  _T_15489; // @[Mux.scala 46:19:@13715.4]
  wire [7:0] _T_15490; // @[Mux.scala 46:16:@13716.4]
  wire  _T_15491; // @[Mux.scala 46:19:@13717.4]
  wire [7:0] _T_15492; // @[Mux.scala 46:16:@13718.4]
  wire  _T_15493; // @[Mux.scala 46:19:@13719.4]
  wire [7:0] _T_15494; // @[Mux.scala 46:16:@13720.4]
  wire  _T_15495; // @[Mux.scala 46:19:@13721.4]
  wire [7:0] _T_15496; // @[Mux.scala 46:16:@13722.4]
  wire  _T_15497; // @[Mux.scala 46:19:@13723.4]
  wire [7:0] _T_15498; // @[Mux.scala 46:16:@13724.4]
  wire  _T_15499; // @[Mux.scala 46:19:@13725.4]
  wire [7:0] _T_15500; // @[Mux.scala 46:16:@13726.4]
  wire  _T_15501; // @[Mux.scala 46:19:@13727.4]
  wire [7:0] _T_15502; // @[Mux.scala 46:16:@13728.4]
  wire  _T_15503; // @[Mux.scala 46:19:@13729.4]
  wire [7:0] _T_15504; // @[Mux.scala 46:16:@13730.4]
  wire  _T_15505; // @[Mux.scala 46:19:@13731.4]
  wire [7:0] _T_15506; // @[Mux.scala 46:16:@13732.4]
  wire  _T_15507; // @[Mux.scala 46:19:@13733.4]
  wire [7:0] _T_15508; // @[Mux.scala 46:16:@13734.4]
  wire  _T_15509; // @[Mux.scala 46:19:@13735.4]
  wire [7:0] _T_15510; // @[Mux.scala 46:16:@13736.4]
  wire  _T_15511; // @[Mux.scala 46:19:@13737.4]
  wire [7:0] _T_15512; // @[Mux.scala 46:16:@13738.4]
  wire  _T_15513; // @[Mux.scala 46:19:@13739.4]
  wire [7:0] _T_15514; // @[Mux.scala 46:16:@13740.4]
  wire  _T_15515; // @[Mux.scala 46:19:@13741.4]
  wire [7:0] _T_15516; // @[Mux.scala 46:16:@13742.4]
  wire  _T_15517; // @[Mux.scala 46:19:@13743.4]
  wire [7:0] _T_15518; // @[Mux.scala 46:16:@13744.4]
  wire  _T_15519; // @[Mux.scala 46:19:@13745.4]
  wire [7:0] _T_15520; // @[Mux.scala 46:16:@13746.4]
  wire  _T_15521; // @[Mux.scala 46:19:@13747.4]
  wire [7:0] _T_15522; // @[Mux.scala 46:16:@13748.4]
  wire  _T_15523; // @[Mux.scala 46:19:@13749.4]
  wire [7:0] _T_15524; // @[Mux.scala 46:16:@13750.4]
  wire  _T_15525; // @[Mux.scala 46:19:@13751.4]
  wire [7:0] _T_15526; // @[Mux.scala 46:16:@13752.4]
  wire  _T_15527; // @[Mux.scala 46:19:@13753.4]
  wire [7:0] _T_15528; // @[Mux.scala 46:16:@13754.4]
  wire  _T_15529; // @[Mux.scala 46:19:@13755.4]
  wire [7:0] _T_15530; // @[Mux.scala 46:16:@13756.4]
  wire  _T_15531; // @[Mux.scala 46:19:@13757.4]
  wire [7:0] _T_15532; // @[Mux.scala 46:16:@13758.4]
  wire  _T_15533; // @[Mux.scala 46:19:@13759.4]
  wire [7:0] _T_15534; // @[Mux.scala 46:16:@13760.4]
  wire  _T_15535; // @[Mux.scala 46:19:@13761.4]
  wire [7:0] _T_15536; // @[Mux.scala 46:16:@13762.4]
  wire  _T_15537; // @[Mux.scala 46:19:@13763.4]
  wire [7:0] _T_15538; // @[Mux.scala 46:16:@13764.4]
  wire  _T_15539; // @[Mux.scala 46:19:@13765.4]
  wire [7:0] _T_15540; // @[Mux.scala 46:16:@13766.4]
  wire  _T_15541; // @[Mux.scala 46:19:@13767.4]
  wire [7:0] _T_15542; // @[Mux.scala 46:16:@13768.4]
  wire  _T_15543; // @[Mux.scala 46:19:@13769.4]
  wire [7:0] _T_15544; // @[Mux.scala 46:16:@13770.4]
  wire  _T_15598; // @[Mux.scala 46:19:@13772.4]
  wire [7:0] _T_15599; // @[Mux.scala 46:16:@13773.4]
  wire  _T_15600; // @[Mux.scala 46:19:@13774.4]
  wire [7:0] _T_15601; // @[Mux.scala 46:16:@13775.4]
  wire  _T_15602; // @[Mux.scala 46:19:@13776.4]
  wire [7:0] _T_15603; // @[Mux.scala 46:16:@13777.4]
  wire  _T_15604; // @[Mux.scala 46:19:@13778.4]
  wire [7:0] _T_15605; // @[Mux.scala 46:16:@13779.4]
  wire  _T_15606; // @[Mux.scala 46:19:@13780.4]
  wire [7:0] _T_15607; // @[Mux.scala 46:16:@13781.4]
  wire  _T_15608; // @[Mux.scala 46:19:@13782.4]
  wire [7:0] _T_15609; // @[Mux.scala 46:16:@13783.4]
  wire  _T_15610; // @[Mux.scala 46:19:@13784.4]
  wire [7:0] _T_15611; // @[Mux.scala 46:16:@13785.4]
  wire  _T_15612; // @[Mux.scala 46:19:@13786.4]
  wire [7:0] _T_15613; // @[Mux.scala 46:16:@13787.4]
  wire  _T_15614; // @[Mux.scala 46:19:@13788.4]
  wire [7:0] _T_15615; // @[Mux.scala 46:16:@13789.4]
  wire  _T_15616; // @[Mux.scala 46:19:@13790.4]
  wire [7:0] _T_15617; // @[Mux.scala 46:16:@13791.4]
  wire  _T_15618; // @[Mux.scala 46:19:@13792.4]
  wire [7:0] _T_15619; // @[Mux.scala 46:16:@13793.4]
  wire  _T_15620; // @[Mux.scala 46:19:@13794.4]
  wire [7:0] _T_15621; // @[Mux.scala 46:16:@13795.4]
  wire  _T_15622; // @[Mux.scala 46:19:@13796.4]
  wire [7:0] _T_15623; // @[Mux.scala 46:16:@13797.4]
  wire  _T_15624; // @[Mux.scala 46:19:@13798.4]
  wire [7:0] _T_15625; // @[Mux.scala 46:16:@13799.4]
  wire  _T_15626; // @[Mux.scala 46:19:@13800.4]
  wire [7:0] _T_15627; // @[Mux.scala 46:16:@13801.4]
  wire  _T_15628; // @[Mux.scala 46:19:@13802.4]
  wire [7:0] _T_15629; // @[Mux.scala 46:16:@13803.4]
  wire  _T_15630; // @[Mux.scala 46:19:@13804.4]
  wire [7:0] _T_15631; // @[Mux.scala 46:16:@13805.4]
  wire  _T_15632; // @[Mux.scala 46:19:@13806.4]
  wire [7:0] _T_15633; // @[Mux.scala 46:16:@13807.4]
  wire  _T_15634; // @[Mux.scala 46:19:@13808.4]
  wire [7:0] _T_15635; // @[Mux.scala 46:16:@13809.4]
  wire  _T_15636; // @[Mux.scala 46:19:@13810.4]
  wire [7:0] _T_15637; // @[Mux.scala 46:16:@13811.4]
  wire  _T_15638; // @[Mux.scala 46:19:@13812.4]
  wire [7:0] _T_15639; // @[Mux.scala 46:16:@13813.4]
  wire  _T_15640; // @[Mux.scala 46:19:@13814.4]
  wire [7:0] _T_15641; // @[Mux.scala 46:16:@13815.4]
  wire  _T_15642; // @[Mux.scala 46:19:@13816.4]
  wire [7:0] _T_15643; // @[Mux.scala 46:16:@13817.4]
  wire  _T_15644; // @[Mux.scala 46:19:@13818.4]
  wire [7:0] _T_15645; // @[Mux.scala 46:16:@13819.4]
  wire  _T_15646; // @[Mux.scala 46:19:@13820.4]
  wire [7:0] _T_15647; // @[Mux.scala 46:16:@13821.4]
  wire  _T_15648; // @[Mux.scala 46:19:@13822.4]
  wire [7:0] _T_15649; // @[Mux.scala 46:16:@13823.4]
  wire  _T_15650; // @[Mux.scala 46:19:@13824.4]
  wire [7:0] _T_15651; // @[Mux.scala 46:16:@13825.4]
  wire  _T_15652; // @[Mux.scala 46:19:@13826.4]
  wire [7:0] _T_15653; // @[Mux.scala 46:16:@13827.4]
  wire  _T_15654; // @[Mux.scala 46:19:@13828.4]
  wire [7:0] _T_15655; // @[Mux.scala 46:16:@13829.4]
  wire  _T_15656; // @[Mux.scala 46:19:@13830.4]
  wire [7:0] _T_15657; // @[Mux.scala 46:16:@13831.4]
  wire  _T_15658; // @[Mux.scala 46:19:@13832.4]
  wire [7:0] _T_15659; // @[Mux.scala 46:16:@13833.4]
  wire  _T_15660; // @[Mux.scala 46:19:@13834.4]
  wire [7:0] _T_15661; // @[Mux.scala 46:16:@13835.4]
  wire  _T_15662; // @[Mux.scala 46:19:@13836.4]
  wire [7:0] _T_15663; // @[Mux.scala 46:16:@13837.4]
  wire  _T_15664; // @[Mux.scala 46:19:@13838.4]
  wire [7:0] _T_15665; // @[Mux.scala 46:16:@13839.4]
  wire  _T_15666; // @[Mux.scala 46:19:@13840.4]
  wire [7:0] _T_15667; // @[Mux.scala 46:16:@13841.4]
  wire  _T_15668; // @[Mux.scala 46:19:@13842.4]
  wire [7:0] _T_15669; // @[Mux.scala 46:16:@13843.4]
  wire  _T_15670; // @[Mux.scala 46:19:@13844.4]
  wire [7:0] _T_15671; // @[Mux.scala 46:16:@13845.4]
  wire  _T_15672; // @[Mux.scala 46:19:@13846.4]
  wire [7:0] _T_15673; // @[Mux.scala 46:16:@13847.4]
  wire  _T_15674; // @[Mux.scala 46:19:@13848.4]
  wire [7:0] _T_15675; // @[Mux.scala 46:16:@13849.4]
  wire  _T_15676; // @[Mux.scala 46:19:@13850.4]
  wire [7:0] _T_15677; // @[Mux.scala 46:16:@13851.4]
  wire  _T_15678; // @[Mux.scala 46:19:@13852.4]
  wire [7:0] _T_15679; // @[Mux.scala 46:16:@13853.4]
  wire  _T_15680; // @[Mux.scala 46:19:@13854.4]
  wire [7:0] _T_15681; // @[Mux.scala 46:16:@13855.4]
  wire  _T_15682; // @[Mux.scala 46:19:@13856.4]
  wire [7:0] _T_15683; // @[Mux.scala 46:16:@13857.4]
  wire  _T_15684; // @[Mux.scala 46:19:@13858.4]
  wire [7:0] _T_15685; // @[Mux.scala 46:16:@13859.4]
  wire  _T_15686; // @[Mux.scala 46:19:@13860.4]
  wire [7:0] _T_15687; // @[Mux.scala 46:16:@13861.4]
  wire  _T_15688; // @[Mux.scala 46:19:@13862.4]
  wire [7:0] _T_15689; // @[Mux.scala 46:16:@13863.4]
  wire  _T_15690; // @[Mux.scala 46:19:@13864.4]
  wire [7:0] _T_15691; // @[Mux.scala 46:16:@13865.4]
  wire  _T_15692; // @[Mux.scala 46:19:@13866.4]
  wire [7:0] _T_15693; // @[Mux.scala 46:16:@13867.4]
  wire  _T_15694; // @[Mux.scala 46:19:@13868.4]
  wire [7:0] _T_15695; // @[Mux.scala 46:16:@13869.4]
  wire  _T_15696; // @[Mux.scala 46:19:@13870.4]
  wire [7:0] _T_15697; // @[Mux.scala 46:16:@13871.4]
  wire  _T_15698; // @[Mux.scala 46:19:@13872.4]
  wire [7:0] _T_15699; // @[Mux.scala 46:16:@13873.4]
  wire  _T_15700; // @[Mux.scala 46:19:@13874.4]
  wire [7:0] _T_15701; // @[Mux.scala 46:16:@13875.4]
  wire  _T_15756; // @[Mux.scala 46:19:@13877.4]
  wire [7:0] _T_15757; // @[Mux.scala 46:16:@13878.4]
  wire  _T_15758; // @[Mux.scala 46:19:@13879.4]
  wire [7:0] _T_15759; // @[Mux.scala 46:16:@13880.4]
  wire  _T_15760; // @[Mux.scala 46:19:@13881.4]
  wire [7:0] _T_15761; // @[Mux.scala 46:16:@13882.4]
  wire  _T_15762; // @[Mux.scala 46:19:@13883.4]
  wire [7:0] _T_15763; // @[Mux.scala 46:16:@13884.4]
  wire  _T_15764; // @[Mux.scala 46:19:@13885.4]
  wire [7:0] _T_15765; // @[Mux.scala 46:16:@13886.4]
  wire  _T_15766; // @[Mux.scala 46:19:@13887.4]
  wire [7:0] _T_15767; // @[Mux.scala 46:16:@13888.4]
  wire  _T_15768; // @[Mux.scala 46:19:@13889.4]
  wire [7:0] _T_15769; // @[Mux.scala 46:16:@13890.4]
  wire  _T_15770; // @[Mux.scala 46:19:@13891.4]
  wire [7:0] _T_15771; // @[Mux.scala 46:16:@13892.4]
  wire  _T_15772; // @[Mux.scala 46:19:@13893.4]
  wire [7:0] _T_15773; // @[Mux.scala 46:16:@13894.4]
  wire  _T_15774; // @[Mux.scala 46:19:@13895.4]
  wire [7:0] _T_15775; // @[Mux.scala 46:16:@13896.4]
  wire  _T_15776; // @[Mux.scala 46:19:@13897.4]
  wire [7:0] _T_15777; // @[Mux.scala 46:16:@13898.4]
  wire  _T_15778; // @[Mux.scala 46:19:@13899.4]
  wire [7:0] _T_15779; // @[Mux.scala 46:16:@13900.4]
  wire  _T_15780; // @[Mux.scala 46:19:@13901.4]
  wire [7:0] _T_15781; // @[Mux.scala 46:16:@13902.4]
  wire  _T_15782; // @[Mux.scala 46:19:@13903.4]
  wire [7:0] _T_15783; // @[Mux.scala 46:16:@13904.4]
  wire  _T_15784; // @[Mux.scala 46:19:@13905.4]
  wire [7:0] _T_15785; // @[Mux.scala 46:16:@13906.4]
  wire  _T_15786; // @[Mux.scala 46:19:@13907.4]
  wire [7:0] _T_15787; // @[Mux.scala 46:16:@13908.4]
  wire  _T_15788; // @[Mux.scala 46:19:@13909.4]
  wire [7:0] _T_15789; // @[Mux.scala 46:16:@13910.4]
  wire  _T_15790; // @[Mux.scala 46:19:@13911.4]
  wire [7:0] _T_15791; // @[Mux.scala 46:16:@13912.4]
  wire  _T_15792; // @[Mux.scala 46:19:@13913.4]
  wire [7:0] _T_15793; // @[Mux.scala 46:16:@13914.4]
  wire  _T_15794; // @[Mux.scala 46:19:@13915.4]
  wire [7:0] _T_15795; // @[Mux.scala 46:16:@13916.4]
  wire  _T_15796; // @[Mux.scala 46:19:@13917.4]
  wire [7:0] _T_15797; // @[Mux.scala 46:16:@13918.4]
  wire  _T_15798; // @[Mux.scala 46:19:@13919.4]
  wire [7:0] _T_15799; // @[Mux.scala 46:16:@13920.4]
  wire  _T_15800; // @[Mux.scala 46:19:@13921.4]
  wire [7:0] _T_15801; // @[Mux.scala 46:16:@13922.4]
  wire  _T_15802; // @[Mux.scala 46:19:@13923.4]
  wire [7:0] _T_15803; // @[Mux.scala 46:16:@13924.4]
  wire  _T_15804; // @[Mux.scala 46:19:@13925.4]
  wire [7:0] _T_15805; // @[Mux.scala 46:16:@13926.4]
  wire  _T_15806; // @[Mux.scala 46:19:@13927.4]
  wire [7:0] _T_15807; // @[Mux.scala 46:16:@13928.4]
  wire  _T_15808; // @[Mux.scala 46:19:@13929.4]
  wire [7:0] _T_15809; // @[Mux.scala 46:16:@13930.4]
  wire  _T_15810; // @[Mux.scala 46:19:@13931.4]
  wire [7:0] _T_15811; // @[Mux.scala 46:16:@13932.4]
  wire  _T_15812; // @[Mux.scala 46:19:@13933.4]
  wire [7:0] _T_15813; // @[Mux.scala 46:16:@13934.4]
  wire  _T_15814; // @[Mux.scala 46:19:@13935.4]
  wire [7:0] _T_15815; // @[Mux.scala 46:16:@13936.4]
  wire  _T_15816; // @[Mux.scala 46:19:@13937.4]
  wire [7:0] _T_15817; // @[Mux.scala 46:16:@13938.4]
  wire  _T_15818; // @[Mux.scala 46:19:@13939.4]
  wire [7:0] _T_15819; // @[Mux.scala 46:16:@13940.4]
  wire  _T_15820; // @[Mux.scala 46:19:@13941.4]
  wire [7:0] _T_15821; // @[Mux.scala 46:16:@13942.4]
  wire  _T_15822; // @[Mux.scala 46:19:@13943.4]
  wire [7:0] _T_15823; // @[Mux.scala 46:16:@13944.4]
  wire  _T_15824; // @[Mux.scala 46:19:@13945.4]
  wire [7:0] _T_15825; // @[Mux.scala 46:16:@13946.4]
  wire  _T_15826; // @[Mux.scala 46:19:@13947.4]
  wire [7:0] _T_15827; // @[Mux.scala 46:16:@13948.4]
  wire  _T_15828; // @[Mux.scala 46:19:@13949.4]
  wire [7:0] _T_15829; // @[Mux.scala 46:16:@13950.4]
  wire  _T_15830; // @[Mux.scala 46:19:@13951.4]
  wire [7:0] _T_15831; // @[Mux.scala 46:16:@13952.4]
  wire  _T_15832; // @[Mux.scala 46:19:@13953.4]
  wire [7:0] _T_15833; // @[Mux.scala 46:16:@13954.4]
  wire  _T_15834; // @[Mux.scala 46:19:@13955.4]
  wire [7:0] _T_15835; // @[Mux.scala 46:16:@13956.4]
  wire  _T_15836; // @[Mux.scala 46:19:@13957.4]
  wire [7:0] _T_15837; // @[Mux.scala 46:16:@13958.4]
  wire  _T_15838; // @[Mux.scala 46:19:@13959.4]
  wire [7:0] _T_15839; // @[Mux.scala 46:16:@13960.4]
  wire  _T_15840; // @[Mux.scala 46:19:@13961.4]
  wire [7:0] _T_15841; // @[Mux.scala 46:16:@13962.4]
  wire  _T_15842; // @[Mux.scala 46:19:@13963.4]
  wire [7:0] _T_15843; // @[Mux.scala 46:16:@13964.4]
  wire  _T_15844; // @[Mux.scala 46:19:@13965.4]
  wire [7:0] _T_15845; // @[Mux.scala 46:16:@13966.4]
  wire  _T_15846; // @[Mux.scala 46:19:@13967.4]
  wire [7:0] _T_15847; // @[Mux.scala 46:16:@13968.4]
  wire  _T_15848; // @[Mux.scala 46:19:@13969.4]
  wire [7:0] _T_15849; // @[Mux.scala 46:16:@13970.4]
  wire  _T_15850; // @[Mux.scala 46:19:@13971.4]
  wire [7:0] _T_15851; // @[Mux.scala 46:16:@13972.4]
  wire  _T_15852; // @[Mux.scala 46:19:@13973.4]
  wire [7:0] _T_15853; // @[Mux.scala 46:16:@13974.4]
  wire  _T_15854; // @[Mux.scala 46:19:@13975.4]
  wire [7:0] _T_15855; // @[Mux.scala 46:16:@13976.4]
  wire  _T_15856; // @[Mux.scala 46:19:@13977.4]
  wire [7:0] _T_15857; // @[Mux.scala 46:16:@13978.4]
  wire  _T_15858; // @[Mux.scala 46:19:@13979.4]
  wire [7:0] _T_15859; // @[Mux.scala 46:16:@13980.4]
  wire  _T_15860; // @[Mux.scala 46:19:@13981.4]
  wire [7:0] _T_15861; // @[Mux.scala 46:16:@13982.4]
  wire  _T_15917; // @[Mux.scala 46:19:@13984.4]
  wire [7:0] _T_15918; // @[Mux.scala 46:16:@13985.4]
  wire  _T_15919; // @[Mux.scala 46:19:@13986.4]
  wire [7:0] _T_15920; // @[Mux.scala 46:16:@13987.4]
  wire  _T_15921; // @[Mux.scala 46:19:@13988.4]
  wire [7:0] _T_15922; // @[Mux.scala 46:16:@13989.4]
  wire  _T_15923; // @[Mux.scala 46:19:@13990.4]
  wire [7:0] _T_15924; // @[Mux.scala 46:16:@13991.4]
  wire  _T_15925; // @[Mux.scala 46:19:@13992.4]
  wire [7:0] _T_15926; // @[Mux.scala 46:16:@13993.4]
  wire  _T_15927; // @[Mux.scala 46:19:@13994.4]
  wire [7:0] _T_15928; // @[Mux.scala 46:16:@13995.4]
  wire  _T_15929; // @[Mux.scala 46:19:@13996.4]
  wire [7:0] _T_15930; // @[Mux.scala 46:16:@13997.4]
  wire  _T_15931; // @[Mux.scala 46:19:@13998.4]
  wire [7:0] _T_15932; // @[Mux.scala 46:16:@13999.4]
  wire  _T_15933; // @[Mux.scala 46:19:@14000.4]
  wire [7:0] _T_15934; // @[Mux.scala 46:16:@14001.4]
  wire  _T_15935; // @[Mux.scala 46:19:@14002.4]
  wire [7:0] _T_15936; // @[Mux.scala 46:16:@14003.4]
  wire  _T_15937; // @[Mux.scala 46:19:@14004.4]
  wire [7:0] _T_15938; // @[Mux.scala 46:16:@14005.4]
  wire  _T_15939; // @[Mux.scala 46:19:@14006.4]
  wire [7:0] _T_15940; // @[Mux.scala 46:16:@14007.4]
  wire  _T_15941; // @[Mux.scala 46:19:@14008.4]
  wire [7:0] _T_15942; // @[Mux.scala 46:16:@14009.4]
  wire  _T_15943; // @[Mux.scala 46:19:@14010.4]
  wire [7:0] _T_15944; // @[Mux.scala 46:16:@14011.4]
  wire  _T_15945; // @[Mux.scala 46:19:@14012.4]
  wire [7:0] _T_15946; // @[Mux.scala 46:16:@14013.4]
  wire  _T_15947; // @[Mux.scala 46:19:@14014.4]
  wire [7:0] _T_15948; // @[Mux.scala 46:16:@14015.4]
  wire  _T_15949; // @[Mux.scala 46:19:@14016.4]
  wire [7:0] _T_15950; // @[Mux.scala 46:16:@14017.4]
  wire  _T_15951; // @[Mux.scala 46:19:@14018.4]
  wire [7:0] _T_15952; // @[Mux.scala 46:16:@14019.4]
  wire  _T_15953; // @[Mux.scala 46:19:@14020.4]
  wire [7:0] _T_15954; // @[Mux.scala 46:16:@14021.4]
  wire  _T_15955; // @[Mux.scala 46:19:@14022.4]
  wire [7:0] _T_15956; // @[Mux.scala 46:16:@14023.4]
  wire  _T_15957; // @[Mux.scala 46:19:@14024.4]
  wire [7:0] _T_15958; // @[Mux.scala 46:16:@14025.4]
  wire  _T_15959; // @[Mux.scala 46:19:@14026.4]
  wire [7:0] _T_15960; // @[Mux.scala 46:16:@14027.4]
  wire  _T_15961; // @[Mux.scala 46:19:@14028.4]
  wire [7:0] _T_15962; // @[Mux.scala 46:16:@14029.4]
  wire  _T_15963; // @[Mux.scala 46:19:@14030.4]
  wire [7:0] _T_15964; // @[Mux.scala 46:16:@14031.4]
  wire  _T_15965; // @[Mux.scala 46:19:@14032.4]
  wire [7:0] _T_15966; // @[Mux.scala 46:16:@14033.4]
  wire  _T_15967; // @[Mux.scala 46:19:@14034.4]
  wire [7:0] _T_15968; // @[Mux.scala 46:16:@14035.4]
  wire  _T_15969; // @[Mux.scala 46:19:@14036.4]
  wire [7:0] _T_15970; // @[Mux.scala 46:16:@14037.4]
  wire  _T_15971; // @[Mux.scala 46:19:@14038.4]
  wire [7:0] _T_15972; // @[Mux.scala 46:16:@14039.4]
  wire  _T_15973; // @[Mux.scala 46:19:@14040.4]
  wire [7:0] _T_15974; // @[Mux.scala 46:16:@14041.4]
  wire  _T_15975; // @[Mux.scala 46:19:@14042.4]
  wire [7:0] _T_15976; // @[Mux.scala 46:16:@14043.4]
  wire  _T_15977; // @[Mux.scala 46:19:@14044.4]
  wire [7:0] _T_15978; // @[Mux.scala 46:16:@14045.4]
  wire  _T_15979; // @[Mux.scala 46:19:@14046.4]
  wire [7:0] _T_15980; // @[Mux.scala 46:16:@14047.4]
  wire  _T_15981; // @[Mux.scala 46:19:@14048.4]
  wire [7:0] _T_15982; // @[Mux.scala 46:16:@14049.4]
  wire  _T_15983; // @[Mux.scala 46:19:@14050.4]
  wire [7:0] _T_15984; // @[Mux.scala 46:16:@14051.4]
  wire  _T_15985; // @[Mux.scala 46:19:@14052.4]
  wire [7:0] _T_15986; // @[Mux.scala 46:16:@14053.4]
  wire  _T_15987; // @[Mux.scala 46:19:@14054.4]
  wire [7:0] _T_15988; // @[Mux.scala 46:16:@14055.4]
  wire  _T_15989; // @[Mux.scala 46:19:@14056.4]
  wire [7:0] _T_15990; // @[Mux.scala 46:16:@14057.4]
  wire  _T_15991; // @[Mux.scala 46:19:@14058.4]
  wire [7:0] _T_15992; // @[Mux.scala 46:16:@14059.4]
  wire  _T_15993; // @[Mux.scala 46:19:@14060.4]
  wire [7:0] _T_15994; // @[Mux.scala 46:16:@14061.4]
  wire  _T_15995; // @[Mux.scala 46:19:@14062.4]
  wire [7:0] _T_15996; // @[Mux.scala 46:16:@14063.4]
  wire  _T_15997; // @[Mux.scala 46:19:@14064.4]
  wire [7:0] _T_15998; // @[Mux.scala 46:16:@14065.4]
  wire  _T_15999; // @[Mux.scala 46:19:@14066.4]
  wire [7:0] _T_16000; // @[Mux.scala 46:16:@14067.4]
  wire  _T_16001; // @[Mux.scala 46:19:@14068.4]
  wire [7:0] _T_16002; // @[Mux.scala 46:16:@14069.4]
  wire  _T_16003; // @[Mux.scala 46:19:@14070.4]
  wire [7:0] _T_16004; // @[Mux.scala 46:16:@14071.4]
  wire  _T_16005; // @[Mux.scala 46:19:@14072.4]
  wire [7:0] _T_16006; // @[Mux.scala 46:16:@14073.4]
  wire  _T_16007; // @[Mux.scala 46:19:@14074.4]
  wire [7:0] _T_16008; // @[Mux.scala 46:16:@14075.4]
  wire  _T_16009; // @[Mux.scala 46:19:@14076.4]
  wire [7:0] _T_16010; // @[Mux.scala 46:16:@14077.4]
  wire  _T_16011; // @[Mux.scala 46:19:@14078.4]
  wire [7:0] _T_16012; // @[Mux.scala 46:16:@14079.4]
  wire  _T_16013; // @[Mux.scala 46:19:@14080.4]
  wire [7:0] _T_16014; // @[Mux.scala 46:16:@14081.4]
  wire  _T_16015; // @[Mux.scala 46:19:@14082.4]
  wire [7:0] _T_16016; // @[Mux.scala 46:16:@14083.4]
  wire  _T_16017; // @[Mux.scala 46:19:@14084.4]
  wire [7:0] _T_16018; // @[Mux.scala 46:16:@14085.4]
  wire  _T_16019; // @[Mux.scala 46:19:@14086.4]
  wire [7:0] _T_16020; // @[Mux.scala 46:16:@14087.4]
  wire  _T_16021; // @[Mux.scala 46:19:@14088.4]
  wire [7:0] _T_16022; // @[Mux.scala 46:16:@14089.4]
  wire  _T_16023; // @[Mux.scala 46:19:@14090.4]
  wire [7:0] _T_16024; // @[Mux.scala 46:16:@14091.4]
  wire  _T_16081; // @[Mux.scala 46:19:@14093.4]
  wire [7:0] _T_16082; // @[Mux.scala 46:16:@14094.4]
  wire  _T_16083; // @[Mux.scala 46:19:@14095.4]
  wire [7:0] _T_16084; // @[Mux.scala 46:16:@14096.4]
  wire  _T_16085; // @[Mux.scala 46:19:@14097.4]
  wire [7:0] _T_16086; // @[Mux.scala 46:16:@14098.4]
  wire  _T_16087; // @[Mux.scala 46:19:@14099.4]
  wire [7:0] _T_16088; // @[Mux.scala 46:16:@14100.4]
  wire  _T_16089; // @[Mux.scala 46:19:@14101.4]
  wire [7:0] _T_16090; // @[Mux.scala 46:16:@14102.4]
  wire  _T_16091; // @[Mux.scala 46:19:@14103.4]
  wire [7:0] _T_16092; // @[Mux.scala 46:16:@14104.4]
  wire  _T_16093; // @[Mux.scala 46:19:@14105.4]
  wire [7:0] _T_16094; // @[Mux.scala 46:16:@14106.4]
  wire  _T_16095; // @[Mux.scala 46:19:@14107.4]
  wire [7:0] _T_16096; // @[Mux.scala 46:16:@14108.4]
  wire  _T_16097; // @[Mux.scala 46:19:@14109.4]
  wire [7:0] _T_16098; // @[Mux.scala 46:16:@14110.4]
  wire  _T_16099; // @[Mux.scala 46:19:@14111.4]
  wire [7:0] _T_16100; // @[Mux.scala 46:16:@14112.4]
  wire  _T_16101; // @[Mux.scala 46:19:@14113.4]
  wire [7:0] _T_16102; // @[Mux.scala 46:16:@14114.4]
  wire  _T_16103; // @[Mux.scala 46:19:@14115.4]
  wire [7:0] _T_16104; // @[Mux.scala 46:16:@14116.4]
  wire  _T_16105; // @[Mux.scala 46:19:@14117.4]
  wire [7:0] _T_16106; // @[Mux.scala 46:16:@14118.4]
  wire  _T_16107; // @[Mux.scala 46:19:@14119.4]
  wire [7:0] _T_16108; // @[Mux.scala 46:16:@14120.4]
  wire  _T_16109; // @[Mux.scala 46:19:@14121.4]
  wire [7:0] _T_16110; // @[Mux.scala 46:16:@14122.4]
  wire  _T_16111; // @[Mux.scala 46:19:@14123.4]
  wire [7:0] _T_16112; // @[Mux.scala 46:16:@14124.4]
  wire  _T_16113; // @[Mux.scala 46:19:@14125.4]
  wire [7:0] _T_16114; // @[Mux.scala 46:16:@14126.4]
  wire  _T_16115; // @[Mux.scala 46:19:@14127.4]
  wire [7:0] _T_16116; // @[Mux.scala 46:16:@14128.4]
  wire  _T_16117; // @[Mux.scala 46:19:@14129.4]
  wire [7:0] _T_16118; // @[Mux.scala 46:16:@14130.4]
  wire  _T_16119; // @[Mux.scala 46:19:@14131.4]
  wire [7:0] _T_16120; // @[Mux.scala 46:16:@14132.4]
  wire  _T_16121; // @[Mux.scala 46:19:@14133.4]
  wire [7:0] _T_16122; // @[Mux.scala 46:16:@14134.4]
  wire  _T_16123; // @[Mux.scala 46:19:@14135.4]
  wire [7:0] _T_16124; // @[Mux.scala 46:16:@14136.4]
  wire  _T_16125; // @[Mux.scala 46:19:@14137.4]
  wire [7:0] _T_16126; // @[Mux.scala 46:16:@14138.4]
  wire  _T_16127; // @[Mux.scala 46:19:@14139.4]
  wire [7:0] _T_16128; // @[Mux.scala 46:16:@14140.4]
  wire  _T_16129; // @[Mux.scala 46:19:@14141.4]
  wire [7:0] _T_16130; // @[Mux.scala 46:16:@14142.4]
  wire  _T_16131; // @[Mux.scala 46:19:@14143.4]
  wire [7:0] _T_16132; // @[Mux.scala 46:16:@14144.4]
  wire  _T_16133; // @[Mux.scala 46:19:@14145.4]
  wire [7:0] _T_16134; // @[Mux.scala 46:16:@14146.4]
  wire  _T_16135; // @[Mux.scala 46:19:@14147.4]
  wire [7:0] _T_16136; // @[Mux.scala 46:16:@14148.4]
  wire  _T_16137; // @[Mux.scala 46:19:@14149.4]
  wire [7:0] _T_16138; // @[Mux.scala 46:16:@14150.4]
  wire  _T_16139; // @[Mux.scala 46:19:@14151.4]
  wire [7:0] _T_16140; // @[Mux.scala 46:16:@14152.4]
  wire  _T_16141; // @[Mux.scala 46:19:@14153.4]
  wire [7:0] _T_16142; // @[Mux.scala 46:16:@14154.4]
  wire  _T_16143; // @[Mux.scala 46:19:@14155.4]
  wire [7:0] _T_16144; // @[Mux.scala 46:16:@14156.4]
  wire  _T_16145; // @[Mux.scala 46:19:@14157.4]
  wire [7:0] _T_16146; // @[Mux.scala 46:16:@14158.4]
  wire  _T_16147; // @[Mux.scala 46:19:@14159.4]
  wire [7:0] _T_16148; // @[Mux.scala 46:16:@14160.4]
  wire  _T_16149; // @[Mux.scala 46:19:@14161.4]
  wire [7:0] _T_16150; // @[Mux.scala 46:16:@14162.4]
  wire  _T_16151; // @[Mux.scala 46:19:@14163.4]
  wire [7:0] _T_16152; // @[Mux.scala 46:16:@14164.4]
  wire  _T_16153; // @[Mux.scala 46:19:@14165.4]
  wire [7:0] _T_16154; // @[Mux.scala 46:16:@14166.4]
  wire  _T_16155; // @[Mux.scala 46:19:@14167.4]
  wire [7:0] _T_16156; // @[Mux.scala 46:16:@14168.4]
  wire  _T_16157; // @[Mux.scala 46:19:@14169.4]
  wire [7:0] _T_16158; // @[Mux.scala 46:16:@14170.4]
  wire  _T_16159; // @[Mux.scala 46:19:@14171.4]
  wire [7:0] _T_16160; // @[Mux.scala 46:16:@14172.4]
  wire  _T_16161; // @[Mux.scala 46:19:@14173.4]
  wire [7:0] _T_16162; // @[Mux.scala 46:16:@14174.4]
  wire  _T_16163; // @[Mux.scala 46:19:@14175.4]
  wire [7:0] _T_16164; // @[Mux.scala 46:16:@14176.4]
  wire  _T_16165; // @[Mux.scala 46:19:@14177.4]
  wire [7:0] _T_16166; // @[Mux.scala 46:16:@14178.4]
  wire  _T_16167; // @[Mux.scala 46:19:@14179.4]
  wire [7:0] _T_16168; // @[Mux.scala 46:16:@14180.4]
  wire  _T_16169; // @[Mux.scala 46:19:@14181.4]
  wire [7:0] _T_16170; // @[Mux.scala 46:16:@14182.4]
  wire  _T_16171; // @[Mux.scala 46:19:@14183.4]
  wire [7:0] _T_16172; // @[Mux.scala 46:16:@14184.4]
  wire  _T_16173; // @[Mux.scala 46:19:@14185.4]
  wire [7:0] _T_16174; // @[Mux.scala 46:16:@14186.4]
  wire  _T_16175; // @[Mux.scala 46:19:@14187.4]
  wire [7:0] _T_16176; // @[Mux.scala 46:16:@14188.4]
  wire  _T_16177; // @[Mux.scala 46:19:@14189.4]
  wire [7:0] _T_16178; // @[Mux.scala 46:16:@14190.4]
  wire  _T_16179; // @[Mux.scala 46:19:@14191.4]
  wire [7:0] _T_16180; // @[Mux.scala 46:16:@14192.4]
  wire  _T_16181; // @[Mux.scala 46:19:@14193.4]
  wire [7:0] _T_16182; // @[Mux.scala 46:16:@14194.4]
  wire  _T_16183; // @[Mux.scala 46:19:@14195.4]
  wire [7:0] _T_16184; // @[Mux.scala 46:16:@14196.4]
  wire  _T_16185; // @[Mux.scala 46:19:@14197.4]
  wire [7:0] _T_16186; // @[Mux.scala 46:16:@14198.4]
  wire  _T_16187; // @[Mux.scala 46:19:@14199.4]
  wire [7:0] _T_16188; // @[Mux.scala 46:16:@14200.4]
  wire  _T_16189; // @[Mux.scala 46:19:@14201.4]
  wire [7:0] _T_16190; // @[Mux.scala 46:16:@14202.4]
  wire  _T_16248; // @[Mux.scala 46:19:@14204.4]
  wire [7:0] _T_16249; // @[Mux.scala 46:16:@14205.4]
  wire  _T_16250; // @[Mux.scala 46:19:@14206.4]
  wire [7:0] _T_16251; // @[Mux.scala 46:16:@14207.4]
  wire  _T_16252; // @[Mux.scala 46:19:@14208.4]
  wire [7:0] _T_16253; // @[Mux.scala 46:16:@14209.4]
  wire  _T_16254; // @[Mux.scala 46:19:@14210.4]
  wire [7:0] _T_16255; // @[Mux.scala 46:16:@14211.4]
  wire  _T_16256; // @[Mux.scala 46:19:@14212.4]
  wire [7:0] _T_16257; // @[Mux.scala 46:16:@14213.4]
  wire  _T_16258; // @[Mux.scala 46:19:@14214.4]
  wire [7:0] _T_16259; // @[Mux.scala 46:16:@14215.4]
  wire  _T_16260; // @[Mux.scala 46:19:@14216.4]
  wire [7:0] _T_16261; // @[Mux.scala 46:16:@14217.4]
  wire  _T_16262; // @[Mux.scala 46:19:@14218.4]
  wire [7:0] _T_16263; // @[Mux.scala 46:16:@14219.4]
  wire  _T_16264; // @[Mux.scala 46:19:@14220.4]
  wire [7:0] _T_16265; // @[Mux.scala 46:16:@14221.4]
  wire  _T_16266; // @[Mux.scala 46:19:@14222.4]
  wire [7:0] _T_16267; // @[Mux.scala 46:16:@14223.4]
  wire  _T_16268; // @[Mux.scala 46:19:@14224.4]
  wire [7:0] _T_16269; // @[Mux.scala 46:16:@14225.4]
  wire  _T_16270; // @[Mux.scala 46:19:@14226.4]
  wire [7:0] _T_16271; // @[Mux.scala 46:16:@14227.4]
  wire  _T_16272; // @[Mux.scala 46:19:@14228.4]
  wire [7:0] _T_16273; // @[Mux.scala 46:16:@14229.4]
  wire  _T_16274; // @[Mux.scala 46:19:@14230.4]
  wire [7:0] _T_16275; // @[Mux.scala 46:16:@14231.4]
  wire  _T_16276; // @[Mux.scala 46:19:@14232.4]
  wire [7:0] _T_16277; // @[Mux.scala 46:16:@14233.4]
  wire  _T_16278; // @[Mux.scala 46:19:@14234.4]
  wire [7:0] _T_16279; // @[Mux.scala 46:16:@14235.4]
  wire  _T_16280; // @[Mux.scala 46:19:@14236.4]
  wire [7:0] _T_16281; // @[Mux.scala 46:16:@14237.4]
  wire  _T_16282; // @[Mux.scala 46:19:@14238.4]
  wire [7:0] _T_16283; // @[Mux.scala 46:16:@14239.4]
  wire  _T_16284; // @[Mux.scala 46:19:@14240.4]
  wire [7:0] _T_16285; // @[Mux.scala 46:16:@14241.4]
  wire  _T_16286; // @[Mux.scala 46:19:@14242.4]
  wire [7:0] _T_16287; // @[Mux.scala 46:16:@14243.4]
  wire  _T_16288; // @[Mux.scala 46:19:@14244.4]
  wire [7:0] _T_16289; // @[Mux.scala 46:16:@14245.4]
  wire  _T_16290; // @[Mux.scala 46:19:@14246.4]
  wire [7:0] _T_16291; // @[Mux.scala 46:16:@14247.4]
  wire  _T_16292; // @[Mux.scala 46:19:@14248.4]
  wire [7:0] _T_16293; // @[Mux.scala 46:16:@14249.4]
  wire  _T_16294; // @[Mux.scala 46:19:@14250.4]
  wire [7:0] _T_16295; // @[Mux.scala 46:16:@14251.4]
  wire  _T_16296; // @[Mux.scala 46:19:@14252.4]
  wire [7:0] _T_16297; // @[Mux.scala 46:16:@14253.4]
  wire  _T_16298; // @[Mux.scala 46:19:@14254.4]
  wire [7:0] _T_16299; // @[Mux.scala 46:16:@14255.4]
  wire  _T_16300; // @[Mux.scala 46:19:@14256.4]
  wire [7:0] _T_16301; // @[Mux.scala 46:16:@14257.4]
  wire  _T_16302; // @[Mux.scala 46:19:@14258.4]
  wire [7:0] _T_16303; // @[Mux.scala 46:16:@14259.4]
  wire  _T_16304; // @[Mux.scala 46:19:@14260.4]
  wire [7:0] _T_16305; // @[Mux.scala 46:16:@14261.4]
  wire  _T_16306; // @[Mux.scala 46:19:@14262.4]
  wire [7:0] _T_16307; // @[Mux.scala 46:16:@14263.4]
  wire  _T_16308; // @[Mux.scala 46:19:@14264.4]
  wire [7:0] _T_16309; // @[Mux.scala 46:16:@14265.4]
  wire  _T_16310; // @[Mux.scala 46:19:@14266.4]
  wire [7:0] _T_16311; // @[Mux.scala 46:16:@14267.4]
  wire  _T_16312; // @[Mux.scala 46:19:@14268.4]
  wire [7:0] _T_16313; // @[Mux.scala 46:16:@14269.4]
  wire  _T_16314; // @[Mux.scala 46:19:@14270.4]
  wire [7:0] _T_16315; // @[Mux.scala 46:16:@14271.4]
  wire  _T_16316; // @[Mux.scala 46:19:@14272.4]
  wire [7:0] _T_16317; // @[Mux.scala 46:16:@14273.4]
  wire  _T_16318; // @[Mux.scala 46:19:@14274.4]
  wire [7:0] _T_16319; // @[Mux.scala 46:16:@14275.4]
  wire  _T_16320; // @[Mux.scala 46:19:@14276.4]
  wire [7:0] _T_16321; // @[Mux.scala 46:16:@14277.4]
  wire  _T_16322; // @[Mux.scala 46:19:@14278.4]
  wire [7:0] _T_16323; // @[Mux.scala 46:16:@14279.4]
  wire  _T_16324; // @[Mux.scala 46:19:@14280.4]
  wire [7:0] _T_16325; // @[Mux.scala 46:16:@14281.4]
  wire  _T_16326; // @[Mux.scala 46:19:@14282.4]
  wire [7:0] _T_16327; // @[Mux.scala 46:16:@14283.4]
  wire  _T_16328; // @[Mux.scala 46:19:@14284.4]
  wire [7:0] _T_16329; // @[Mux.scala 46:16:@14285.4]
  wire  _T_16330; // @[Mux.scala 46:19:@14286.4]
  wire [7:0] _T_16331; // @[Mux.scala 46:16:@14287.4]
  wire  _T_16332; // @[Mux.scala 46:19:@14288.4]
  wire [7:0] _T_16333; // @[Mux.scala 46:16:@14289.4]
  wire  _T_16334; // @[Mux.scala 46:19:@14290.4]
  wire [7:0] _T_16335; // @[Mux.scala 46:16:@14291.4]
  wire  _T_16336; // @[Mux.scala 46:19:@14292.4]
  wire [7:0] _T_16337; // @[Mux.scala 46:16:@14293.4]
  wire  _T_16338; // @[Mux.scala 46:19:@14294.4]
  wire [7:0] _T_16339; // @[Mux.scala 46:16:@14295.4]
  wire  _T_16340; // @[Mux.scala 46:19:@14296.4]
  wire [7:0] _T_16341; // @[Mux.scala 46:16:@14297.4]
  wire  _T_16342; // @[Mux.scala 46:19:@14298.4]
  wire [7:0] _T_16343; // @[Mux.scala 46:16:@14299.4]
  wire  _T_16344; // @[Mux.scala 46:19:@14300.4]
  wire [7:0] _T_16345; // @[Mux.scala 46:16:@14301.4]
  wire  _T_16346; // @[Mux.scala 46:19:@14302.4]
  wire [7:0] _T_16347; // @[Mux.scala 46:16:@14303.4]
  wire  _T_16348; // @[Mux.scala 46:19:@14304.4]
  wire [7:0] _T_16349; // @[Mux.scala 46:16:@14305.4]
  wire  _T_16350; // @[Mux.scala 46:19:@14306.4]
  wire [7:0] _T_16351; // @[Mux.scala 46:16:@14307.4]
  wire  _T_16352; // @[Mux.scala 46:19:@14308.4]
  wire [7:0] _T_16353; // @[Mux.scala 46:16:@14309.4]
  wire  _T_16354; // @[Mux.scala 46:19:@14310.4]
  wire [7:0] _T_16355; // @[Mux.scala 46:16:@14311.4]
  wire  _T_16356; // @[Mux.scala 46:19:@14312.4]
  wire [7:0] _T_16357; // @[Mux.scala 46:16:@14313.4]
  wire  _T_16358; // @[Mux.scala 46:19:@14314.4]
  wire [7:0] _T_16359; // @[Mux.scala 46:16:@14315.4]
  wire  _T_16418; // @[Mux.scala 46:19:@14317.4]
  wire [7:0] _T_16419; // @[Mux.scala 46:16:@14318.4]
  wire  _T_16420; // @[Mux.scala 46:19:@14319.4]
  wire [7:0] _T_16421; // @[Mux.scala 46:16:@14320.4]
  wire  _T_16422; // @[Mux.scala 46:19:@14321.4]
  wire [7:0] _T_16423; // @[Mux.scala 46:16:@14322.4]
  wire  _T_16424; // @[Mux.scala 46:19:@14323.4]
  wire [7:0] _T_16425; // @[Mux.scala 46:16:@14324.4]
  wire  _T_16426; // @[Mux.scala 46:19:@14325.4]
  wire [7:0] _T_16427; // @[Mux.scala 46:16:@14326.4]
  wire  _T_16428; // @[Mux.scala 46:19:@14327.4]
  wire [7:0] _T_16429; // @[Mux.scala 46:16:@14328.4]
  wire  _T_16430; // @[Mux.scala 46:19:@14329.4]
  wire [7:0] _T_16431; // @[Mux.scala 46:16:@14330.4]
  wire  _T_16432; // @[Mux.scala 46:19:@14331.4]
  wire [7:0] _T_16433; // @[Mux.scala 46:16:@14332.4]
  wire  _T_16434; // @[Mux.scala 46:19:@14333.4]
  wire [7:0] _T_16435; // @[Mux.scala 46:16:@14334.4]
  wire  _T_16436; // @[Mux.scala 46:19:@14335.4]
  wire [7:0] _T_16437; // @[Mux.scala 46:16:@14336.4]
  wire  _T_16438; // @[Mux.scala 46:19:@14337.4]
  wire [7:0] _T_16439; // @[Mux.scala 46:16:@14338.4]
  wire  _T_16440; // @[Mux.scala 46:19:@14339.4]
  wire [7:0] _T_16441; // @[Mux.scala 46:16:@14340.4]
  wire  _T_16442; // @[Mux.scala 46:19:@14341.4]
  wire [7:0] _T_16443; // @[Mux.scala 46:16:@14342.4]
  wire  _T_16444; // @[Mux.scala 46:19:@14343.4]
  wire [7:0] _T_16445; // @[Mux.scala 46:16:@14344.4]
  wire  _T_16446; // @[Mux.scala 46:19:@14345.4]
  wire [7:0] _T_16447; // @[Mux.scala 46:16:@14346.4]
  wire  _T_16448; // @[Mux.scala 46:19:@14347.4]
  wire [7:0] _T_16449; // @[Mux.scala 46:16:@14348.4]
  wire  _T_16450; // @[Mux.scala 46:19:@14349.4]
  wire [7:0] _T_16451; // @[Mux.scala 46:16:@14350.4]
  wire  _T_16452; // @[Mux.scala 46:19:@14351.4]
  wire [7:0] _T_16453; // @[Mux.scala 46:16:@14352.4]
  wire  _T_16454; // @[Mux.scala 46:19:@14353.4]
  wire [7:0] _T_16455; // @[Mux.scala 46:16:@14354.4]
  wire  _T_16456; // @[Mux.scala 46:19:@14355.4]
  wire [7:0] _T_16457; // @[Mux.scala 46:16:@14356.4]
  wire  _T_16458; // @[Mux.scala 46:19:@14357.4]
  wire [7:0] _T_16459; // @[Mux.scala 46:16:@14358.4]
  wire  _T_16460; // @[Mux.scala 46:19:@14359.4]
  wire [7:0] _T_16461; // @[Mux.scala 46:16:@14360.4]
  wire  _T_16462; // @[Mux.scala 46:19:@14361.4]
  wire [7:0] _T_16463; // @[Mux.scala 46:16:@14362.4]
  wire  _T_16464; // @[Mux.scala 46:19:@14363.4]
  wire [7:0] _T_16465; // @[Mux.scala 46:16:@14364.4]
  wire  _T_16466; // @[Mux.scala 46:19:@14365.4]
  wire [7:0] _T_16467; // @[Mux.scala 46:16:@14366.4]
  wire  _T_16468; // @[Mux.scala 46:19:@14367.4]
  wire [7:0] _T_16469; // @[Mux.scala 46:16:@14368.4]
  wire  _T_16470; // @[Mux.scala 46:19:@14369.4]
  wire [7:0] _T_16471; // @[Mux.scala 46:16:@14370.4]
  wire  _T_16472; // @[Mux.scala 46:19:@14371.4]
  wire [7:0] _T_16473; // @[Mux.scala 46:16:@14372.4]
  wire  _T_16474; // @[Mux.scala 46:19:@14373.4]
  wire [7:0] _T_16475; // @[Mux.scala 46:16:@14374.4]
  wire  _T_16476; // @[Mux.scala 46:19:@14375.4]
  wire [7:0] _T_16477; // @[Mux.scala 46:16:@14376.4]
  wire  _T_16478; // @[Mux.scala 46:19:@14377.4]
  wire [7:0] _T_16479; // @[Mux.scala 46:16:@14378.4]
  wire  _T_16480; // @[Mux.scala 46:19:@14379.4]
  wire [7:0] _T_16481; // @[Mux.scala 46:16:@14380.4]
  wire  _T_16482; // @[Mux.scala 46:19:@14381.4]
  wire [7:0] _T_16483; // @[Mux.scala 46:16:@14382.4]
  wire  _T_16484; // @[Mux.scala 46:19:@14383.4]
  wire [7:0] _T_16485; // @[Mux.scala 46:16:@14384.4]
  wire  _T_16486; // @[Mux.scala 46:19:@14385.4]
  wire [7:0] _T_16487; // @[Mux.scala 46:16:@14386.4]
  wire  _T_16488; // @[Mux.scala 46:19:@14387.4]
  wire [7:0] _T_16489; // @[Mux.scala 46:16:@14388.4]
  wire  _T_16490; // @[Mux.scala 46:19:@14389.4]
  wire [7:0] _T_16491; // @[Mux.scala 46:16:@14390.4]
  wire  _T_16492; // @[Mux.scala 46:19:@14391.4]
  wire [7:0] _T_16493; // @[Mux.scala 46:16:@14392.4]
  wire  _T_16494; // @[Mux.scala 46:19:@14393.4]
  wire [7:0] _T_16495; // @[Mux.scala 46:16:@14394.4]
  wire  _T_16496; // @[Mux.scala 46:19:@14395.4]
  wire [7:0] _T_16497; // @[Mux.scala 46:16:@14396.4]
  wire  _T_16498; // @[Mux.scala 46:19:@14397.4]
  wire [7:0] _T_16499; // @[Mux.scala 46:16:@14398.4]
  wire  _T_16500; // @[Mux.scala 46:19:@14399.4]
  wire [7:0] _T_16501; // @[Mux.scala 46:16:@14400.4]
  wire  _T_16502; // @[Mux.scala 46:19:@14401.4]
  wire [7:0] _T_16503; // @[Mux.scala 46:16:@14402.4]
  wire  _T_16504; // @[Mux.scala 46:19:@14403.4]
  wire [7:0] _T_16505; // @[Mux.scala 46:16:@14404.4]
  wire  _T_16506; // @[Mux.scala 46:19:@14405.4]
  wire [7:0] _T_16507; // @[Mux.scala 46:16:@14406.4]
  wire  _T_16508; // @[Mux.scala 46:19:@14407.4]
  wire [7:0] _T_16509; // @[Mux.scala 46:16:@14408.4]
  wire  _T_16510; // @[Mux.scala 46:19:@14409.4]
  wire [7:0] _T_16511; // @[Mux.scala 46:16:@14410.4]
  wire  _T_16512; // @[Mux.scala 46:19:@14411.4]
  wire [7:0] _T_16513; // @[Mux.scala 46:16:@14412.4]
  wire  _T_16514; // @[Mux.scala 46:19:@14413.4]
  wire [7:0] _T_16515; // @[Mux.scala 46:16:@14414.4]
  wire  _T_16516; // @[Mux.scala 46:19:@14415.4]
  wire [7:0] _T_16517; // @[Mux.scala 46:16:@14416.4]
  wire  _T_16518; // @[Mux.scala 46:19:@14417.4]
  wire [7:0] _T_16519; // @[Mux.scala 46:16:@14418.4]
  wire  _T_16520; // @[Mux.scala 46:19:@14419.4]
  wire [7:0] _T_16521; // @[Mux.scala 46:16:@14420.4]
  wire  _T_16522; // @[Mux.scala 46:19:@14421.4]
  wire [7:0] _T_16523; // @[Mux.scala 46:16:@14422.4]
  wire  _T_16524; // @[Mux.scala 46:19:@14423.4]
  wire [7:0] _T_16525; // @[Mux.scala 46:16:@14424.4]
  wire  _T_16526; // @[Mux.scala 46:19:@14425.4]
  wire [7:0] _T_16527; // @[Mux.scala 46:16:@14426.4]
  wire  _T_16528; // @[Mux.scala 46:19:@14427.4]
  wire [7:0] _T_16529; // @[Mux.scala 46:16:@14428.4]
  wire  _T_16530; // @[Mux.scala 46:19:@14429.4]
  wire [7:0] _T_16531; // @[Mux.scala 46:16:@14430.4]
  wire  _T_16591; // @[Mux.scala 46:19:@14432.4]
  wire [7:0] _T_16592; // @[Mux.scala 46:16:@14433.4]
  wire  _T_16593; // @[Mux.scala 46:19:@14434.4]
  wire [7:0] _T_16594; // @[Mux.scala 46:16:@14435.4]
  wire  _T_16595; // @[Mux.scala 46:19:@14436.4]
  wire [7:0] _T_16596; // @[Mux.scala 46:16:@14437.4]
  wire  _T_16597; // @[Mux.scala 46:19:@14438.4]
  wire [7:0] _T_16598; // @[Mux.scala 46:16:@14439.4]
  wire  _T_16599; // @[Mux.scala 46:19:@14440.4]
  wire [7:0] _T_16600; // @[Mux.scala 46:16:@14441.4]
  wire  _T_16601; // @[Mux.scala 46:19:@14442.4]
  wire [7:0] _T_16602; // @[Mux.scala 46:16:@14443.4]
  wire  _T_16603; // @[Mux.scala 46:19:@14444.4]
  wire [7:0] _T_16604; // @[Mux.scala 46:16:@14445.4]
  wire  _T_16605; // @[Mux.scala 46:19:@14446.4]
  wire [7:0] _T_16606; // @[Mux.scala 46:16:@14447.4]
  wire  _T_16607; // @[Mux.scala 46:19:@14448.4]
  wire [7:0] _T_16608; // @[Mux.scala 46:16:@14449.4]
  wire  _T_16609; // @[Mux.scala 46:19:@14450.4]
  wire [7:0] _T_16610; // @[Mux.scala 46:16:@14451.4]
  wire  _T_16611; // @[Mux.scala 46:19:@14452.4]
  wire [7:0] _T_16612; // @[Mux.scala 46:16:@14453.4]
  wire  _T_16613; // @[Mux.scala 46:19:@14454.4]
  wire [7:0] _T_16614; // @[Mux.scala 46:16:@14455.4]
  wire  _T_16615; // @[Mux.scala 46:19:@14456.4]
  wire [7:0] _T_16616; // @[Mux.scala 46:16:@14457.4]
  wire  _T_16617; // @[Mux.scala 46:19:@14458.4]
  wire [7:0] _T_16618; // @[Mux.scala 46:16:@14459.4]
  wire  _T_16619; // @[Mux.scala 46:19:@14460.4]
  wire [7:0] _T_16620; // @[Mux.scala 46:16:@14461.4]
  wire  _T_16621; // @[Mux.scala 46:19:@14462.4]
  wire [7:0] _T_16622; // @[Mux.scala 46:16:@14463.4]
  wire  _T_16623; // @[Mux.scala 46:19:@14464.4]
  wire [7:0] _T_16624; // @[Mux.scala 46:16:@14465.4]
  wire  _T_16625; // @[Mux.scala 46:19:@14466.4]
  wire [7:0] _T_16626; // @[Mux.scala 46:16:@14467.4]
  wire  _T_16627; // @[Mux.scala 46:19:@14468.4]
  wire [7:0] _T_16628; // @[Mux.scala 46:16:@14469.4]
  wire  _T_16629; // @[Mux.scala 46:19:@14470.4]
  wire [7:0] _T_16630; // @[Mux.scala 46:16:@14471.4]
  wire  _T_16631; // @[Mux.scala 46:19:@14472.4]
  wire [7:0] _T_16632; // @[Mux.scala 46:16:@14473.4]
  wire  _T_16633; // @[Mux.scala 46:19:@14474.4]
  wire [7:0] _T_16634; // @[Mux.scala 46:16:@14475.4]
  wire  _T_16635; // @[Mux.scala 46:19:@14476.4]
  wire [7:0] _T_16636; // @[Mux.scala 46:16:@14477.4]
  wire  _T_16637; // @[Mux.scala 46:19:@14478.4]
  wire [7:0] _T_16638; // @[Mux.scala 46:16:@14479.4]
  wire  _T_16639; // @[Mux.scala 46:19:@14480.4]
  wire [7:0] _T_16640; // @[Mux.scala 46:16:@14481.4]
  wire  _T_16641; // @[Mux.scala 46:19:@14482.4]
  wire [7:0] _T_16642; // @[Mux.scala 46:16:@14483.4]
  wire  _T_16643; // @[Mux.scala 46:19:@14484.4]
  wire [7:0] _T_16644; // @[Mux.scala 46:16:@14485.4]
  wire  _T_16645; // @[Mux.scala 46:19:@14486.4]
  wire [7:0] _T_16646; // @[Mux.scala 46:16:@14487.4]
  wire  _T_16647; // @[Mux.scala 46:19:@14488.4]
  wire [7:0] _T_16648; // @[Mux.scala 46:16:@14489.4]
  wire  _T_16649; // @[Mux.scala 46:19:@14490.4]
  wire [7:0] _T_16650; // @[Mux.scala 46:16:@14491.4]
  wire  _T_16651; // @[Mux.scala 46:19:@14492.4]
  wire [7:0] _T_16652; // @[Mux.scala 46:16:@14493.4]
  wire  _T_16653; // @[Mux.scala 46:19:@14494.4]
  wire [7:0] _T_16654; // @[Mux.scala 46:16:@14495.4]
  wire  _T_16655; // @[Mux.scala 46:19:@14496.4]
  wire [7:0] _T_16656; // @[Mux.scala 46:16:@14497.4]
  wire  _T_16657; // @[Mux.scala 46:19:@14498.4]
  wire [7:0] _T_16658; // @[Mux.scala 46:16:@14499.4]
  wire  _T_16659; // @[Mux.scala 46:19:@14500.4]
  wire [7:0] _T_16660; // @[Mux.scala 46:16:@14501.4]
  wire  _T_16661; // @[Mux.scala 46:19:@14502.4]
  wire [7:0] _T_16662; // @[Mux.scala 46:16:@14503.4]
  wire  _T_16663; // @[Mux.scala 46:19:@14504.4]
  wire [7:0] _T_16664; // @[Mux.scala 46:16:@14505.4]
  wire  _T_16665; // @[Mux.scala 46:19:@14506.4]
  wire [7:0] _T_16666; // @[Mux.scala 46:16:@14507.4]
  wire  _T_16667; // @[Mux.scala 46:19:@14508.4]
  wire [7:0] _T_16668; // @[Mux.scala 46:16:@14509.4]
  wire  _T_16669; // @[Mux.scala 46:19:@14510.4]
  wire [7:0] _T_16670; // @[Mux.scala 46:16:@14511.4]
  wire  _T_16671; // @[Mux.scala 46:19:@14512.4]
  wire [7:0] _T_16672; // @[Mux.scala 46:16:@14513.4]
  wire  _T_16673; // @[Mux.scala 46:19:@14514.4]
  wire [7:0] _T_16674; // @[Mux.scala 46:16:@14515.4]
  wire  _T_16675; // @[Mux.scala 46:19:@14516.4]
  wire [7:0] _T_16676; // @[Mux.scala 46:16:@14517.4]
  wire  _T_16677; // @[Mux.scala 46:19:@14518.4]
  wire [7:0] _T_16678; // @[Mux.scala 46:16:@14519.4]
  wire  _T_16679; // @[Mux.scala 46:19:@14520.4]
  wire [7:0] _T_16680; // @[Mux.scala 46:16:@14521.4]
  wire  _T_16681; // @[Mux.scala 46:19:@14522.4]
  wire [7:0] _T_16682; // @[Mux.scala 46:16:@14523.4]
  wire  _T_16683; // @[Mux.scala 46:19:@14524.4]
  wire [7:0] _T_16684; // @[Mux.scala 46:16:@14525.4]
  wire  _T_16685; // @[Mux.scala 46:19:@14526.4]
  wire [7:0] _T_16686; // @[Mux.scala 46:16:@14527.4]
  wire  _T_16687; // @[Mux.scala 46:19:@14528.4]
  wire [7:0] _T_16688; // @[Mux.scala 46:16:@14529.4]
  wire  _T_16689; // @[Mux.scala 46:19:@14530.4]
  wire [7:0] _T_16690; // @[Mux.scala 46:16:@14531.4]
  wire  _T_16691; // @[Mux.scala 46:19:@14532.4]
  wire [7:0] _T_16692; // @[Mux.scala 46:16:@14533.4]
  wire  _T_16693; // @[Mux.scala 46:19:@14534.4]
  wire [7:0] _T_16694; // @[Mux.scala 46:16:@14535.4]
  wire  _T_16695; // @[Mux.scala 46:19:@14536.4]
  wire [7:0] _T_16696; // @[Mux.scala 46:16:@14537.4]
  wire  _T_16697; // @[Mux.scala 46:19:@14538.4]
  wire [7:0] _T_16698; // @[Mux.scala 46:16:@14539.4]
  wire  _T_16699; // @[Mux.scala 46:19:@14540.4]
  wire [7:0] _T_16700; // @[Mux.scala 46:16:@14541.4]
  wire  _T_16701; // @[Mux.scala 46:19:@14542.4]
  wire [7:0] _T_16702; // @[Mux.scala 46:16:@14543.4]
  wire  _T_16703; // @[Mux.scala 46:19:@14544.4]
  wire [7:0] _T_16704; // @[Mux.scala 46:16:@14545.4]
  wire  _T_16705; // @[Mux.scala 46:19:@14546.4]
  wire [7:0] _T_16706; // @[Mux.scala 46:16:@14547.4]
  wire  _T_16767; // @[Mux.scala 46:19:@14549.4]
  wire [7:0] _T_16768; // @[Mux.scala 46:16:@14550.4]
  wire  _T_16769; // @[Mux.scala 46:19:@14551.4]
  wire [7:0] _T_16770; // @[Mux.scala 46:16:@14552.4]
  wire  _T_16771; // @[Mux.scala 46:19:@14553.4]
  wire [7:0] _T_16772; // @[Mux.scala 46:16:@14554.4]
  wire  _T_16773; // @[Mux.scala 46:19:@14555.4]
  wire [7:0] _T_16774; // @[Mux.scala 46:16:@14556.4]
  wire  _T_16775; // @[Mux.scala 46:19:@14557.4]
  wire [7:0] _T_16776; // @[Mux.scala 46:16:@14558.4]
  wire  _T_16777; // @[Mux.scala 46:19:@14559.4]
  wire [7:0] _T_16778; // @[Mux.scala 46:16:@14560.4]
  wire  _T_16779; // @[Mux.scala 46:19:@14561.4]
  wire [7:0] _T_16780; // @[Mux.scala 46:16:@14562.4]
  wire  _T_16781; // @[Mux.scala 46:19:@14563.4]
  wire [7:0] _T_16782; // @[Mux.scala 46:16:@14564.4]
  wire  _T_16783; // @[Mux.scala 46:19:@14565.4]
  wire [7:0] _T_16784; // @[Mux.scala 46:16:@14566.4]
  wire  _T_16785; // @[Mux.scala 46:19:@14567.4]
  wire [7:0] _T_16786; // @[Mux.scala 46:16:@14568.4]
  wire  _T_16787; // @[Mux.scala 46:19:@14569.4]
  wire [7:0] _T_16788; // @[Mux.scala 46:16:@14570.4]
  wire  _T_16789; // @[Mux.scala 46:19:@14571.4]
  wire [7:0] _T_16790; // @[Mux.scala 46:16:@14572.4]
  wire  _T_16791; // @[Mux.scala 46:19:@14573.4]
  wire [7:0] _T_16792; // @[Mux.scala 46:16:@14574.4]
  wire  _T_16793; // @[Mux.scala 46:19:@14575.4]
  wire [7:0] _T_16794; // @[Mux.scala 46:16:@14576.4]
  wire  _T_16795; // @[Mux.scala 46:19:@14577.4]
  wire [7:0] _T_16796; // @[Mux.scala 46:16:@14578.4]
  wire  _T_16797; // @[Mux.scala 46:19:@14579.4]
  wire [7:0] _T_16798; // @[Mux.scala 46:16:@14580.4]
  wire  _T_16799; // @[Mux.scala 46:19:@14581.4]
  wire [7:0] _T_16800; // @[Mux.scala 46:16:@14582.4]
  wire  _T_16801; // @[Mux.scala 46:19:@14583.4]
  wire [7:0] _T_16802; // @[Mux.scala 46:16:@14584.4]
  wire  _T_16803; // @[Mux.scala 46:19:@14585.4]
  wire [7:0] _T_16804; // @[Mux.scala 46:16:@14586.4]
  wire  _T_16805; // @[Mux.scala 46:19:@14587.4]
  wire [7:0] _T_16806; // @[Mux.scala 46:16:@14588.4]
  wire  _T_16807; // @[Mux.scala 46:19:@14589.4]
  wire [7:0] _T_16808; // @[Mux.scala 46:16:@14590.4]
  wire  _T_16809; // @[Mux.scala 46:19:@14591.4]
  wire [7:0] _T_16810; // @[Mux.scala 46:16:@14592.4]
  wire  _T_16811; // @[Mux.scala 46:19:@14593.4]
  wire [7:0] _T_16812; // @[Mux.scala 46:16:@14594.4]
  wire  _T_16813; // @[Mux.scala 46:19:@14595.4]
  wire [7:0] _T_16814; // @[Mux.scala 46:16:@14596.4]
  wire  _T_16815; // @[Mux.scala 46:19:@14597.4]
  wire [7:0] _T_16816; // @[Mux.scala 46:16:@14598.4]
  wire  _T_16817; // @[Mux.scala 46:19:@14599.4]
  wire [7:0] _T_16818; // @[Mux.scala 46:16:@14600.4]
  wire  _T_16819; // @[Mux.scala 46:19:@14601.4]
  wire [7:0] _T_16820; // @[Mux.scala 46:16:@14602.4]
  wire  _T_16821; // @[Mux.scala 46:19:@14603.4]
  wire [7:0] _T_16822; // @[Mux.scala 46:16:@14604.4]
  wire  _T_16823; // @[Mux.scala 46:19:@14605.4]
  wire [7:0] _T_16824; // @[Mux.scala 46:16:@14606.4]
  wire  _T_16825; // @[Mux.scala 46:19:@14607.4]
  wire [7:0] _T_16826; // @[Mux.scala 46:16:@14608.4]
  wire  _T_16827; // @[Mux.scala 46:19:@14609.4]
  wire [7:0] _T_16828; // @[Mux.scala 46:16:@14610.4]
  wire  _T_16829; // @[Mux.scala 46:19:@14611.4]
  wire [7:0] _T_16830; // @[Mux.scala 46:16:@14612.4]
  wire  _T_16831; // @[Mux.scala 46:19:@14613.4]
  wire [7:0] _T_16832; // @[Mux.scala 46:16:@14614.4]
  wire  _T_16833; // @[Mux.scala 46:19:@14615.4]
  wire [7:0] _T_16834; // @[Mux.scala 46:16:@14616.4]
  wire  _T_16835; // @[Mux.scala 46:19:@14617.4]
  wire [7:0] _T_16836; // @[Mux.scala 46:16:@14618.4]
  wire  _T_16837; // @[Mux.scala 46:19:@14619.4]
  wire [7:0] _T_16838; // @[Mux.scala 46:16:@14620.4]
  wire  _T_16839; // @[Mux.scala 46:19:@14621.4]
  wire [7:0] _T_16840; // @[Mux.scala 46:16:@14622.4]
  wire  _T_16841; // @[Mux.scala 46:19:@14623.4]
  wire [7:0] _T_16842; // @[Mux.scala 46:16:@14624.4]
  wire  _T_16843; // @[Mux.scala 46:19:@14625.4]
  wire [7:0] _T_16844; // @[Mux.scala 46:16:@14626.4]
  wire  _T_16845; // @[Mux.scala 46:19:@14627.4]
  wire [7:0] _T_16846; // @[Mux.scala 46:16:@14628.4]
  wire  _T_16847; // @[Mux.scala 46:19:@14629.4]
  wire [7:0] _T_16848; // @[Mux.scala 46:16:@14630.4]
  wire  _T_16849; // @[Mux.scala 46:19:@14631.4]
  wire [7:0] _T_16850; // @[Mux.scala 46:16:@14632.4]
  wire  _T_16851; // @[Mux.scala 46:19:@14633.4]
  wire [7:0] _T_16852; // @[Mux.scala 46:16:@14634.4]
  wire  _T_16853; // @[Mux.scala 46:19:@14635.4]
  wire [7:0] _T_16854; // @[Mux.scala 46:16:@14636.4]
  wire  _T_16855; // @[Mux.scala 46:19:@14637.4]
  wire [7:0] _T_16856; // @[Mux.scala 46:16:@14638.4]
  wire  _T_16857; // @[Mux.scala 46:19:@14639.4]
  wire [7:0] _T_16858; // @[Mux.scala 46:16:@14640.4]
  wire  _T_16859; // @[Mux.scala 46:19:@14641.4]
  wire [7:0] _T_16860; // @[Mux.scala 46:16:@14642.4]
  wire  _T_16861; // @[Mux.scala 46:19:@14643.4]
  wire [7:0] _T_16862; // @[Mux.scala 46:16:@14644.4]
  wire  _T_16863; // @[Mux.scala 46:19:@14645.4]
  wire [7:0] _T_16864; // @[Mux.scala 46:16:@14646.4]
  wire  _T_16865; // @[Mux.scala 46:19:@14647.4]
  wire [7:0] _T_16866; // @[Mux.scala 46:16:@14648.4]
  wire  _T_16867; // @[Mux.scala 46:19:@14649.4]
  wire [7:0] _T_16868; // @[Mux.scala 46:16:@14650.4]
  wire  _T_16869; // @[Mux.scala 46:19:@14651.4]
  wire [7:0] _T_16870; // @[Mux.scala 46:16:@14652.4]
  wire  _T_16871; // @[Mux.scala 46:19:@14653.4]
  wire [7:0] _T_16872; // @[Mux.scala 46:16:@14654.4]
  wire  _T_16873; // @[Mux.scala 46:19:@14655.4]
  wire [7:0] _T_16874; // @[Mux.scala 46:16:@14656.4]
  wire  _T_16875; // @[Mux.scala 46:19:@14657.4]
  wire [7:0] _T_16876; // @[Mux.scala 46:16:@14658.4]
  wire  _T_16877; // @[Mux.scala 46:19:@14659.4]
  wire [7:0] _T_16878; // @[Mux.scala 46:16:@14660.4]
  wire  _T_16879; // @[Mux.scala 46:19:@14661.4]
  wire [7:0] _T_16880; // @[Mux.scala 46:16:@14662.4]
  wire  _T_16881; // @[Mux.scala 46:19:@14663.4]
  wire [7:0] _T_16882; // @[Mux.scala 46:16:@14664.4]
  wire  _T_16883; // @[Mux.scala 46:19:@14665.4]
  wire [7:0] _T_16884; // @[Mux.scala 46:16:@14666.4]
  wire  _T_16946; // @[Mux.scala 46:19:@14668.4]
  wire [7:0] _T_16947; // @[Mux.scala 46:16:@14669.4]
  wire  _T_16948; // @[Mux.scala 46:19:@14670.4]
  wire [7:0] _T_16949; // @[Mux.scala 46:16:@14671.4]
  wire  _T_16950; // @[Mux.scala 46:19:@14672.4]
  wire [7:0] _T_16951; // @[Mux.scala 46:16:@14673.4]
  wire  _T_16952; // @[Mux.scala 46:19:@14674.4]
  wire [7:0] _T_16953; // @[Mux.scala 46:16:@14675.4]
  wire  _T_16954; // @[Mux.scala 46:19:@14676.4]
  wire [7:0] _T_16955; // @[Mux.scala 46:16:@14677.4]
  wire  _T_16956; // @[Mux.scala 46:19:@14678.4]
  wire [7:0] _T_16957; // @[Mux.scala 46:16:@14679.4]
  wire  _T_16958; // @[Mux.scala 46:19:@14680.4]
  wire [7:0] _T_16959; // @[Mux.scala 46:16:@14681.4]
  wire  _T_16960; // @[Mux.scala 46:19:@14682.4]
  wire [7:0] _T_16961; // @[Mux.scala 46:16:@14683.4]
  wire  _T_16962; // @[Mux.scala 46:19:@14684.4]
  wire [7:0] _T_16963; // @[Mux.scala 46:16:@14685.4]
  wire  _T_16964; // @[Mux.scala 46:19:@14686.4]
  wire [7:0] _T_16965; // @[Mux.scala 46:16:@14687.4]
  wire  _T_16966; // @[Mux.scala 46:19:@14688.4]
  wire [7:0] _T_16967; // @[Mux.scala 46:16:@14689.4]
  wire  _T_16968; // @[Mux.scala 46:19:@14690.4]
  wire [7:0] _T_16969; // @[Mux.scala 46:16:@14691.4]
  wire  _T_16970; // @[Mux.scala 46:19:@14692.4]
  wire [7:0] _T_16971; // @[Mux.scala 46:16:@14693.4]
  wire  _T_16972; // @[Mux.scala 46:19:@14694.4]
  wire [7:0] _T_16973; // @[Mux.scala 46:16:@14695.4]
  wire  _T_16974; // @[Mux.scala 46:19:@14696.4]
  wire [7:0] _T_16975; // @[Mux.scala 46:16:@14697.4]
  wire  _T_16976; // @[Mux.scala 46:19:@14698.4]
  wire [7:0] _T_16977; // @[Mux.scala 46:16:@14699.4]
  wire  _T_16978; // @[Mux.scala 46:19:@14700.4]
  wire [7:0] _T_16979; // @[Mux.scala 46:16:@14701.4]
  wire  _T_16980; // @[Mux.scala 46:19:@14702.4]
  wire [7:0] _T_16981; // @[Mux.scala 46:16:@14703.4]
  wire  _T_16982; // @[Mux.scala 46:19:@14704.4]
  wire [7:0] _T_16983; // @[Mux.scala 46:16:@14705.4]
  wire  _T_16984; // @[Mux.scala 46:19:@14706.4]
  wire [7:0] _T_16985; // @[Mux.scala 46:16:@14707.4]
  wire  _T_16986; // @[Mux.scala 46:19:@14708.4]
  wire [7:0] _T_16987; // @[Mux.scala 46:16:@14709.4]
  wire  _T_16988; // @[Mux.scala 46:19:@14710.4]
  wire [7:0] _T_16989; // @[Mux.scala 46:16:@14711.4]
  wire  _T_16990; // @[Mux.scala 46:19:@14712.4]
  wire [7:0] _T_16991; // @[Mux.scala 46:16:@14713.4]
  wire  _T_16992; // @[Mux.scala 46:19:@14714.4]
  wire [7:0] _T_16993; // @[Mux.scala 46:16:@14715.4]
  wire  _T_16994; // @[Mux.scala 46:19:@14716.4]
  wire [7:0] _T_16995; // @[Mux.scala 46:16:@14717.4]
  wire  _T_16996; // @[Mux.scala 46:19:@14718.4]
  wire [7:0] _T_16997; // @[Mux.scala 46:16:@14719.4]
  wire  _T_16998; // @[Mux.scala 46:19:@14720.4]
  wire [7:0] _T_16999; // @[Mux.scala 46:16:@14721.4]
  wire  _T_17000; // @[Mux.scala 46:19:@14722.4]
  wire [7:0] _T_17001; // @[Mux.scala 46:16:@14723.4]
  wire  _T_17002; // @[Mux.scala 46:19:@14724.4]
  wire [7:0] _T_17003; // @[Mux.scala 46:16:@14725.4]
  wire  _T_17004; // @[Mux.scala 46:19:@14726.4]
  wire [7:0] _T_17005; // @[Mux.scala 46:16:@14727.4]
  wire  _T_17006; // @[Mux.scala 46:19:@14728.4]
  wire [7:0] _T_17007; // @[Mux.scala 46:16:@14729.4]
  wire  _T_17008; // @[Mux.scala 46:19:@14730.4]
  wire [7:0] _T_17009; // @[Mux.scala 46:16:@14731.4]
  wire  _T_17010; // @[Mux.scala 46:19:@14732.4]
  wire [7:0] _T_17011; // @[Mux.scala 46:16:@14733.4]
  wire  _T_17012; // @[Mux.scala 46:19:@14734.4]
  wire [7:0] _T_17013; // @[Mux.scala 46:16:@14735.4]
  wire  _T_17014; // @[Mux.scala 46:19:@14736.4]
  wire [7:0] _T_17015; // @[Mux.scala 46:16:@14737.4]
  wire  _T_17016; // @[Mux.scala 46:19:@14738.4]
  wire [7:0] _T_17017; // @[Mux.scala 46:16:@14739.4]
  wire  _T_17018; // @[Mux.scala 46:19:@14740.4]
  wire [7:0] _T_17019; // @[Mux.scala 46:16:@14741.4]
  wire  _T_17020; // @[Mux.scala 46:19:@14742.4]
  wire [7:0] _T_17021; // @[Mux.scala 46:16:@14743.4]
  wire  _T_17022; // @[Mux.scala 46:19:@14744.4]
  wire [7:0] _T_17023; // @[Mux.scala 46:16:@14745.4]
  wire  _T_17024; // @[Mux.scala 46:19:@14746.4]
  wire [7:0] _T_17025; // @[Mux.scala 46:16:@14747.4]
  wire  _T_17026; // @[Mux.scala 46:19:@14748.4]
  wire [7:0] _T_17027; // @[Mux.scala 46:16:@14749.4]
  wire  _T_17028; // @[Mux.scala 46:19:@14750.4]
  wire [7:0] _T_17029; // @[Mux.scala 46:16:@14751.4]
  wire  _T_17030; // @[Mux.scala 46:19:@14752.4]
  wire [7:0] _T_17031; // @[Mux.scala 46:16:@14753.4]
  wire  _T_17032; // @[Mux.scala 46:19:@14754.4]
  wire [7:0] _T_17033; // @[Mux.scala 46:16:@14755.4]
  wire  _T_17034; // @[Mux.scala 46:19:@14756.4]
  wire [7:0] _T_17035; // @[Mux.scala 46:16:@14757.4]
  wire  _T_17036; // @[Mux.scala 46:19:@14758.4]
  wire [7:0] _T_17037; // @[Mux.scala 46:16:@14759.4]
  wire  _T_17038; // @[Mux.scala 46:19:@14760.4]
  wire [7:0] _T_17039; // @[Mux.scala 46:16:@14761.4]
  wire  _T_17040; // @[Mux.scala 46:19:@14762.4]
  wire [7:0] _T_17041; // @[Mux.scala 46:16:@14763.4]
  wire  _T_17042; // @[Mux.scala 46:19:@14764.4]
  wire [7:0] _T_17043; // @[Mux.scala 46:16:@14765.4]
  wire  _T_17044; // @[Mux.scala 46:19:@14766.4]
  wire [7:0] _T_17045; // @[Mux.scala 46:16:@14767.4]
  wire  _T_17046; // @[Mux.scala 46:19:@14768.4]
  wire [7:0] _T_17047; // @[Mux.scala 46:16:@14769.4]
  wire  _T_17048; // @[Mux.scala 46:19:@14770.4]
  wire [7:0] _T_17049; // @[Mux.scala 46:16:@14771.4]
  wire  _T_17050; // @[Mux.scala 46:19:@14772.4]
  wire [7:0] _T_17051; // @[Mux.scala 46:16:@14773.4]
  wire  _T_17052; // @[Mux.scala 46:19:@14774.4]
  wire [7:0] _T_17053; // @[Mux.scala 46:16:@14775.4]
  wire  _T_17054; // @[Mux.scala 46:19:@14776.4]
  wire [7:0] _T_17055; // @[Mux.scala 46:16:@14777.4]
  wire  _T_17056; // @[Mux.scala 46:19:@14778.4]
  wire [7:0] _T_17057; // @[Mux.scala 46:16:@14779.4]
  wire  _T_17058; // @[Mux.scala 46:19:@14780.4]
  wire [7:0] _T_17059; // @[Mux.scala 46:16:@14781.4]
  wire  _T_17060; // @[Mux.scala 46:19:@14782.4]
  wire [7:0] _T_17061; // @[Mux.scala 46:16:@14783.4]
  wire  _T_17062; // @[Mux.scala 46:19:@14784.4]
  wire [7:0] _T_17063; // @[Mux.scala 46:16:@14785.4]
  wire  _T_17064; // @[Mux.scala 46:19:@14786.4]
  wire [7:0] _T_17065; // @[Mux.scala 46:16:@14787.4]
  wire  _T_17128; // @[Mux.scala 46:19:@14789.4]
  wire [7:0] _T_17129; // @[Mux.scala 46:16:@14790.4]
  wire  _T_17130; // @[Mux.scala 46:19:@14791.4]
  wire [7:0] _T_17131; // @[Mux.scala 46:16:@14792.4]
  wire  _T_17132; // @[Mux.scala 46:19:@14793.4]
  wire [7:0] _T_17133; // @[Mux.scala 46:16:@14794.4]
  wire  _T_17134; // @[Mux.scala 46:19:@14795.4]
  wire [7:0] _T_17135; // @[Mux.scala 46:16:@14796.4]
  wire  _T_17136; // @[Mux.scala 46:19:@14797.4]
  wire [7:0] _T_17137; // @[Mux.scala 46:16:@14798.4]
  wire  _T_17138; // @[Mux.scala 46:19:@14799.4]
  wire [7:0] _T_17139; // @[Mux.scala 46:16:@14800.4]
  wire  _T_17140; // @[Mux.scala 46:19:@14801.4]
  wire [7:0] _T_17141; // @[Mux.scala 46:16:@14802.4]
  wire  _T_17142; // @[Mux.scala 46:19:@14803.4]
  wire [7:0] _T_17143; // @[Mux.scala 46:16:@14804.4]
  wire  _T_17144; // @[Mux.scala 46:19:@14805.4]
  wire [7:0] _T_17145; // @[Mux.scala 46:16:@14806.4]
  wire  _T_17146; // @[Mux.scala 46:19:@14807.4]
  wire [7:0] _T_17147; // @[Mux.scala 46:16:@14808.4]
  wire  _T_17148; // @[Mux.scala 46:19:@14809.4]
  wire [7:0] _T_17149; // @[Mux.scala 46:16:@14810.4]
  wire  _T_17150; // @[Mux.scala 46:19:@14811.4]
  wire [7:0] _T_17151; // @[Mux.scala 46:16:@14812.4]
  wire  _T_17152; // @[Mux.scala 46:19:@14813.4]
  wire [7:0] _T_17153; // @[Mux.scala 46:16:@14814.4]
  wire  _T_17154; // @[Mux.scala 46:19:@14815.4]
  wire [7:0] _T_17155; // @[Mux.scala 46:16:@14816.4]
  wire  _T_17156; // @[Mux.scala 46:19:@14817.4]
  wire [7:0] _T_17157; // @[Mux.scala 46:16:@14818.4]
  wire  _T_17158; // @[Mux.scala 46:19:@14819.4]
  wire [7:0] _T_17159; // @[Mux.scala 46:16:@14820.4]
  wire  _T_17160; // @[Mux.scala 46:19:@14821.4]
  wire [7:0] _T_17161; // @[Mux.scala 46:16:@14822.4]
  wire  _T_17162; // @[Mux.scala 46:19:@14823.4]
  wire [7:0] _T_17163; // @[Mux.scala 46:16:@14824.4]
  wire  _T_17164; // @[Mux.scala 46:19:@14825.4]
  wire [7:0] _T_17165; // @[Mux.scala 46:16:@14826.4]
  wire  _T_17166; // @[Mux.scala 46:19:@14827.4]
  wire [7:0] _T_17167; // @[Mux.scala 46:16:@14828.4]
  wire  _T_17168; // @[Mux.scala 46:19:@14829.4]
  wire [7:0] _T_17169; // @[Mux.scala 46:16:@14830.4]
  wire  _T_17170; // @[Mux.scala 46:19:@14831.4]
  wire [7:0] _T_17171; // @[Mux.scala 46:16:@14832.4]
  wire  _T_17172; // @[Mux.scala 46:19:@14833.4]
  wire [7:0] _T_17173; // @[Mux.scala 46:16:@14834.4]
  wire  _T_17174; // @[Mux.scala 46:19:@14835.4]
  wire [7:0] _T_17175; // @[Mux.scala 46:16:@14836.4]
  wire  _T_17176; // @[Mux.scala 46:19:@14837.4]
  wire [7:0] _T_17177; // @[Mux.scala 46:16:@14838.4]
  wire  _T_17178; // @[Mux.scala 46:19:@14839.4]
  wire [7:0] _T_17179; // @[Mux.scala 46:16:@14840.4]
  wire  _T_17180; // @[Mux.scala 46:19:@14841.4]
  wire [7:0] _T_17181; // @[Mux.scala 46:16:@14842.4]
  wire  _T_17182; // @[Mux.scala 46:19:@14843.4]
  wire [7:0] _T_17183; // @[Mux.scala 46:16:@14844.4]
  wire  _T_17184; // @[Mux.scala 46:19:@14845.4]
  wire [7:0] _T_17185; // @[Mux.scala 46:16:@14846.4]
  wire  _T_17186; // @[Mux.scala 46:19:@14847.4]
  wire [7:0] _T_17187; // @[Mux.scala 46:16:@14848.4]
  wire  _T_17188; // @[Mux.scala 46:19:@14849.4]
  wire [7:0] _T_17189; // @[Mux.scala 46:16:@14850.4]
  wire  _T_17190; // @[Mux.scala 46:19:@14851.4]
  wire [7:0] _T_17191; // @[Mux.scala 46:16:@14852.4]
  wire  _T_17192; // @[Mux.scala 46:19:@14853.4]
  wire [7:0] _T_17193; // @[Mux.scala 46:16:@14854.4]
  wire  _T_17194; // @[Mux.scala 46:19:@14855.4]
  wire [7:0] _T_17195; // @[Mux.scala 46:16:@14856.4]
  wire  _T_17196; // @[Mux.scala 46:19:@14857.4]
  wire [7:0] _T_17197; // @[Mux.scala 46:16:@14858.4]
  wire  _T_17198; // @[Mux.scala 46:19:@14859.4]
  wire [7:0] _T_17199; // @[Mux.scala 46:16:@14860.4]
  wire  _T_17200; // @[Mux.scala 46:19:@14861.4]
  wire [7:0] _T_17201; // @[Mux.scala 46:16:@14862.4]
  wire  _T_17202; // @[Mux.scala 46:19:@14863.4]
  wire [7:0] _T_17203; // @[Mux.scala 46:16:@14864.4]
  wire  _T_17204; // @[Mux.scala 46:19:@14865.4]
  wire [7:0] _T_17205; // @[Mux.scala 46:16:@14866.4]
  wire  _T_17206; // @[Mux.scala 46:19:@14867.4]
  wire [7:0] _T_17207; // @[Mux.scala 46:16:@14868.4]
  wire  _T_17208; // @[Mux.scala 46:19:@14869.4]
  wire [7:0] _T_17209; // @[Mux.scala 46:16:@14870.4]
  wire  _T_17210; // @[Mux.scala 46:19:@14871.4]
  wire [7:0] _T_17211; // @[Mux.scala 46:16:@14872.4]
  wire  _T_17212; // @[Mux.scala 46:19:@14873.4]
  wire [7:0] _T_17213; // @[Mux.scala 46:16:@14874.4]
  wire  _T_17214; // @[Mux.scala 46:19:@14875.4]
  wire [7:0] _T_17215; // @[Mux.scala 46:16:@14876.4]
  wire  _T_17216; // @[Mux.scala 46:19:@14877.4]
  wire [7:0] _T_17217; // @[Mux.scala 46:16:@14878.4]
  wire  _T_17218; // @[Mux.scala 46:19:@14879.4]
  wire [7:0] _T_17219; // @[Mux.scala 46:16:@14880.4]
  wire  _T_17220; // @[Mux.scala 46:19:@14881.4]
  wire [7:0] _T_17221; // @[Mux.scala 46:16:@14882.4]
  wire  _T_17222; // @[Mux.scala 46:19:@14883.4]
  wire [7:0] _T_17223; // @[Mux.scala 46:16:@14884.4]
  wire  _T_17224; // @[Mux.scala 46:19:@14885.4]
  wire [7:0] _T_17225; // @[Mux.scala 46:16:@14886.4]
  wire  _T_17226; // @[Mux.scala 46:19:@14887.4]
  wire [7:0] _T_17227; // @[Mux.scala 46:16:@14888.4]
  wire  _T_17228; // @[Mux.scala 46:19:@14889.4]
  wire [7:0] _T_17229; // @[Mux.scala 46:16:@14890.4]
  wire  _T_17230; // @[Mux.scala 46:19:@14891.4]
  wire [7:0] _T_17231; // @[Mux.scala 46:16:@14892.4]
  wire  _T_17232; // @[Mux.scala 46:19:@14893.4]
  wire [7:0] _T_17233; // @[Mux.scala 46:16:@14894.4]
  wire  _T_17234; // @[Mux.scala 46:19:@14895.4]
  wire [7:0] _T_17235; // @[Mux.scala 46:16:@14896.4]
  wire  _T_17236; // @[Mux.scala 46:19:@14897.4]
  wire [7:0] _T_17237; // @[Mux.scala 46:16:@14898.4]
  wire  _T_17238; // @[Mux.scala 46:19:@14899.4]
  wire [7:0] _T_17239; // @[Mux.scala 46:16:@14900.4]
  wire  _T_17240; // @[Mux.scala 46:19:@14901.4]
  wire [7:0] _T_17241; // @[Mux.scala 46:16:@14902.4]
  wire  _T_17242; // @[Mux.scala 46:19:@14903.4]
  wire [7:0] _T_17243; // @[Mux.scala 46:16:@14904.4]
  wire  _T_17244; // @[Mux.scala 46:19:@14905.4]
  wire [7:0] _T_17245; // @[Mux.scala 46:16:@14906.4]
  wire  _T_17246; // @[Mux.scala 46:19:@14907.4]
  wire [7:0] _T_17247; // @[Mux.scala 46:16:@14908.4]
  wire  _T_17248; // @[Mux.scala 46:19:@14909.4]
  wire [7:0] _T_17249; // @[Mux.scala 46:16:@14910.4]
  wire  _T_17313; // @[Mux.scala 46:19:@14912.4]
  wire [7:0] _T_17314; // @[Mux.scala 46:16:@14913.4]
  wire  _T_17315; // @[Mux.scala 46:19:@14914.4]
  wire [7:0] _T_17316; // @[Mux.scala 46:16:@14915.4]
  wire  _T_17317; // @[Mux.scala 46:19:@14916.4]
  wire [7:0] _T_17318; // @[Mux.scala 46:16:@14917.4]
  wire  _T_17319; // @[Mux.scala 46:19:@14918.4]
  wire [7:0] _T_17320; // @[Mux.scala 46:16:@14919.4]
  wire  _T_17321; // @[Mux.scala 46:19:@14920.4]
  wire [7:0] _T_17322; // @[Mux.scala 46:16:@14921.4]
  wire  _T_17323; // @[Mux.scala 46:19:@14922.4]
  wire [7:0] _T_17324; // @[Mux.scala 46:16:@14923.4]
  wire  _T_17325; // @[Mux.scala 46:19:@14924.4]
  wire [7:0] _T_17326; // @[Mux.scala 46:16:@14925.4]
  wire  _T_17327; // @[Mux.scala 46:19:@14926.4]
  wire [7:0] _T_17328; // @[Mux.scala 46:16:@14927.4]
  wire  _T_17329; // @[Mux.scala 46:19:@14928.4]
  wire [7:0] _T_17330; // @[Mux.scala 46:16:@14929.4]
  wire  _T_17331; // @[Mux.scala 46:19:@14930.4]
  wire [7:0] _T_17332; // @[Mux.scala 46:16:@14931.4]
  wire  _T_17333; // @[Mux.scala 46:19:@14932.4]
  wire [7:0] _T_17334; // @[Mux.scala 46:16:@14933.4]
  wire  _T_17335; // @[Mux.scala 46:19:@14934.4]
  wire [7:0] _T_17336; // @[Mux.scala 46:16:@14935.4]
  wire  _T_17337; // @[Mux.scala 46:19:@14936.4]
  wire [7:0] _T_17338; // @[Mux.scala 46:16:@14937.4]
  wire  _T_17339; // @[Mux.scala 46:19:@14938.4]
  wire [7:0] _T_17340; // @[Mux.scala 46:16:@14939.4]
  wire  _T_17341; // @[Mux.scala 46:19:@14940.4]
  wire [7:0] _T_17342; // @[Mux.scala 46:16:@14941.4]
  wire  _T_17343; // @[Mux.scala 46:19:@14942.4]
  wire [7:0] _T_17344; // @[Mux.scala 46:16:@14943.4]
  wire  _T_17345; // @[Mux.scala 46:19:@14944.4]
  wire [7:0] _T_17346; // @[Mux.scala 46:16:@14945.4]
  wire  _T_17347; // @[Mux.scala 46:19:@14946.4]
  wire [7:0] _T_17348; // @[Mux.scala 46:16:@14947.4]
  wire  _T_17349; // @[Mux.scala 46:19:@14948.4]
  wire [7:0] _T_17350; // @[Mux.scala 46:16:@14949.4]
  wire  _T_17351; // @[Mux.scala 46:19:@14950.4]
  wire [7:0] _T_17352; // @[Mux.scala 46:16:@14951.4]
  wire  _T_17353; // @[Mux.scala 46:19:@14952.4]
  wire [7:0] _T_17354; // @[Mux.scala 46:16:@14953.4]
  wire  _T_17355; // @[Mux.scala 46:19:@14954.4]
  wire [7:0] _T_17356; // @[Mux.scala 46:16:@14955.4]
  wire  _T_17357; // @[Mux.scala 46:19:@14956.4]
  wire [7:0] _T_17358; // @[Mux.scala 46:16:@14957.4]
  wire  _T_17359; // @[Mux.scala 46:19:@14958.4]
  wire [7:0] _T_17360; // @[Mux.scala 46:16:@14959.4]
  wire  _T_17361; // @[Mux.scala 46:19:@14960.4]
  wire [7:0] _T_17362; // @[Mux.scala 46:16:@14961.4]
  wire  _T_17363; // @[Mux.scala 46:19:@14962.4]
  wire [7:0] _T_17364; // @[Mux.scala 46:16:@14963.4]
  wire  _T_17365; // @[Mux.scala 46:19:@14964.4]
  wire [7:0] _T_17366; // @[Mux.scala 46:16:@14965.4]
  wire  _T_17367; // @[Mux.scala 46:19:@14966.4]
  wire [7:0] _T_17368; // @[Mux.scala 46:16:@14967.4]
  wire  _T_17369; // @[Mux.scala 46:19:@14968.4]
  wire [7:0] _T_17370; // @[Mux.scala 46:16:@14969.4]
  wire  _T_17371; // @[Mux.scala 46:19:@14970.4]
  wire [7:0] _T_17372; // @[Mux.scala 46:16:@14971.4]
  wire  _T_17373; // @[Mux.scala 46:19:@14972.4]
  wire [7:0] _T_17374; // @[Mux.scala 46:16:@14973.4]
  wire  _T_17375; // @[Mux.scala 46:19:@14974.4]
  wire [7:0] _T_17376; // @[Mux.scala 46:16:@14975.4]
  wire  _T_17377; // @[Mux.scala 46:19:@14976.4]
  wire [7:0] _T_17378; // @[Mux.scala 46:16:@14977.4]
  wire  _T_17379; // @[Mux.scala 46:19:@14978.4]
  wire [7:0] _T_17380; // @[Mux.scala 46:16:@14979.4]
  wire  _T_17381; // @[Mux.scala 46:19:@14980.4]
  wire [7:0] _T_17382; // @[Mux.scala 46:16:@14981.4]
  wire  _T_17383; // @[Mux.scala 46:19:@14982.4]
  wire [7:0] _T_17384; // @[Mux.scala 46:16:@14983.4]
  wire  _T_17385; // @[Mux.scala 46:19:@14984.4]
  wire [7:0] _T_17386; // @[Mux.scala 46:16:@14985.4]
  wire  _T_17387; // @[Mux.scala 46:19:@14986.4]
  wire [7:0] _T_17388; // @[Mux.scala 46:16:@14987.4]
  wire  _T_17389; // @[Mux.scala 46:19:@14988.4]
  wire [7:0] _T_17390; // @[Mux.scala 46:16:@14989.4]
  wire  _T_17391; // @[Mux.scala 46:19:@14990.4]
  wire [7:0] _T_17392; // @[Mux.scala 46:16:@14991.4]
  wire  _T_17393; // @[Mux.scala 46:19:@14992.4]
  wire [7:0] _T_17394; // @[Mux.scala 46:16:@14993.4]
  wire  _T_17395; // @[Mux.scala 46:19:@14994.4]
  wire [7:0] _T_17396; // @[Mux.scala 46:16:@14995.4]
  wire  _T_17397; // @[Mux.scala 46:19:@14996.4]
  wire [7:0] _T_17398; // @[Mux.scala 46:16:@14997.4]
  wire  _T_17399; // @[Mux.scala 46:19:@14998.4]
  wire [7:0] _T_17400; // @[Mux.scala 46:16:@14999.4]
  wire  _T_17401; // @[Mux.scala 46:19:@15000.4]
  wire [7:0] _T_17402; // @[Mux.scala 46:16:@15001.4]
  wire  _T_17403; // @[Mux.scala 46:19:@15002.4]
  wire [7:0] _T_17404; // @[Mux.scala 46:16:@15003.4]
  wire  _T_17405; // @[Mux.scala 46:19:@15004.4]
  wire [7:0] _T_17406; // @[Mux.scala 46:16:@15005.4]
  wire  _T_17407; // @[Mux.scala 46:19:@15006.4]
  wire [7:0] _T_17408; // @[Mux.scala 46:16:@15007.4]
  wire  _T_17409; // @[Mux.scala 46:19:@15008.4]
  wire [7:0] _T_17410; // @[Mux.scala 46:16:@15009.4]
  wire  _T_17411; // @[Mux.scala 46:19:@15010.4]
  wire [7:0] _T_17412; // @[Mux.scala 46:16:@15011.4]
  wire  _T_17413; // @[Mux.scala 46:19:@15012.4]
  wire [7:0] _T_17414; // @[Mux.scala 46:16:@15013.4]
  wire  _T_17415; // @[Mux.scala 46:19:@15014.4]
  wire [7:0] _T_17416; // @[Mux.scala 46:16:@15015.4]
  wire  _T_17417; // @[Mux.scala 46:19:@15016.4]
  wire [7:0] _T_17418; // @[Mux.scala 46:16:@15017.4]
  wire  _T_17419; // @[Mux.scala 46:19:@15018.4]
  wire [7:0] _T_17420; // @[Mux.scala 46:16:@15019.4]
  wire  _T_17421; // @[Mux.scala 46:19:@15020.4]
  wire [7:0] _T_17422; // @[Mux.scala 46:16:@15021.4]
  wire  _T_17423; // @[Mux.scala 46:19:@15022.4]
  wire [7:0] _T_17424; // @[Mux.scala 46:16:@15023.4]
  wire  _T_17425; // @[Mux.scala 46:19:@15024.4]
  wire [7:0] _T_17426; // @[Mux.scala 46:16:@15025.4]
  wire  _T_17427; // @[Mux.scala 46:19:@15026.4]
  wire [7:0] _T_17428; // @[Mux.scala 46:16:@15027.4]
  wire  _T_17429; // @[Mux.scala 46:19:@15028.4]
  wire [7:0] _T_17430; // @[Mux.scala 46:16:@15029.4]
  wire  _T_17431; // @[Mux.scala 46:19:@15030.4]
  wire [7:0] _T_17432; // @[Mux.scala 46:16:@15031.4]
  wire  _T_17433; // @[Mux.scala 46:19:@15032.4]
  wire [7:0] _T_17434; // @[Mux.scala 46:16:@15033.4]
  wire  _T_17435; // @[Mux.scala 46:19:@15034.4]
  wire [7:0] _T_17436; // @[Mux.scala 46:16:@15035.4]
  wire  _T_17501; // @[Mux.scala 46:19:@15037.4]
  wire [7:0] _T_17502; // @[Mux.scala 46:16:@15038.4]
  wire  _T_17503; // @[Mux.scala 46:19:@15039.4]
  wire [7:0] _T_17504; // @[Mux.scala 46:16:@15040.4]
  wire  _T_17505; // @[Mux.scala 46:19:@15041.4]
  wire [7:0] _T_17506; // @[Mux.scala 46:16:@15042.4]
  wire  _T_17507; // @[Mux.scala 46:19:@15043.4]
  wire [7:0] _T_17508; // @[Mux.scala 46:16:@15044.4]
  wire  _T_17509; // @[Mux.scala 46:19:@15045.4]
  wire [7:0] _T_17510; // @[Mux.scala 46:16:@15046.4]
  wire  _T_17511; // @[Mux.scala 46:19:@15047.4]
  wire [7:0] _T_17512; // @[Mux.scala 46:16:@15048.4]
  wire  _T_17513; // @[Mux.scala 46:19:@15049.4]
  wire [7:0] _T_17514; // @[Mux.scala 46:16:@15050.4]
  wire  _T_17515; // @[Mux.scala 46:19:@15051.4]
  wire [7:0] _T_17516; // @[Mux.scala 46:16:@15052.4]
  wire  _T_17517; // @[Mux.scala 46:19:@15053.4]
  wire [7:0] _T_17518; // @[Mux.scala 46:16:@15054.4]
  wire  _T_17519; // @[Mux.scala 46:19:@15055.4]
  wire [7:0] _T_17520; // @[Mux.scala 46:16:@15056.4]
  wire  _T_17521; // @[Mux.scala 46:19:@15057.4]
  wire [7:0] _T_17522; // @[Mux.scala 46:16:@15058.4]
  wire  _T_17523; // @[Mux.scala 46:19:@15059.4]
  wire [7:0] _T_17524; // @[Mux.scala 46:16:@15060.4]
  wire  _T_17525; // @[Mux.scala 46:19:@15061.4]
  wire [7:0] _T_17526; // @[Mux.scala 46:16:@15062.4]
  wire  _T_17527; // @[Mux.scala 46:19:@15063.4]
  wire [7:0] _T_17528; // @[Mux.scala 46:16:@15064.4]
  wire  _T_17529; // @[Mux.scala 46:19:@15065.4]
  wire [7:0] _T_17530; // @[Mux.scala 46:16:@15066.4]
  wire  _T_17531; // @[Mux.scala 46:19:@15067.4]
  wire [7:0] _T_17532; // @[Mux.scala 46:16:@15068.4]
  wire  _T_17533; // @[Mux.scala 46:19:@15069.4]
  wire [7:0] _T_17534; // @[Mux.scala 46:16:@15070.4]
  wire  _T_17535; // @[Mux.scala 46:19:@15071.4]
  wire [7:0] _T_17536; // @[Mux.scala 46:16:@15072.4]
  wire  _T_17537; // @[Mux.scala 46:19:@15073.4]
  wire [7:0] _T_17538; // @[Mux.scala 46:16:@15074.4]
  wire  _T_17539; // @[Mux.scala 46:19:@15075.4]
  wire [7:0] _T_17540; // @[Mux.scala 46:16:@15076.4]
  wire  _T_17541; // @[Mux.scala 46:19:@15077.4]
  wire [7:0] _T_17542; // @[Mux.scala 46:16:@15078.4]
  wire  _T_17543; // @[Mux.scala 46:19:@15079.4]
  wire [7:0] _T_17544; // @[Mux.scala 46:16:@15080.4]
  wire  _T_17545; // @[Mux.scala 46:19:@15081.4]
  wire [7:0] _T_17546; // @[Mux.scala 46:16:@15082.4]
  wire  _T_17547; // @[Mux.scala 46:19:@15083.4]
  wire [7:0] _T_17548; // @[Mux.scala 46:16:@15084.4]
  wire  _T_17549; // @[Mux.scala 46:19:@15085.4]
  wire [7:0] _T_17550; // @[Mux.scala 46:16:@15086.4]
  wire  _T_17551; // @[Mux.scala 46:19:@15087.4]
  wire [7:0] _T_17552; // @[Mux.scala 46:16:@15088.4]
  wire  _T_17553; // @[Mux.scala 46:19:@15089.4]
  wire [7:0] _T_17554; // @[Mux.scala 46:16:@15090.4]
  wire  _T_17555; // @[Mux.scala 46:19:@15091.4]
  wire [7:0] _T_17556; // @[Mux.scala 46:16:@15092.4]
  wire  _T_17557; // @[Mux.scala 46:19:@15093.4]
  wire [7:0] _T_17558; // @[Mux.scala 46:16:@15094.4]
  wire  _T_17559; // @[Mux.scala 46:19:@15095.4]
  wire [7:0] _T_17560; // @[Mux.scala 46:16:@15096.4]
  wire  _T_17561; // @[Mux.scala 46:19:@15097.4]
  wire [7:0] _T_17562; // @[Mux.scala 46:16:@15098.4]
  wire  _T_17563; // @[Mux.scala 46:19:@15099.4]
  wire [7:0] _T_17564; // @[Mux.scala 46:16:@15100.4]
  wire  _T_17565; // @[Mux.scala 46:19:@15101.4]
  wire [7:0] _T_17566; // @[Mux.scala 46:16:@15102.4]
  wire  _T_17567; // @[Mux.scala 46:19:@15103.4]
  wire [7:0] _T_17568; // @[Mux.scala 46:16:@15104.4]
  wire  _T_17569; // @[Mux.scala 46:19:@15105.4]
  wire [7:0] _T_17570; // @[Mux.scala 46:16:@15106.4]
  wire  _T_17571; // @[Mux.scala 46:19:@15107.4]
  wire [7:0] _T_17572; // @[Mux.scala 46:16:@15108.4]
  wire  _T_17573; // @[Mux.scala 46:19:@15109.4]
  wire [7:0] _T_17574; // @[Mux.scala 46:16:@15110.4]
  wire  _T_17575; // @[Mux.scala 46:19:@15111.4]
  wire [7:0] _T_17576; // @[Mux.scala 46:16:@15112.4]
  wire  _T_17577; // @[Mux.scala 46:19:@15113.4]
  wire [7:0] _T_17578; // @[Mux.scala 46:16:@15114.4]
  wire  _T_17579; // @[Mux.scala 46:19:@15115.4]
  wire [7:0] _T_17580; // @[Mux.scala 46:16:@15116.4]
  wire  _T_17581; // @[Mux.scala 46:19:@15117.4]
  wire [7:0] _T_17582; // @[Mux.scala 46:16:@15118.4]
  wire  _T_17583; // @[Mux.scala 46:19:@15119.4]
  wire [7:0] _T_17584; // @[Mux.scala 46:16:@15120.4]
  wire  _T_17585; // @[Mux.scala 46:19:@15121.4]
  wire [7:0] _T_17586; // @[Mux.scala 46:16:@15122.4]
  wire  _T_17587; // @[Mux.scala 46:19:@15123.4]
  wire [7:0] _T_17588; // @[Mux.scala 46:16:@15124.4]
  wire  _T_17589; // @[Mux.scala 46:19:@15125.4]
  wire [7:0] _T_17590; // @[Mux.scala 46:16:@15126.4]
  wire  _T_17591; // @[Mux.scala 46:19:@15127.4]
  wire [7:0] _T_17592; // @[Mux.scala 46:16:@15128.4]
  wire  _T_17593; // @[Mux.scala 46:19:@15129.4]
  wire [7:0] _T_17594; // @[Mux.scala 46:16:@15130.4]
  wire  _T_17595; // @[Mux.scala 46:19:@15131.4]
  wire [7:0] _T_17596; // @[Mux.scala 46:16:@15132.4]
  wire  _T_17597; // @[Mux.scala 46:19:@15133.4]
  wire [7:0] _T_17598; // @[Mux.scala 46:16:@15134.4]
  wire  _T_17599; // @[Mux.scala 46:19:@15135.4]
  wire [7:0] _T_17600; // @[Mux.scala 46:16:@15136.4]
  wire  _T_17601; // @[Mux.scala 46:19:@15137.4]
  wire [7:0] _T_17602; // @[Mux.scala 46:16:@15138.4]
  wire  _T_17603; // @[Mux.scala 46:19:@15139.4]
  wire [7:0] _T_17604; // @[Mux.scala 46:16:@15140.4]
  wire  _T_17605; // @[Mux.scala 46:19:@15141.4]
  wire [7:0] _T_17606; // @[Mux.scala 46:16:@15142.4]
  wire  _T_17607; // @[Mux.scala 46:19:@15143.4]
  wire [7:0] _T_17608; // @[Mux.scala 46:16:@15144.4]
  wire  _T_17609; // @[Mux.scala 46:19:@15145.4]
  wire [7:0] _T_17610; // @[Mux.scala 46:16:@15146.4]
  wire  _T_17611; // @[Mux.scala 46:19:@15147.4]
  wire [7:0] _T_17612; // @[Mux.scala 46:16:@15148.4]
  wire  _T_17613; // @[Mux.scala 46:19:@15149.4]
  wire [7:0] _T_17614; // @[Mux.scala 46:16:@15150.4]
  wire  _T_17615; // @[Mux.scala 46:19:@15151.4]
  wire [7:0] _T_17616; // @[Mux.scala 46:16:@15152.4]
  wire  _T_17617; // @[Mux.scala 46:19:@15153.4]
  wire [7:0] _T_17618; // @[Mux.scala 46:16:@15154.4]
  wire  _T_17619; // @[Mux.scala 46:19:@15155.4]
  wire [7:0] _T_17620; // @[Mux.scala 46:16:@15156.4]
  wire  _T_17621; // @[Mux.scala 46:19:@15157.4]
  wire [7:0] _T_17622; // @[Mux.scala 46:16:@15158.4]
  wire  _T_17623; // @[Mux.scala 46:19:@15159.4]
  wire [7:0] _T_17624; // @[Mux.scala 46:16:@15160.4]
  wire  _T_17625; // @[Mux.scala 46:19:@15161.4]
  wire [7:0] _T_17626; // @[Mux.scala 46:16:@15162.4]
  wire  _T_17692; // @[Mux.scala 46:19:@15164.4]
  wire [7:0] _T_17693; // @[Mux.scala 46:16:@15165.4]
  wire  _T_17694; // @[Mux.scala 46:19:@15166.4]
  wire [7:0] _T_17695; // @[Mux.scala 46:16:@15167.4]
  wire  _T_17696; // @[Mux.scala 46:19:@15168.4]
  wire [7:0] _T_17697; // @[Mux.scala 46:16:@15169.4]
  wire  _T_17698; // @[Mux.scala 46:19:@15170.4]
  wire [7:0] _T_17699; // @[Mux.scala 46:16:@15171.4]
  wire  _T_17700; // @[Mux.scala 46:19:@15172.4]
  wire [7:0] _T_17701; // @[Mux.scala 46:16:@15173.4]
  wire  _T_17702; // @[Mux.scala 46:19:@15174.4]
  wire [7:0] _T_17703; // @[Mux.scala 46:16:@15175.4]
  wire  _T_17704; // @[Mux.scala 46:19:@15176.4]
  wire [7:0] _T_17705; // @[Mux.scala 46:16:@15177.4]
  wire  _T_17706; // @[Mux.scala 46:19:@15178.4]
  wire [7:0] _T_17707; // @[Mux.scala 46:16:@15179.4]
  wire  _T_17708; // @[Mux.scala 46:19:@15180.4]
  wire [7:0] _T_17709; // @[Mux.scala 46:16:@15181.4]
  wire  _T_17710; // @[Mux.scala 46:19:@15182.4]
  wire [7:0] _T_17711; // @[Mux.scala 46:16:@15183.4]
  wire  _T_17712; // @[Mux.scala 46:19:@15184.4]
  wire [7:0] _T_17713; // @[Mux.scala 46:16:@15185.4]
  wire  _T_17714; // @[Mux.scala 46:19:@15186.4]
  wire [7:0] _T_17715; // @[Mux.scala 46:16:@15187.4]
  wire  _T_17716; // @[Mux.scala 46:19:@15188.4]
  wire [7:0] _T_17717; // @[Mux.scala 46:16:@15189.4]
  wire  _T_17718; // @[Mux.scala 46:19:@15190.4]
  wire [7:0] _T_17719; // @[Mux.scala 46:16:@15191.4]
  wire  _T_17720; // @[Mux.scala 46:19:@15192.4]
  wire [7:0] _T_17721; // @[Mux.scala 46:16:@15193.4]
  wire  _T_17722; // @[Mux.scala 46:19:@15194.4]
  wire [7:0] _T_17723; // @[Mux.scala 46:16:@15195.4]
  wire  _T_17724; // @[Mux.scala 46:19:@15196.4]
  wire [7:0] _T_17725; // @[Mux.scala 46:16:@15197.4]
  wire  _T_17726; // @[Mux.scala 46:19:@15198.4]
  wire [7:0] _T_17727; // @[Mux.scala 46:16:@15199.4]
  wire  _T_17728; // @[Mux.scala 46:19:@15200.4]
  wire [7:0] _T_17729; // @[Mux.scala 46:16:@15201.4]
  wire  _T_17730; // @[Mux.scala 46:19:@15202.4]
  wire [7:0] _T_17731; // @[Mux.scala 46:16:@15203.4]
  wire  _T_17732; // @[Mux.scala 46:19:@15204.4]
  wire [7:0] _T_17733; // @[Mux.scala 46:16:@15205.4]
  wire  _T_17734; // @[Mux.scala 46:19:@15206.4]
  wire [7:0] _T_17735; // @[Mux.scala 46:16:@15207.4]
  wire  _T_17736; // @[Mux.scala 46:19:@15208.4]
  wire [7:0] _T_17737; // @[Mux.scala 46:16:@15209.4]
  wire  _T_17738; // @[Mux.scala 46:19:@15210.4]
  wire [7:0] _T_17739; // @[Mux.scala 46:16:@15211.4]
  wire  _T_17740; // @[Mux.scala 46:19:@15212.4]
  wire [7:0] _T_17741; // @[Mux.scala 46:16:@15213.4]
  wire  _T_17742; // @[Mux.scala 46:19:@15214.4]
  wire [7:0] _T_17743; // @[Mux.scala 46:16:@15215.4]
  wire  _T_17744; // @[Mux.scala 46:19:@15216.4]
  wire [7:0] _T_17745; // @[Mux.scala 46:16:@15217.4]
  wire  _T_17746; // @[Mux.scala 46:19:@15218.4]
  wire [7:0] _T_17747; // @[Mux.scala 46:16:@15219.4]
  wire  _T_17748; // @[Mux.scala 46:19:@15220.4]
  wire [7:0] _T_17749; // @[Mux.scala 46:16:@15221.4]
  wire  _T_17750; // @[Mux.scala 46:19:@15222.4]
  wire [7:0] _T_17751; // @[Mux.scala 46:16:@15223.4]
  wire  _T_17752; // @[Mux.scala 46:19:@15224.4]
  wire [7:0] _T_17753; // @[Mux.scala 46:16:@15225.4]
  wire  _T_17754; // @[Mux.scala 46:19:@15226.4]
  wire [7:0] _T_17755; // @[Mux.scala 46:16:@15227.4]
  wire  _T_17756; // @[Mux.scala 46:19:@15228.4]
  wire [7:0] _T_17757; // @[Mux.scala 46:16:@15229.4]
  wire  _T_17758; // @[Mux.scala 46:19:@15230.4]
  wire [7:0] _T_17759; // @[Mux.scala 46:16:@15231.4]
  wire  _T_17760; // @[Mux.scala 46:19:@15232.4]
  wire [7:0] _T_17761; // @[Mux.scala 46:16:@15233.4]
  wire  _T_17762; // @[Mux.scala 46:19:@15234.4]
  wire [7:0] _T_17763; // @[Mux.scala 46:16:@15235.4]
  wire  _T_17764; // @[Mux.scala 46:19:@15236.4]
  wire [7:0] _T_17765; // @[Mux.scala 46:16:@15237.4]
  wire  _T_17766; // @[Mux.scala 46:19:@15238.4]
  wire [7:0] _T_17767; // @[Mux.scala 46:16:@15239.4]
  wire  _T_17768; // @[Mux.scala 46:19:@15240.4]
  wire [7:0] _T_17769; // @[Mux.scala 46:16:@15241.4]
  wire  _T_17770; // @[Mux.scala 46:19:@15242.4]
  wire [7:0] _T_17771; // @[Mux.scala 46:16:@15243.4]
  wire  _T_17772; // @[Mux.scala 46:19:@15244.4]
  wire [7:0] _T_17773; // @[Mux.scala 46:16:@15245.4]
  wire  _T_17774; // @[Mux.scala 46:19:@15246.4]
  wire [7:0] _T_17775; // @[Mux.scala 46:16:@15247.4]
  wire  _T_17776; // @[Mux.scala 46:19:@15248.4]
  wire [7:0] _T_17777; // @[Mux.scala 46:16:@15249.4]
  wire  _T_17778; // @[Mux.scala 46:19:@15250.4]
  wire [7:0] _T_17779; // @[Mux.scala 46:16:@15251.4]
  wire  _T_17780; // @[Mux.scala 46:19:@15252.4]
  wire [7:0] _T_17781; // @[Mux.scala 46:16:@15253.4]
  wire  _T_17782; // @[Mux.scala 46:19:@15254.4]
  wire [7:0] _T_17783; // @[Mux.scala 46:16:@15255.4]
  wire  _T_17784; // @[Mux.scala 46:19:@15256.4]
  wire [7:0] _T_17785; // @[Mux.scala 46:16:@15257.4]
  wire  _T_17786; // @[Mux.scala 46:19:@15258.4]
  wire [7:0] _T_17787; // @[Mux.scala 46:16:@15259.4]
  wire  _T_17788; // @[Mux.scala 46:19:@15260.4]
  wire [7:0] _T_17789; // @[Mux.scala 46:16:@15261.4]
  wire  _T_17790; // @[Mux.scala 46:19:@15262.4]
  wire [7:0] _T_17791; // @[Mux.scala 46:16:@15263.4]
  wire  _T_17792; // @[Mux.scala 46:19:@15264.4]
  wire [7:0] _T_17793; // @[Mux.scala 46:16:@15265.4]
  wire  _T_17794; // @[Mux.scala 46:19:@15266.4]
  wire [7:0] _T_17795; // @[Mux.scala 46:16:@15267.4]
  wire  _T_17796; // @[Mux.scala 46:19:@15268.4]
  wire [7:0] _T_17797; // @[Mux.scala 46:16:@15269.4]
  wire  _T_17798; // @[Mux.scala 46:19:@15270.4]
  wire [7:0] _T_17799; // @[Mux.scala 46:16:@15271.4]
  wire  _T_17800; // @[Mux.scala 46:19:@15272.4]
  wire [7:0] _T_17801; // @[Mux.scala 46:16:@15273.4]
  wire  _T_17802; // @[Mux.scala 46:19:@15274.4]
  wire [7:0] _T_17803; // @[Mux.scala 46:16:@15275.4]
  wire  _T_17804; // @[Mux.scala 46:19:@15276.4]
  wire [7:0] _T_17805; // @[Mux.scala 46:16:@15277.4]
  wire  _T_17806; // @[Mux.scala 46:19:@15278.4]
  wire [7:0] _T_17807; // @[Mux.scala 46:16:@15279.4]
  wire  _T_17808; // @[Mux.scala 46:19:@15280.4]
  wire [7:0] _T_17809; // @[Mux.scala 46:16:@15281.4]
  wire  _T_17810; // @[Mux.scala 46:19:@15282.4]
  wire [7:0] _T_17811; // @[Mux.scala 46:16:@15283.4]
  wire  _T_17812; // @[Mux.scala 46:19:@15284.4]
  wire [7:0] _T_17813; // @[Mux.scala 46:16:@15285.4]
  wire  _T_17814; // @[Mux.scala 46:19:@15286.4]
  wire [7:0] _T_17815; // @[Mux.scala 46:16:@15287.4]
  wire  _T_17816; // @[Mux.scala 46:19:@15288.4]
  wire [7:0] _T_17817; // @[Mux.scala 46:16:@15289.4]
  wire  _T_17818; // @[Mux.scala 46:19:@15290.4]
  wire [7:0] _T_17819; // @[Mux.scala 46:16:@15291.4]
  reg  _T_17822; // @[NV_NVDLA_CSC_WL_dec.scala 94:27:@15293.4]
  reg [31:0] _RAND_225;
  reg  _T_17961_0; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_226;
  reg  _T_17961_1; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_227;
  reg  _T_17961_2; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_228;
  reg  _T_17961_3; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_229;
  reg  _T_17961_4; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_230;
  reg  _T_17961_5; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_231;
  reg  _T_17961_6; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_232;
  reg  _T_17961_7; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_233;
  reg  _T_17961_8; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_234;
  reg  _T_17961_9; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_235;
  reg  _T_17961_10; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_236;
  reg  _T_17961_11; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_237;
  reg  _T_17961_12; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_238;
  reg  _T_17961_13; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_239;
  reg  _T_17961_14; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_240;
  reg  _T_17961_15; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_241;
  reg  _T_17961_16; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_242;
  reg  _T_17961_17; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_243;
  reg  _T_17961_18; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_244;
  reg  _T_17961_19; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_245;
  reg  _T_17961_20; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_246;
  reg  _T_17961_21; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_247;
  reg  _T_17961_22; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_248;
  reg  _T_17961_23; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_249;
  reg  _T_17961_24; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_250;
  reg  _T_17961_25; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_251;
  reg  _T_17961_26; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_252;
  reg  _T_17961_27; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_253;
  reg  _T_17961_28; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_254;
  reg  _T_17961_29; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_255;
  reg  _T_17961_30; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_256;
  reg  _T_17961_31; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@15327.4]
  reg [31:0] _RAND_257;
  reg [7:0] _T_18065_0; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_258;
  reg [7:0] _T_18065_1; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_259;
  reg [7:0] _T_18065_2; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_260;
  reg [7:0] _T_18065_3; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_261;
  reg [7:0] _T_18065_4; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_262;
  reg [7:0] _T_18065_5; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_263;
  reg [7:0] _T_18065_6; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_264;
  reg [7:0] _T_18065_7; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_265;
  reg [7:0] _T_18065_8; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_266;
  reg [7:0] _T_18065_9; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_267;
  reg [7:0] _T_18065_10; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_268;
  reg [7:0] _T_18065_11; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_269;
  reg [7:0] _T_18065_12; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_270;
  reg [7:0] _T_18065_13; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_271;
  reg [7:0] _T_18065_14; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_272;
  reg [7:0] _T_18065_15; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_273;
  reg [7:0] _T_18065_16; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_274;
  reg [7:0] _T_18065_17; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_275;
  reg [7:0] _T_18065_18; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_276;
  reg [7:0] _T_18065_19; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_277;
  reg [7:0] _T_18065_20; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_278;
  reg [7:0] _T_18065_21; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_279;
  reg [7:0] _T_18065_22; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_280;
  reg [7:0] _T_18065_23; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_281;
  reg [7:0] _T_18065_24; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_282;
  reg [7:0] _T_18065_25; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_283;
  reg [7:0] _T_18065_26; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_284;
  reg [7:0] _T_18065_27; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_285;
  reg [7:0] _T_18065_28; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_286;
  reg [7:0] _T_18065_29; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_287;
  reg [7:0] _T_18065_30; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_288;
  reg [7:0] _T_18065_31; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_289;
  reg [7:0] _T_18065_32; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_290;
  reg [7:0] _T_18065_33; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_291;
  reg [7:0] _T_18065_34; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_292;
  reg [7:0] _T_18065_35; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_293;
  reg [7:0] _T_18065_36; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_294;
  reg [7:0] _T_18065_37; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_295;
  reg [7:0] _T_18065_38; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_296;
  reg [7:0] _T_18065_39; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_297;
  reg [7:0] _T_18065_40; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_298;
  reg [7:0] _T_18065_41; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_299;
  reg [7:0] _T_18065_42; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_300;
  reg [7:0] _T_18065_43; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_301;
  reg [7:0] _T_18065_44; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_302;
  reg [7:0] _T_18065_45; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_303;
  reg [7:0] _T_18065_46; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_304;
  reg [7:0] _T_18065_47; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_305;
  reg [7:0] _T_18065_48; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_306;
  reg [7:0] _T_18065_49; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_307;
  reg [7:0] _T_18065_50; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_308;
  reg [7:0] _T_18065_51; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_309;
  reg [7:0] _T_18065_52; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_310;
  reg [7:0] _T_18065_53; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_311;
  reg [7:0] _T_18065_54; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_312;
  reg [7:0] _T_18065_55; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_313;
  reg [7:0] _T_18065_56; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_314;
  reg [7:0] _T_18065_57; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_315;
  reg [7:0] _T_18065_58; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_316;
  reg [7:0] _T_18065_59; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_317;
  reg [7:0] _T_18065_60; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_318;
  reg [7:0] _T_18065_61; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_319;
  reg [7:0] _T_18065_62; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_320;
  reg [7:0] _T_18065_63; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@15328.4]
  reg [31:0] _RAND_321;
  wire  _GEN_224; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_225; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_226; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_227; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_228; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_229; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_230; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_231; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_232; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_233; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_234; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_235; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_236; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_237; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_238; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_239; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_240; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_241; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_242; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_243; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_244; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_245; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_246; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_247; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_248; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_249; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_250; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_251; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_252; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_253; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_254; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire  _GEN_255; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  wire [7:0] _GEN_256; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15365.6]
  wire [7:0] _GEN_258; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15373.6]
  wire [7:0] _GEN_260; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15381.6]
  wire [7:0] _GEN_262; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15389.6]
  wire [7:0] _GEN_264; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15397.6]
  wire [7:0] _GEN_266; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15405.6]
  wire [7:0] _GEN_268; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15413.6]
  wire [7:0] _GEN_270; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15421.6]
  wire [7:0] _GEN_272; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15429.6]
  wire [7:0] _GEN_274; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15437.6]
  wire [7:0] _GEN_276; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15445.6]
  wire [7:0] _GEN_278; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15453.6]
  wire [7:0] _GEN_280; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15461.6]
  wire [7:0] _GEN_282; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15469.6]
  wire [7:0] _GEN_284; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15477.6]
  wire [7:0] _GEN_286; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15485.6]
  wire [7:0] _GEN_288; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15493.6]
  wire [7:0] _GEN_290; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15501.6]
  wire [7:0] _GEN_292; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15509.6]
  wire [7:0] _GEN_294; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15517.6]
  wire [7:0] _GEN_296; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15525.6]
  wire [7:0] _GEN_298; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15533.6]
  wire [7:0] _GEN_300; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15541.6]
  wire [7:0] _GEN_302; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15549.6]
  wire [7:0] _GEN_304; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15557.6]
  wire [7:0] _GEN_306; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15565.6]
  wire [7:0] _GEN_308; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15573.6]
  wire [7:0] _GEN_310; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15581.6]
  wire [7:0] _GEN_312; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15589.6]
  wire [7:0] _GEN_314; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15597.6]
  wire [7:0] _GEN_316; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15605.6]
  wire [7:0] _GEN_318; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15613.6]
  wire [7:0] _GEN_320; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15621.6]
  wire [7:0] _GEN_322; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15629.6]
  wire [7:0] _GEN_324; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15637.6]
  wire [7:0] _GEN_326; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15645.6]
  wire [7:0] _GEN_328; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15653.6]
  wire [7:0] _GEN_330; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15661.6]
  wire [7:0] _GEN_332; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15669.6]
  wire [7:0] _GEN_334; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15677.6]
  wire [7:0] _GEN_336; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15685.6]
  wire [7:0] _GEN_338; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15693.6]
  wire [7:0] _GEN_340; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15701.6]
  wire [7:0] _GEN_342; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15709.6]
  wire [7:0] _GEN_344; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15717.6]
  wire [7:0] _GEN_346; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15725.6]
  wire [7:0] _GEN_348; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15733.6]
  wire [7:0] _GEN_350; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15741.6]
  wire [7:0] _GEN_352; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15749.6]
  wire [7:0] _GEN_354; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15757.6]
  wire [7:0] _GEN_356; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15765.6]
  wire [7:0] _GEN_358; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15773.6]
  wire [7:0] _GEN_360; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15781.6]
  wire [7:0] _GEN_362; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15789.6]
  wire [7:0] _GEN_364; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15797.6]
  wire [7:0] _GEN_366; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15805.6]
  wire [7:0] _GEN_368; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15813.6]
  wire [7:0] _GEN_370; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15821.6]
  wire [7:0] _GEN_372; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15829.6]
  wire [7:0] _GEN_374; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15837.6]
  wire [7:0] _GEN_376; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15845.6]
  wire [7:0] _GEN_378; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15853.6]
  wire [7:0] _GEN_380; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15861.6]
  wire [7:0] _GEN_382; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15869.6]
  wire  _T_18267; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15877.4]
  wire  _T_18269; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15879.4]
  wire  _T_18271; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15881.4]
  wire  _T_18273; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15883.4]
  wire  _T_18275; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15885.4]
  wire  _T_18277; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15887.4]
  wire  _T_18279; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15889.4]
  wire  _T_18281; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15891.4]
  wire  _T_18283; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15893.4]
  wire  _T_18285; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15895.4]
  wire  _T_18287; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15897.4]
  wire  _T_18289; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15899.4]
  wire  _T_18291; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15901.4]
  wire  _T_18293; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15903.4]
  wire  _T_18295; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15905.4]
  wire  _T_18297; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15907.4]
  wire  _T_18299; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15909.4]
  wire  _T_18301; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15911.4]
  wire  _T_18303; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15913.4]
  wire  _T_18305; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15915.4]
  wire  _T_18307; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15917.4]
  wire  _T_18309; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15919.4]
  wire  _T_18311; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15921.4]
  wire  _T_18313; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15923.4]
  wire  _T_18315; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15925.4]
  wire  _T_18317; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15927.4]
  wire  _T_18319; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15929.4]
  wire  _T_18321; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15931.4]
  wire  _T_18323; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15933.4]
  wire  _T_18325; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15935.4]
  wire  _T_18327; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15937.4]
  wire  _T_18329; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15939.4]
  wire  _T_18331; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15941.4]
  wire  _T_18333; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15943.4]
  wire  _T_18335; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15945.4]
  wire  _T_18337; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15947.4]
  wire  _T_18339; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15949.4]
  wire  _T_18341; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15951.4]
  wire  _T_18343; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15953.4]
  wire  _T_18345; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15955.4]
  wire  _T_18347; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15957.4]
  wire  _T_18349; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15959.4]
  wire  _T_18351; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15961.4]
  wire  _T_18353; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15963.4]
  wire  _T_18355; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15965.4]
  wire  _T_18357; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15967.4]
  wire  _T_18359; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15969.4]
  wire  _T_18361; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15971.4]
  wire  _T_18363; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15973.4]
  wire  _T_18365; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15975.4]
  wire  _T_18367; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15977.4]
  wire  _T_18369; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15979.4]
  wire  _T_18371; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15981.4]
  wire  _T_18373; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15983.4]
  wire  _T_18375; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15985.4]
  wire  _T_18377; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15987.4]
  wire  _T_18379; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15989.4]
  wire  _T_18381; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15991.4]
  wire  _T_18383; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15993.4]
  wire  _T_18385; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15995.4]
  wire  _T_18387; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15997.4]
  wire  _T_18389; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15999.4]
  wire  _T_18391; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@16001.4]
  wire  _T_18393; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@16003.4]
  reg  _T_18396; // @[NV_NVDLA_CSC_WL_dec.scala 122:27:@16005.4]
  reg [31:0] _RAND_322;
  reg  _T_18400_0; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_323;
  reg  _T_18400_1; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_324;
  reg  _T_18400_2; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_325;
  reg  _T_18400_3; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_326;
  reg  _T_18400_4; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_327;
  reg  _T_18400_5; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_328;
  reg  _T_18400_6; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_329;
  reg  _T_18400_7; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_330;
  reg  _T_18400_8; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_331;
  reg  _T_18400_9; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_332;
  reg  _T_18400_10; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_333;
  reg  _T_18400_11; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_334;
  reg  _T_18400_12; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_335;
  reg  _T_18400_13; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_336;
  reg  _T_18400_14; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_337;
  reg  _T_18400_15; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_338;
  reg  _T_18400_16; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_339;
  reg  _T_18400_17; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_340;
  reg  _T_18400_18; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_341;
  reg  _T_18400_19; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_342;
  reg  _T_18400_20; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_343;
  reg  _T_18400_21; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_344;
  reg  _T_18400_22; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_345;
  reg  _T_18400_23; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_346;
  reg  _T_18400_24; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_347;
  reg  _T_18400_25; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_348;
  reg  _T_18400_26; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_349;
  reg  _T_18400_27; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_350;
  reg  _T_18400_28; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_351;
  reg  _T_18400_29; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_352;
  reg  _T_18400_30; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_353;
  reg  _T_18400_31; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_354;
  reg  _T_18400_32; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_355;
  reg  _T_18400_33; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_356;
  reg  _T_18400_34; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_357;
  reg  _T_18400_35; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_358;
  reg  _T_18400_36; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_359;
  reg  _T_18400_37; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_360;
  reg  _T_18400_38; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_361;
  reg  _T_18400_39; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_362;
  reg  _T_18400_40; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_363;
  reg  _T_18400_41; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_364;
  reg  _T_18400_42; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_365;
  reg  _T_18400_43; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_366;
  reg  _T_18400_44; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_367;
  reg  _T_18400_45; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_368;
  reg  _T_18400_46; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_369;
  reg  _T_18400_47; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_370;
  reg  _T_18400_48; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_371;
  reg  _T_18400_49; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_372;
  reg  _T_18400_50; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_373;
  reg  _T_18400_51; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_374;
  reg  _T_18400_52; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_375;
  reg  _T_18400_53; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_376;
  reg  _T_18400_54; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_377;
  reg  _T_18400_55; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_378;
  reg  _T_18400_56; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_379;
  reg  _T_18400_57; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_380;
  reg  _T_18400_58; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_381;
  reg  _T_18400_59; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_382;
  reg  _T_18400_60; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_383;
  reg  _T_18400_61; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_384;
  reg  _T_18400_62; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_385;
  reg  _T_18400_63; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@16006.4]
  reg [31:0] _RAND_386;
  reg  _T_18605_0; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_387;
  reg  _T_18605_1; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_388;
  reg  _T_18605_2; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_389;
  reg  _T_18605_3; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_390;
  reg  _T_18605_4; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_391;
  reg  _T_18605_5; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_392;
  reg  _T_18605_6; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_393;
  reg  _T_18605_7; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_394;
  reg  _T_18605_8; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_395;
  reg  _T_18605_9; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_396;
  reg  _T_18605_10; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_397;
  reg  _T_18605_11; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_398;
  reg  _T_18605_12; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_399;
  reg  _T_18605_13; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_400;
  reg  _T_18605_14; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_401;
  reg  _T_18605_15; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_402;
  reg  _T_18605_16; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_403;
  reg  _T_18605_17; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_404;
  reg  _T_18605_18; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_405;
  reg  _T_18605_19; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_406;
  reg  _T_18605_20; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_407;
  reg  _T_18605_21; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_408;
  reg  _T_18605_22; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_409;
  reg  _T_18605_23; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_410;
  reg  _T_18605_24; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_411;
  reg  _T_18605_25; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_412;
  reg  _T_18605_26; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_413;
  reg  _T_18605_27; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_414;
  reg  _T_18605_28; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_415;
  reg  _T_18605_29; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_416;
  reg  _T_18605_30; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_417;
  reg  _T_18605_31; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@16040.4]
  reg [31:0] _RAND_418;
  reg [7:0] _T_18709_0; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_419;
  reg [7:0] _T_18709_1; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_420;
  reg [7:0] _T_18709_2; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_421;
  reg [7:0] _T_18709_3; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_422;
  reg [7:0] _T_18709_4; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_423;
  reg [7:0] _T_18709_5; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_424;
  reg [7:0] _T_18709_6; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_425;
  reg [7:0] _T_18709_7; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_426;
  reg [7:0] _T_18709_8; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_427;
  reg [7:0] _T_18709_9; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_428;
  reg [7:0] _T_18709_10; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_429;
  reg [7:0] _T_18709_11; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_430;
  reg [7:0] _T_18709_12; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_431;
  reg [7:0] _T_18709_13; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_432;
  reg [7:0] _T_18709_14; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_433;
  reg [7:0] _T_18709_15; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_434;
  reg [7:0] _T_18709_16; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_435;
  reg [7:0] _T_18709_17; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_436;
  reg [7:0] _T_18709_18; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_437;
  reg [7:0] _T_18709_19; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_438;
  reg [7:0] _T_18709_20; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_439;
  reg [7:0] _T_18709_21; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_440;
  reg [7:0] _T_18709_22; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_441;
  reg [7:0] _T_18709_23; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_442;
  reg [7:0] _T_18709_24; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_443;
  reg [7:0] _T_18709_25; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_444;
  reg [7:0] _T_18709_26; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_445;
  reg [7:0] _T_18709_27; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_446;
  reg [7:0] _T_18709_28; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_447;
  reg [7:0] _T_18709_29; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_448;
  reg [7:0] _T_18709_30; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_449;
  reg [7:0] _T_18709_31; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_450;
  reg [7:0] _T_18709_32; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_451;
  reg [7:0] _T_18709_33; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_452;
  reg [7:0] _T_18709_34; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_453;
  reg [7:0] _T_18709_35; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_454;
  reg [7:0] _T_18709_36; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_455;
  reg [7:0] _T_18709_37; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_456;
  reg [7:0] _T_18709_38; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_457;
  reg [7:0] _T_18709_39; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_458;
  reg [7:0] _T_18709_40; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_459;
  reg [7:0] _T_18709_41; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_460;
  reg [7:0] _T_18709_42; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_461;
  reg [7:0] _T_18709_43; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_462;
  reg [7:0] _T_18709_44; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_463;
  reg [7:0] _T_18709_45; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_464;
  reg [7:0] _T_18709_46; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_465;
  reg [7:0] _T_18709_47; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_466;
  reg [7:0] _T_18709_48; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_467;
  reg [7:0] _T_18709_49; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_468;
  reg [7:0] _T_18709_50; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_469;
  reg [7:0] _T_18709_51; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_470;
  reg [7:0] _T_18709_52; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_471;
  reg [7:0] _T_18709_53; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_472;
  reg [7:0] _T_18709_54; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_473;
  reg [7:0] _T_18709_55; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_474;
  reg [7:0] _T_18709_56; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_475;
  reg [7:0] _T_18709_57; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_476;
  reg [7:0] _T_18709_58; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_477;
  reg [7:0] _T_18709_59; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_478;
  reg [7:0] _T_18709_60; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_479;
  reg [7:0] _T_18709_61; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_480;
  reg [7:0] _T_18709_62; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_481;
  reg [7:0] _T_18709_63; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@16041.4]
  reg [31:0] _RAND_482;
  wire  _GEN_448; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_449; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_450; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_451; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_452; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_453; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_454; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_455; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_456; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_457; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_458; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_459; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_460; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_461; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_462; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_463; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_464; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_465; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_466; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_467; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_468; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_469; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_470; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_471; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_472; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_473; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_474; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_475; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_476; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_477; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_478; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  wire  _GEN_479; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _T_1771 = io_input_mask_en[8]; // @[NV_NVDLA_CSC_WL_dec.scala 56:48:@2095.4]
  assign _T_1906_0 = _T_1771 ? io_input_bits_mask_0 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_1 = _T_1771 ? io_input_bits_mask_1 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_2 = _T_1771 ? io_input_bits_mask_2 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_3 = _T_1771 ? io_input_bits_mask_3 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_4 = _T_1771 ? io_input_bits_mask_4 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_5 = _T_1771 ? io_input_bits_mask_5 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_6 = _T_1771 ? io_input_bits_mask_6 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_7 = _T_1771 ? io_input_bits_mask_7 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_8 = _T_1771 ? io_input_bits_mask_8 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_9 = _T_1771 ? io_input_bits_mask_9 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_10 = _T_1771 ? io_input_bits_mask_10 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_11 = _T_1771 ? io_input_bits_mask_11 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_12 = _T_1771 ? io_input_bits_mask_12 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_13 = _T_1771 ? io_input_bits_mask_13 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_14 = _T_1771 ? io_input_bits_mask_14 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_15 = _T_1771 ? io_input_bits_mask_15 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_16 = _T_1771 ? io_input_bits_mask_16 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_17 = _T_1771 ? io_input_bits_mask_17 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_18 = _T_1771 ? io_input_bits_mask_18 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_19 = _T_1771 ? io_input_bits_mask_19 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_20 = _T_1771 ? io_input_bits_mask_20 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_21 = _T_1771 ? io_input_bits_mask_21 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_22 = _T_1771 ? io_input_bits_mask_22 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_23 = _T_1771 ? io_input_bits_mask_23 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_24 = _T_1771 ? io_input_bits_mask_24 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_25 = _T_1771 ? io_input_bits_mask_25 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_26 = _T_1771 ? io_input_bits_mask_26 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_27 = _T_1771 ? io_input_bits_mask_27 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_28 = _T_1771 ? io_input_bits_mask_28 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_29 = _T_1771 ? io_input_bits_mask_29 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_30 = _T_1771 ? io_input_bits_mask_30 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_31 = _T_1771 ? io_input_bits_mask_31 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_32 = _T_1771 ? io_input_bits_mask_32 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_33 = _T_1771 ? io_input_bits_mask_33 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_34 = _T_1771 ? io_input_bits_mask_34 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_35 = _T_1771 ? io_input_bits_mask_35 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_36 = _T_1771 ? io_input_bits_mask_36 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_37 = _T_1771 ? io_input_bits_mask_37 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_38 = _T_1771 ? io_input_bits_mask_38 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_39 = _T_1771 ? io_input_bits_mask_39 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_40 = _T_1771 ? io_input_bits_mask_40 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_41 = _T_1771 ? io_input_bits_mask_41 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_42 = _T_1771 ? io_input_bits_mask_42 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_43 = _T_1771 ? io_input_bits_mask_43 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_44 = _T_1771 ? io_input_bits_mask_44 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_45 = _T_1771 ? io_input_bits_mask_45 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_46 = _T_1771 ? io_input_bits_mask_46 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_47 = _T_1771 ? io_input_bits_mask_47 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_48 = _T_1771 ? io_input_bits_mask_48 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_49 = _T_1771 ? io_input_bits_mask_49 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_50 = _T_1771 ? io_input_bits_mask_50 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_51 = _T_1771 ? io_input_bits_mask_51 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_52 = _T_1771 ? io_input_bits_mask_52 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_53 = _T_1771 ? io_input_bits_mask_53 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_54 = _T_1771 ? io_input_bits_mask_54 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_55 = _T_1771 ? io_input_bits_mask_55 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_56 = _T_1771 ? io_input_bits_mask_56 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_57 = _T_1771 ? io_input_bits_mask_57 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_58 = _T_1771 ? io_input_bits_mask_58 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_59 = _T_1771 ? io_input_bits_mask_59 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_60 = _T_1771 ? io_input_bits_mask_60 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_61 = _T_1771 ? io_input_bits_mask_61 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_62 = _T_1771 ? io_input_bits_mask_62 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_1906_63 = _T_1771 ? io_input_bits_mask_63 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@2161.4]
  assign _T_2174 = {_T_1906_7,_T_1906_6,_T_1906_5,_T_1906_4,_T_1906_3,_T_1906_2,_T_1906_1,_T_1906_0}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2169.4]
  assign _T_2182 = {_T_1906_15,_T_1906_14,_T_1906_13,_T_1906_12,_T_1906_11,_T_1906_10,_T_1906_9,_T_1906_8,_T_2174}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2177.4]
  assign _T_2189 = {_T_1906_23,_T_1906_22,_T_1906_21,_T_1906_20,_T_1906_19,_T_1906_18,_T_1906_17,_T_1906_16}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2184.4]
  assign _T_2198 = {_T_1906_31,_T_1906_30,_T_1906_29,_T_1906_28,_T_1906_27,_T_1906_26,_T_1906_25,_T_1906_24,_T_2189,_T_2182}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2193.4]
  assign _T_2205 = {_T_1906_39,_T_1906_38,_T_1906_37,_T_1906_36,_T_1906_35,_T_1906_34,_T_1906_33,_T_1906_32}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2200.4]
  assign _T_2213 = {_T_1906_47,_T_1906_46,_T_1906_45,_T_1906_44,_T_1906_43,_T_1906_42,_T_1906_41,_T_1906_40,_T_2205}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2208.4]
  assign _T_2220 = {_T_1906_55,_T_1906_54,_T_1906_53,_T_1906_52,_T_1906_51,_T_1906_50,_T_1906_49,_T_1906_48}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2215.4]
  assign _T_2229 = {_T_1906_63,_T_1906_62,_T_1906_61,_T_1906_60,_T_1906_59,_T_1906_58,_T_1906_57,_T_1906_56,_T_2220,_T_2213}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2224.4]
  assign _T_2230 = {_T_2229,_T_2198}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@2225.4]
  assign _T_2231 = _T_2230[0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2226.4]
  assign _T_2296 = _T_2230[1:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2292.4]
  assign _T_2297 = _T_2296[0]; // @[Bitwise.scala 50:65:@2293.4]
  assign _T_2298 = _T_2296[1]; // @[Bitwise.scala 50:65:@2294.4]
  assign _T_2299 = _T_2297 + _T_2298; // @[Bitwise.scala 48:55:@2295.4]
  assign _T_2363 = _T_2230[2:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2360.4]
  assign _T_2364 = _T_2363[0]; // @[Bitwise.scala 50:65:@2361.4]
  assign _T_2365 = _T_2363[1]; // @[Bitwise.scala 50:65:@2362.4]
  assign _T_2366 = _T_2363[2]; // @[Bitwise.scala 50:65:@2363.4]
  assign _T_2367 = _T_2365 + _T_2366; // @[Bitwise.scala 48:55:@2364.4]
  assign _GEN_544 = {{1'd0}, _T_2364}; // @[Bitwise.scala 48:55:@2365.4]
  assign _T_2368 = _GEN_544 + _T_2367; // @[Bitwise.scala 48:55:@2365.4]
  assign _T_2432 = _T_2230[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2430.4]
  assign _T_2433 = _T_2432[0]; // @[Bitwise.scala 50:65:@2431.4]
  assign _T_2434 = _T_2432[1]; // @[Bitwise.scala 50:65:@2432.4]
  assign _T_2435 = _T_2432[2]; // @[Bitwise.scala 50:65:@2433.4]
  assign _T_2436 = _T_2432[3]; // @[Bitwise.scala 50:65:@2434.4]
  assign _T_2437 = _T_2433 + _T_2434; // @[Bitwise.scala 48:55:@2435.4]
  assign _T_2438 = _T_2435 + _T_2436; // @[Bitwise.scala 48:55:@2436.4]
  assign _T_2439 = _T_2437 + _T_2438; // @[Bitwise.scala 48:55:@2437.4]
  assign _T_2503 = _T_2230[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2502.4]
  assign _T_2504 = _T_2503[0]; // @[Bitwise.scala 50:65:@2503.4]
  assign _T_2505 = _T_2503[1]; // @[Bitwise.scala 50:65:@2504.4]
  assign _T_2506 = _T_2503[2]; // @[Bitwise.scala 50:65:@2505.4]
  assign _T_2507 = _T_2503[3]; // @[Bitwise.scala 50:65:@2506.4]
  assign _T_2508 = _T_2503[4]; // @[Bitwise.scala 50:65:@2507.4]
  assign _T_2509 = _T_2504 + _T_2505; // @[Bitwise.scala 48:55:@2508.4]
  assign _T_2510 = _T_2507 + _T_2508; // @[Bitwise.scala 48:55:@2509.4]
  assign _GEN_545 = {{1'd0}, _T_2506}; // @[Bitwise.scala 48:55:@2510.4]
  assign _T_2511 = _GEN_545 + _T_2510; // @[Bitwise.scala 48:55:@2510.4]
  assign _GEN_546 = {{1'd0}, _T_2509}; // @[Bitwise.scala 48:55:@2511.4]
  assign _T_2512 = _GEN_546 + _T_2511; // @[Bitwise.scala 48:55:@2511.4]
  assign _T_2576 = _T_2230[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2576.4]
  assign _T_2577 = _T_2576[0]; // @[Bitwise.scala 50:65:@2577.4]
  assign _T_2578 = _T_2576[1]; // @[Bitwise.scala 50:65:@2578.4]
  assign _T_2579 = _T_2576[2]; // @[Bitwise.scala 50:65:@2579.4]
  assign _T_2580 = _T_2576[3]; // @[Bitwise.scala 50:65:@2580.4]
  assign _T_2581 = _T_2576[4]; // @[Bitwise.scala 50:65:@2581.4]
  assign _T_2582 = _T_2576[5]; // @[Bitwise.scala 50:65:@2582.4]
  assign _T_2583 = _T_2578 + _T_2579; // @[Bitwise.scala 48:55:@2583.4]
  assign _GEN_547 = {{1'd0}, _T_2577}; // @[Bitwise.scala 48:55:@2584.4]
  assign _T_2584 = _GEN_547 + _T_2583; // @[Bitwise.scala 48:55:@2584.4]
  assign _T_2585 = _T_2581 + _T_2582; // @[Bitwise.scala 48:55:@2585.4]
  assign _GEN_548 = {{1'd0}, _T_2580}; // @[Bitwise.scala 48:55:@2586.4]
  assign _T_2586 = _GEN_548 + _T_2585; // @[Bitwise.scala 48:55:@2586.4]
  assign _T_2587 = _T_2584 + _T_2586; // @[Bitwise.scala 48:55:@2587.4]
  assign _T_2651 = _T_2230[6:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2652.4]
  assign _T_2652 = _T_2651[0]; // @[Bitwise.scala 50:65:@2653.4]
  assign _T_2653 = _T_2651[1]; // @[Bitwise.scala 50:65:@2654.4]
  assign _T_2654 = _T_2651[2]; // @[Bitwise.scala 50:65:@2655.4]
  assign _T_2655 = _T_2651[3]; // @[Bitwise.scala 50:65:@2656.4]
  assign _T_2656 = _T_2651[4]; // @[Bitwise.scala 50:65:@2657.4]
  assign _T_2657 = _T_2651[5]; // @[Bitwise.scala 50:65:@2658.4]
  assign _T_2658 = _T_2651[6]; // @[Bitwise.scala 50:65:@2659.4]
  assign _T_2659 = _T_2653 + _T_2654; // @[Bitwise.scala 48:55:@2660.4]
  assign _GEN_549 = {{1'd0}, _T_2652}; // @[Bitwise.scala 48:55:@2661.4]
  assign _T_2660 = _GEN_549 + _T_2659; // @[Bitwise.scala 48:55:@2661.4]
  assign _T_2661 = _T_2655 + _T_2656; // @[Bitwise.scala 48:55:@2662.4]
  assign _T_2662 = _T_2657 + _T_2658; // @[Bitwise.scala 48:55:@2663.4]
  assign _T_2663 = _T_2661 + _T_2662; // @[Bitwise.scala 48:55:@2664.4]
  assign _T_2664 = _T_2660 + _T_2663; // @[Bitwise.scala 48:55:@2665.4]
  assign _T_2728 = _T_2230[7:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2730.4]
  assign _T_2729 = _T_2728[0]; // @[Bitwise.scala 50:65:@2731.4]
  assign _T_2730 = _T_2728[1]; // @[Bitwise.scala 50:65:@2732.4]
  assign _T_2731 = _T_2728[2]; // @[Bitwise.scala 50:65:@2733.4]
  assign _T_2732 = _T_2728[3]; // @[Bitwise.scala 50:65:@2734.4]
  assign _T_2733 = _T_2728[4]; // @[Bitwise.scala 50:65:@2735.4]
  assign _T_2734 = _T_2728[5]; // @[Bitwise.scala 50:65:@2736.4]
  assign _T_2735 = _T_2728[6]; // @[Bitwise.scala 50:65:@2737.4]
  assign _T_2736 = _T_2728[7]; // @[Bitwise.scala 50:65:@2738.4]
  assign _T_2737 = _T_2729 + _T_2730; // @[Bitwise.scala 48:55:@2739.4]
  assign _T_2738 = _T_2731 + _T_2732; // @[Bitwise.scala 48:55:@2740.4]
  assign _T_2739 = _T_2737 + _T_2738; // @[Bitwise.scala 48:55:@2741.4]
  assign _T_2740 = _T_2733 + _T_2734; // @[Bitwise.scala 48:55:@2742.4]
  assign _T_2741 = _T_2735 + _T_2736; // @[Bitwise.scala 48:55:@2743.4]
  assign _T_2742 = _T_2740 + _T_2741; // @[Bitwise.scala 48:55:@2744.4]
  assign _T_2743 = _T_2739 + _T_2742; // @[Bitwise.scala 48:55:@2745.4]
  assign _T_2807 = _T_2230[8:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2810.4]
  assign _T_2808 = _T_2807[0]; // @[Bitwise.scala 50:65:@2811.4]
  assign _T_2809 = _T_2807[1]; // @[Bitwise.scala 50:65:@2812.4]
  assign _T_2810 = _T_2807[2]; // @[Bitwise.scala 50:65:@2813.4]
  assign _T_2811 = _T_2807[3]; // @[Bitwise.scala 50:65:@2814.4]
  assign _T_2812 = _T_2807[4]; // @[Bitwise.scala 50:65:@2815.4]
  assign _T_2813 = _T_2807[5]; // @[Bitwise.scala 50:65:@2816.4]
  assign _T_2814 = _T_2807[6]; // @[Bitwise.scala 50:65:@2817.4]
  assign _T_2815 = _T_2807[7]; // @[Bitwise.scala 50:65:@2818.4]
  assign _T_2816 = _T_2807[8]; // @[Bitwise.scala 50:65:@2819.4]
  assign _T_2817 = _T_2808 + _T_2809; // @[Bitwise.scala 48:55:@2820.4]
  assign _T_2818 = _T_2810 + _T_2811; // @[Bitwise.scala 48:55:@2821.4]
  assign _T_2819 = _T_2817 + _T_2818; // @[Bitwise.scala 48:55:@2822.4]
  assign _T_2820 = _T_2812 + _T_2813; // @[Bitwise.scala 48:55:@2823.4]
  assign _T_2821 = _T_2815 + _T_2816; // @[Bitwise.scala 48:55:@2824.4]
  assign _GEN_550 = {{1'd0}, _T_2814}; // @[Bitwise.scala 48:55:@2825.4]
  assign _T_2822 = _GEN_550 + _T_2821; // @[Bitwise.scala 48:55:@2825.4]
  assign _GEN_551 = {{1'd0}, _T_2820}; // @[Bitwise.scala 48:55:@2826.4]
  assign _T_2823 = _GEN_551 + _T_2822; // @[Bitwise.scala 48:55:@2826.4]
  assign _GEN_552 = {{1'd0}, _T_2819}; // @[Bitwise.scala 48:55:@2827.4]
  assign _T_2824 = _GEN_552 + _T_2823; // @[Bitwise.scala 48:55:@2827.4]
  assign _T_2888 = _T_2230[9:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2892.4]
  assign _T_2889 = _T_2888[0]; // @[Bitwise.scala 50:65:@2893.4]
  assign _T_2890 = _T_2888[1]; // @[Bitwise.scala 50:65:@2894.4]
  assign _T_2891 = _T_2888[2]; // @[Bitwise.scala 50:65:@2895.4]
  assign _T_2892 = _T_2888[3]; // @[Bitwise.scala 50:65:@2896.4]
  assign _T_2893 = _T_2888[4]; // @[Bitwise.scala 50:65:@2897.4]
  assign _T_2894 = _T_2888[5]; // @[Bitwise.scala 50:65:@2898.4]
  assign _T_2895 = _T_2888[6]; // @[Bitwise.scala 50:65:@2899.4]
  assign _T_2896 = _T_2888[7]; // @[Bitwise.scala 50:65:@2900.4]
  assign _T_2897 = _T_2888[8]; // @[Bitwise.scala 50:65:@2901.4]
  assign _T_2898 = _T_2888[9]; // @[Bitwise.scala 50:65:@2902.4]
  assign _T_2899 = _T_2889 + _T_2890; // @[Bitwise.scala 48:55:@2903.4]
  assign _T_2900 = _T_2892 + _T_2893; // @[Bitwise.scala 48:55:@2904.4]
  assign _GEN_553 = {{1'd0}, _T_2891}; // @[Bitwise.scala 48:55:@2905.4]
  assign _T_2901 = _GEN_553 + _T_2900; // @[Bitwise.scala 48:55:@2905.4]
  assign _GEN_554 = {{1'd0}, _T_2899}; // @[Bitwise.scala 48:55:@2906.4]
  assign _T_2902 = _GEN_554 + _T_2901; // @[Bitwise.scala 48:55:@2906.4]
  assign _T_2903 = _T_2894 + _T_2895; // @[Bitwise.scala 48:55:@2907.4]
  assign _T_2904 = _T_2897 + _T_2898; // @[Bitwise.scala 48:55:@2908.4]
  assign _GEN_555 = {{1'd0}, _T_2896}; // @[Bitwise.scala 48:55:@2909.4]
  assign _T_2905 = _GEN_555 + _T_2904; // @[Bitwise.scala 48:55:@2909.4]
  assign _GEN_556 = {{1'd0}, _T_2903}; // @[Bitwise.scala 48:55:@2910.4]
  assign _T_2906 = _GEN_556 + _T_2905; // @[Bitwise.scala 48:55:@2910.4]
  assign _T_2907 = _T_2902 + _T_2906; // @[Bitwise.scala 48:55:@2911.4]
  assign _T_2971 = _T_2230[10:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2976.4]
  assign _T_2972 = _T_2971[0]; // @[Bitwise.scala 50:65:@2977.4]
  assign _T_2973 = _T_2971[1]; // @[Bitwise.scala 50:65:@2978.4]
  assign _T_2974 = _T_2971[2]; // @[Bitwise.scala 50:65:@2979.4]
  assign _T_2975 = _T_2971[3]; // @[Bitwise.scala 50:65:@2980.4]
  assign _T_2976 = _T_2971[4]; // @[Bitwise.scala 50:65:@2981.4]
  assign _T_2977 = _T_2971[5]; // @[Bitwise.scala 50:65:@2982.4]
  assign _T_2978 = _T_2971[6]; // @[Bitwise.scala 50:65:@2983.4]
  assign _T_2979 = _T_2971[7]; // @[Bitwise.scala 50:65:@2984.4]
  assign _T_2980 = _T_2971[8]; // @[Bitwise.scala 50:65:@2985.4]
  assign _T_2981 = _T_2971[9]; // @[Bitwise.scala 50:65:@2986.4]
  assign _T_2982 = _T_2971[10]; // @[Bitwise.scala 50:65:@2987.4]
  assign _T_2983 = _T_2972 + _T_2973; // @[Bitwise.scala 48:55:@2988.4]
  assign _T_2984 = _T_2975 + _T_2976; // @[Bitwise.scala 48:55:@2989.4]
  assign _GEN_557 = {{1'd0}, _T_2974}; // @[Bitwise.scala 48:55:@2990.4]
  assign _T_2985 = _GEN_557 + _T_2984; // @[Bitwise.scala 48:55:@2990.4]
  assign _GEN_558 = {{1'd0}, _T_2983}; // @[Bitwise.scala 48:55:@2991.4]
  assign _T_2986 = _GEN_558 + _T_2985; // @[Bitwise.scala 48:55:@2991.4]
  assign _T_2987 = _T_2978 + _T_2979; // @[Bitwise.scala 48:55:@2992.4]
  assign _GEN_559 = {{1'd0}, _T_2977}; // @[Bitwise.scala 48:55:@2993.4]
  assign _T_2988 = _GEN_559 + _T_2987; // @[Bitwise.scala 48:55:@2993.4]
  assign _T_2989 = _T_2981 + _T_2982; // @[Bitwise.scala 48:55:@2994.4]
  assign _GEN_560 = {{1'd0}, _T_2980}; // @[Bitwise.scala 48:55:@2995.4]
  assign _T_2990 = _GEN_560 + _T_2989; // @[Bitwise.scala 48:55:@2995.4]
  assign _T_2991 = _T_2988 + _T_2990; // @[Bitwise.scala 48:55:@2996.4]
  assign _T_2992 = _T_2986 + _T_2991; // @[Bitwise.scala 48:55:@2997.4]
  assign _T_3056 = _T_2230[11:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3062.4]
  assign _T_3057 = _T_3056[0]; // @[Bitwise.scala 50:65:@3063.4]
  assign _T_3058 = _T_3056[1]; // @[Bitwise.scala 50:65:@3064.4]
  assign _T_3059 = _T_3056[2]; // @[Bitwise.scala 50:65:@3065.4]
  assign _T_3060 = _T_3056[3]; // @[Bitwise.scala 50:65:@3066.4]
  assign _T_3061 = _T_3056[4]; // @[Bitwise.scala 50:65:@3067.4]
  assign _T_3062 = _T_3056[5]; // @[Bitwise.scala 50:65:@3068.4]
  assign _T_3063 = _T_3056[6]; // @[Bitwise.scala 50:65:@3069.4]
  assign _T_3064 = _T_3056[7]; // @[Bitwise.scala 50:65:@3070.4]
  assign _T_3065 = _T_3056[8]; // @[Bitwise.scala 50:65:@3071.4]
  assign _T_3066 = _T_3056[9]; // @[Bitwise.scala 50:65:@3072.4]
  assign _T_3067 = _T_3056[10]; // @[Bitwise.scala 50:65:@3073.4]
  assign _T_3068 = _T_3056[11]; // @[Bitwise.scala 50:65:@3074.4]
  assign _T_3069 = _T_3058 + _T_3059; // @[Bitwise.scala 48:55:@3075.4]
  assign _GEN_561 = {{1'd0}, _T_3057}; // @[Bitwise.scala 48:55:@3076.4]
  assign _T_3070 = _GEN_561 + _T_3069; // @[Bitwise.scala 48:55:@3076.4]
  assign _T_3071 = _T_3061 + _T_3062; // @[Bitwise.scala 48:55:@3077.4]
  assign _GEN_562 = {{1'd0}, _T_3060}; // @[Bitwise.scala 48:55:@3078.4]
  assign _T_3072 = _GEN_562 + _T_3071; // @[Bitwise.scala 48:55:@3078.4]
  assign _T_3073 = _T_3070 + _T_3072; // @[Bitwise.scala 48:55:@3079.4]
  assign _T_3074 = _T_3064 + _T_3065; // @[Bitwise.scala 48:55:@3080.4]
  assign _GEN_563 = {{1'd0}, _T_3063}; // @[Bitwise.scala 48:55:@3081.4]
  assign _T_3075 = _GEN_563 + _T_3074; // @[Bitwise.scala 48:55:@3081.4]
  assign _T_3076 = _T_3067 + _T_3068; // @[Bitwise.scala 48:55:@3082.4]
  assign _GEN_564 = {{1'd0}, _T_3066}; // @[Bitwise.scala 48:55:@3083.4]
  assign _T_3077 = _GEN_564 + _T_3076; // @[Bitwise.scala 48:55:@3083.4]
  assign _T_3078 = _T_3075 + _T_3077; // @[Bitwise.scala 48:55:@3084.4]
  assign _T_3079 = _T_3073 + _T_3078; // @[Bitwise.scala 48:55:@3085.4]
  assign _T_3143 = _T_2230[12:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3150.4]
  assign _T_3144 = _T_3143[0]; // @[Bitwise.scala 50:65:@3151.4]
  assign _T_3145 = _T_3143[1]; // @[Bitwise.scala 50:65:@3152.4]
  assign _T_3146 = _T_3143[2]; // @[Bitwise.scala 50:65:@3153.4]
  assign _T_3147 = _T_3143[3]; // @[Bitwise.scala 50:65:@3154.4]
  assign _T_3148 = _T_3143[4]; // @[Bitwise.scala 50:65:@3155.4]
  assign _T_3149 = _T_3143[5]; // @[Bitwise.scala 50:65:@3156.4]
  assign _T_3150 = _T_3143[6]; // @[Bitwise.scala 50:65:@3157.4]
  assign _T_3151 = _T_3143[7]; // @[Bitwise.scala 50:65:@3158.4]
  assign _T_3152 = _T_3143[8]; // @[Bitwise.scala 50:65:@3159.4]
  assign _T_3153 = _T_3143[9]; // @[Bitwise.scala 50:65:@3160.4]
  assign _T_3154 = _T_3143[10]; // @[Bitwise.scala 50:65:@3161.4]
  assign _T_3155 = _T_3143[11]; // @[Bitwise.scala 50:65:@3162.4]
  assign _T_3156 = _T_3143[12]; // @[Bitwise.scala 50:65:@3163.4]
  assign _T_3157 = _T_3145 + _T_3146; // @[Bitwise.scala 48:55:@3164.4]
  assign _GEN_565 = {{1'd0}, _T_3144}; // @[Bitwise.scala 48:55:@3165.4]
  assign _T_3158 = _GEN_565 + _T_3157; // @[Bitwise.scala 48:55:@3165.4]
  assign _T_3159 = _T_3148 + _T_3149; // @[Bitwise.scala 48:55:@3166.4]
  assign _GEN_566 = {{1'd0}, _T_3147}; // @[Bitwise.scala 48:55:@3167.4]
  assign _T_3160 = _GEN_566 + _T_3159; // @[Bitwise.scala 48:55:@3167.4]
  assign _T_3161 = _T_3158 + _T_3160; // @[Bitwise.scala 48:55:@3168.4]
  assign _T_3162 = _T_3151 + _T_3152; // @[Bitwise.scala 48:55:@3169.4]
  assign _GEN_567 = {{1'd0}, _T_3150}; // @[Bitwise.scala 48:55:@3170.4]
  assign _T_3163 = _GEN_567 + _T_3162; // @[Bitwise.scala 48:55:@3170.4]
  assign _T_3164 = _T_3153 + _T_3154; // @[Bitwise.scala 48:55:@3171.4]
  assign _T_3165 = _T_3155 + _T_3156; // @[Bitwise.scala 48:55:@3172.4]
  assign _T_3166 = _T_3164 + _T_3165; // @[Bitwise.scala 48:55:@3173.4]
  assign _T_3167 = _T_3163 + _T_3166; // @[Bitwise.scala 48:55:@3174.4]
  assign _T_3168 = _T_3161 + _T_3167; // @[Bitwise.scala 48:55:@3175.4]
  assign _T_3232 = _T_2230[13:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3240.4]
  assign _T_3233 = _T_3232[0]; // @[Bitwise.scala 50:65:@3241.4]
  assign _T_3234 = _T_3232[1]; // @[Bitwise.scala 50:65:@3242.4]
  assign _T_3235 = _T_3232[2]; // @[Bitwise.scala 50:65:@3243.4]
  assign _T_3236 = _T_3232[3]; // @[Bitwise.scala 50:65:@3244.4]
  assign _T_3237 = _T_3232[4]; // @[Bitwise.scala 50:65:@3245.4]
  assign _T_3238 = _T_3232[5]; // @[Bitwise.scala 50:65:@3246.4]
  assign _T_3239 = _T_3232[6]; // @[Bitwise.scala 50:65:@3247.4]
  assign _T_3240 = _T_3232[7]; // @[Bitwise.scala 50:65:@3248.4]
  assign _T_3241 = _T_3232[8]; // @[Bitwise.scala 50:65:@3249.4]
  assign _T_3242 = _T_3232[9]; // @[Bitwise.scala 50:65:@3250.4]
  assign _T_3243 = _T_3232[10]; // @[Bitwise.scala 50:65:@3251.4]
  assign _T_3244 = _T_3232[11]; // @[Bitwise.scala 50:65:@3252.4]
  assign _T_3245 = _T_3232[12]; // @[Bitwise.scala 50:65:@3253.4]
  assign _T_3246 = _T_3232[13]; // @[Bitwise.scala 50:65:@3254.4]
  assign _T_3247 = _T_3234 + _T_3235; // @[Bitwise.scala 48:55:@3255.4]
  assign _GEN_568 = {{1'd0}, _T_3233}; // @[Bitwise.scala 48:55:@3256.4]
  assign _T_3248 = _GEN_568 + _T_3247; // @[Bitwise.scala 48:55:@3256.4]
  assign _T_3249 = _T_3236 + _T_3237; // @[Bitwise.scala 48:55:@3257.4]
  assign _T_3250 = _T_3238 + _T_3239; // @[Bitwise.scala 48:55:@3258.4]
  assign _T_3251 = _T_3249 + _T_3250; // @[Bitwise.scala 48:55:@3259.4]
  assign _T_3252 = _T_3248 + _T_3251; // @[Bitwise.scala 48:55:@3260.4]
  assign _T_3253 = _T_3241 + _T_3242; // @[Bitwise.scala 48:55:@3261.4]
  assign _GEN_569 = {{1'd0}, _T_3240}; // @[Bitwise.scala 48:55:@3262.4]
  assign _T_3254 = _GEN_569 + _T_3253; // @[Bitwise.scala 48:55:@3262.4]
  assign _T_3255 = _T_3243 + _T_3244; // @[Bitwise.scala 48:55:@3263.4]
  assign _T_3256 = _T_3245 + _T_3246; // @[Bitwise.scala 48:55:@3264.4]
  assign _T_3257 = _T_3255 + _T_3256; // @[Bitwise.scala 48:55:@3265.4]
  assign _T_3258 = _T_3254 + _T_3257; // @[Bitwise.scala 48:55:@3266.4]
  assign _T_3259 = _T_3252 + _T_3258; // @[Bitwise.scala 48:55:@3267.4]
  assign _T_3323 = _T_2230[14:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3332.4]
  assign _T_3324 = _T_3323[0]; // @[Bitwise.scala 50:65:@3333.4]
  assign _T_3325 = _T_3323[1]; // @[Bitwise.scala 50:65:@3334.4]
  assign _T_3326 = _T_3323[2]; // @[Bitwise.scala 50:65:@3335.4]
  assign _T_3327 = _T_3323[3]; // @[Bitwise.scala 50:65:@3336.4]
  assign _T_3328 = _T_3323[4]; // @[Bitwise.scala 50:65:@3337.4]
  assign _T_3329 = _T_3323[5]; // @[Bitwise.scala 50:65:@3338.4]
  assign _T_3330 = _T_3323[6]; // @[Bitwise.scala 50:65:@3339.4]
  assign _T_3331 = _T_3323[7]; // @[Bitwise.scala 50:65:@3340.4]
  assign _T_3332 = _T_3323[8]; // @[Bitwise.scala 50:65:@3341.4]
  assign _T_3333 = _T_3323[9]; // @[Bitwise.scala 50:65:@3342.4]
  assign _T_3334 = _T_3323[10]; // @[Bitwise.scala 50:65:@3343.4]
  assign _T_3335 = _T_3323[11]; // @[Bitwise.scala 50:65:@3344.4]
  assign _T_3336 = _T_3323[12]; // @[Bitwise.scala 50:65:@3345.4]
  assign _T_3337 = _T_3323[13]; // @[Bitwise.scala 50:65:@3346.4]
  assign _T_3338 = _T_3323[14]; // @[Bitwise.scala 50:65:@3347.4]
  assign _T_3339 = _T_3325 + _T_3326; // @[Bitwise.scala 48:55:@3348.4]
  assign _GEN_570 = {{1'd0}, _T_3324}; // @[Bitwise.scala 48:55:@3349.4]
  assign _T_3340 = _GEN_570 + _T_3339; // @[Bitwise.scala 48:55:@3349.4]
  assign _T_3341 = _T_3327 + _T_3328; // @[Bitwise.scala 48:55:@3350.4]
  assign _T_3342 = _T_3329 + _T_3330; // @[Bitwise.scala 48:55:@3351.4]
  assign _T_3343 = _T_3341 + _T_3342; // @[Bitwise.scala 48:55:@3352.4]
  assign _T_3344 = _T_3340 + _T_3343; // @[Bitwise.scala 48:55:@3353.4]
  assign _T_3345 = _T_3331 + _T_3332; // @[Bitwise.scala 48:55:@3354.4]
  assign _T_3346 = _T_3333 + _T_3334; // @[Bitwise.scala 48:55:@3355.4]
  assign _T_3347 = _T_3345 + _T_3346; // @[Bitwise.scala 48:55:@3356.4]
  assign _T_3348 = _T_3335 + _T_3336; // @[Bitwise.scala 48:55:@3357.4]
  assign _T_3349 = _T_3337 + _T_3338; // @[Bitwise.scala 48:55:@3358.4]
  assign _T_3350 = _T_3348 + _T_3349; // @[Bitwise.scala 48:55:@3359.4]
  assign _T_3351 = _T_3347 + _T_3350; // @[Bitwise.scala 48:55:@3360.4]
  assign _T_3352 = _T_3344 + _T_3351; // @[Bitwise.scala 48:55:@3361.4]
  assign _T_3416 = _T_2230[15:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3426.4]
  assign _T_3417 = _T_3416[0]; // @[Bitwise.scala 50:65:@3427.4]
  assign _T_3418 = _T_3416[1]; // @[Bitwise.scala 50:65:@3428.4]
  assign _T_3419 = _T_3416[2]; // @[Bitwise.scala 50:65:@3429.4]
  assign _T_3420 = _T_3416[3]; // @[Bitwise.scala 50:65:@3430.4]
  assign _T_3421 = _T_3416[4]; // @[Bitwise.scala 50:65:@3431.4]
  assign _T_3422 = _T_3416[5]; // @[Bitwise.scala 50:65:@3432.4]
  assign _T_3423 = _T_3416[6]; // @[Bitwise.scala 50:65:@3433.4]
  assign _T_3424 = _T_3416[7]; // @[Bitwise.scala 50:65:@3434.4]
  assign _T_3425 = _T_3416[8]; // @[Bitwise.scala 50:65:@3435.4]
  assign _T_3426 = _T_3416[9]; // @[Bitwise.scala 50:65:@3436.4]
  assign _T_3427 = _T_3416[10]; // @[Bitwise.scala 50:65:@3437.4]
  assign _T_3428 = _T_3416[11]; // @[Bitwise.scala 50:65:@3438.4]
  assign _T_3429 = _T_3416[12]; // @[Bitwise.scala 50:65:@3439.4]
  assign _T_3430 = _T_3416[13]; // @[Bitwise.scala 50:65:@3440.4]
  assign _T_3431 = _T_3416[14]; // @[Bitwise.scala 50:65:@3441.4]
  assign _T_3432 = _T_3416[15]; // @[Bitwise.scala 50:65:@3442.4]
  assign _T_3433 = _T_3417 + _T_3418; // @[Bitwise.scala 48:55:@3443.4]
  assign _T_3434 = _T_3419 + _T_3420; // @[Bitwise.scala 48:55:@3444.4]
  assign _T_3435 = _T_3433 + _T_3434; // @[Bitwise.scala 48:55:@3445.4]
  assign _T_3436 = _T_3421 + _T_3422; // @[Bitwise.scala 48:55:@3446.4]
  assign _T_3437 = _T_3423 + _T_3424; // @[Bitwise.scala 48:55:@3447.4]
  assign _T_3438 = _T_3436 + _T_3437; // @[Bitwise.scala 48:55:@3448.4]
  assign _T_3439 = _T_3435 + _T_3438; // @[Bitwise.scala 48:55:@3449.4]
  assign _T_3440 = _T_3425 + _T_3426; // @[Bitwise.scala 48:55:@3450.4]
  assign _T_3441 = _T_3427 + _T_3428; // @[Bitwise.scala 48:55:@3451.4]
  assign _T_3442 = _T_3440 + _T_3441; // @[Bitwise.scala 48:55:@3452.4]
  assign _T_3443 = _T_3429 + _T_3430; // @[Bitwise.scala 48:55:@3453.4]
  assign _T_3444 = _T_3431 + _T_3432; // @[Bitwise.scala 48:55:@3454.4]
  assign _T_3445 = _T_3443 + _T_3444; // @[Bitwise.scala 48:55:@3455.4]
  assign _T_3446 = _T_3442 + _T_3445; // @[Bitwise.scala 48:55:@3456.4]
  assign _T_3447 = _T_3439 + _T_3446; // @[Bitwise.scala 48:55:@3457.4]
  assign _T_3511 = _T_2230[16:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3522.4]
  assign _T_3512 = _T_3511[0]; // @[Bitwise.scala 50:65:@3523.4]
  assign _T_3513 = _T_3511[1]; // @[Bitwise.scala 50:65:@3524.4]
  assign _T_3514 = _T_3511[2]; // @[Bitwise.scala 50:65:@3525.4]
  assign _T_3515 = _T_3511[3]; // @[Bitwise.scala 50:65:@3526.4]
  assign _T_3516 = _T_3511[4]; // @[Bitwise.scala 50:65:@3527.4]
  assign _T_3517 = _T_3511[5]; // @[Bitwise.scala 50:65:@3528.4]
  assign _T_3518 = _T_3511[6]; // @[Bitwise.scala 50:65:@3529.4]
  assign _T_3519 = _T_3511[7]; // @[Bitwise.scala 50:65:@3530.4]
  assign _T_3520 = _T_3511[8]; // @[Bitwise.scala 50:65:@3531.4]
  assign _T_3521 = _T_3511[9]; // @[Bitwise.scala 50:65:@3532.4]
  assign _T_3522 = _T_3511[10]; // @[Bitwise.scala 50:65:@3533.4]
  assign _T_3523 = _T_3511[11]; // @[Bitwise.scala 50:65:@3534.4]
  assign _T_3524 = _T_3511[12]; // @[Bitwise.scala 50:65:@3535.4]
  assign _T_3525 = _T_3511[13]; // @[Bitwise.scala 50:65:@3536.4]
  assign _T_3526 = _T_3511[14]; // @[Bitwise.scala 50:65:@3537.4]
  assign _T_3527 = _T_3511[15]; // @[Bitwise.scala 50:65:@3538.4]
  assign _T_3528 = _T_3511[16]; // @[Bitwise.scala 50:65:@3539.4]
  assign _T_3529 = _T_3512 + _T_3513; // @[Bitwise.scala 48:55:@3540.4]
  assign _T_3530 = _T_3514 + _T_3515; // @[Bitwise.scala 48:55:@3541.4]
  assign _T_3531 = _T_3529 + _T_3530; // @[Bitwise.scala 48:55:@3542.4]
  assign _T_3532 = _T_3516 + _T_3517; // @[Bitwise.scala 48:55:@3543.4]
  assign _T_3533 = _T_3518 + _T_3519; // @[Bitwise.scala 48:55:@3544.4]
  assign _T_3534 = _T_3532 + _T_3533; // @[Bitwise.scala 48:55:@3545.4]
  assign _T_3535 = _T_3531 + _T_3534; // @[Bitwise.scala 48:55:@3546.4]
  assign _T_3536 = _T_3520 + _T_3521; // @[Bitwise.scala 48:55:@3547.4]
  assign _T_3537 = _T_3522 + _T_3523; // @[Bitwise.scala 48:55:@3548.4]
  assign _T_3538 = _T_3536 + _T_3537; // @[Bitwise.scala 48:55:@3549.4]
  assign _T_3539 = _T_3524 + _T_3525; // @[Bitwise.scala 48:55:@3550.4]
  assign _T_3540 = _T_3527 + _T_3528; // @[Bitwise.scala 48:55:@3551.4]
  assign _GEN_571 = {{1'd0}, _T_3526}; // @[Bitwise.scala 48:55:@3552.4]
  assign _T_3541 = _GEN_571 + _T_3540; // @[Bitwise.scala 48:55:@3552.4]
  assign _GEN_572 = {{1'd0}, _T_3539}; // @[Bitwise.scala 48:55:@3553.4]
  assign _T_3542 = _GEN_572 + _T_3541; // @[Bitwise.scala 48:55:@3553.4]
  assign _GEN_573 = {{1'd0}, _T_3538}; // @[Bitwise.scala 48:55:@3554.4]
  assign _T_3543 = _GEN_573 + _T_3542; // @[Bitwise.scala 48:55:@3554.4]
  assign _GEN_574 = {{1'd0}, _T_3535}; // @[Bitwise.scala 48:55:@3555.4]
  assign _T_3544 = _GEN_574 + _T_3543; // @[Bitwise.scala 48:55:@3555.4]
  assign _T_3608 = _T_2230[17:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3620.4]
  assign _T_3609 = _T_3608[0]; // @[Bitwise.scala 50:65:@3621.4]
  assign _T_3610 = _T_3608[1]; // @[Bitwise.scala 50:65:@3622.4]
  assign _T_3611 = _T_3608[2]; // @[Bitwise.scala 50:65:@3623.4]
  assign _T_3612 = _T_3608[3]; // @[Bitwise.scala 50:65:@3624.4]
  assign _T_3613 = _T_3608[4]; // @[Bitwise.scala 50:65:@3625.4]
  assign _T_3614 = _T_3608[5]; // @[Bitwise.scala 50:65:@3626.4]
  assign _T_3615 = _T_3608[6]; // @[Bitwise.scala 50:65:@3627.4]
  assign _T_3616 = _T_3608[7]; // @[Bitwise.scala 50:65:@3628.4]
  assign _T_3617 = _T_3608[8]; // @[Bitwise.scala 50:65:@3629.4]
  assign _T_3618 = _T_3608[9]; // @[Bitwise.scala 50:65:@3630.4]
  assign _T_3619 = _T_3608[10]; // @[Bitwise.scala 50:65:@3631.4]
  assign _T_3620 = _T_3608[11]; // @[Bitwise.scala 50:65:@3632.4]
  assign _T_3621 = _T_3608[12]; // @[Bitwise.scala 50:65:@3633.4]
  assign _T_3622 = _T_3608[13]; // @[Bitwise.scala 50:65:@3634.4]
  assign _T_3623 = _T_3608[14]; // @[Bitwise.scala 50:65:@3635.4]
  assign _T_3624 = _T_3608[15]; // @[Bitwise.scala 50:65:@3636.4]
  assign _T_3625 = _T_3608[16]; // @[Bitwise.scala 50:65:@3637.4]
  assign _T_3626 = _T_3608[17]; // @[Bitwise.scala 50:65:@3638.4]
  assign _T_3627 = _T_3609 + _T_3610; // @[Bitwise.scala 48:55:@3639.4]
  assign _T_3628 = _T_3611 + _T_3612; // @[Bitwise.scala 48:55:@3640.4]
  assign _T_3629 = _T_3627 + _T_3628; // @[Bitwise.scala 48:55:@3641.4]
  assign _T_3630 = _T_3613 + _T_3614; // @[Bitwise.scala 48:55:@3642.4]
  assign _T_3631 = _T_3616 + _T_3617; // @[Bitwise.scala 48:55:@3643.4]
  assign _GEN_575 = {{1'd0}, _T_3615}; // @[Bitwise.scala 48:55:@3644.4]
  assign _T_3632 = _GEN_575 + _T_3631; // @[Bitwise.scala 48:55:@3644.4]
  assign _GEN_576 = {{1'd0}, _T_3630}; // @[Bitwise.scala 48:55:@3645.4]
  assign _T_3633 = _GEN_576 + _T_3632; // @[Bitwise.scala 48:55:@3645.4]
  assign _GEN_577 = {{1'd0}, _T_3629}; // @[Bitwise.scala 48:55:@3646.4]
  assign _T_3634 = _GEN_577 + _T_3633; // @[Bitwise.scala 48:55:@3646.4]
  assign _T_3635 = _T_3618 + _T_3619; // @[Bitwise.scala 48:55:@3647.4]
  assign _T_3636 = _T_3620 + _T_3621; // @[Bitwise.scala 48:55:@3648.4]
  assign _T_3637 = _T_3635 + _T_3636; // @[Bitwise.scala 48:55:@3649.4]
  assign _T_3638 = _T_3622 + _T_3623; // @[Bitwise.scala 48:55:@3650.4]
  assign _T_3639 = _T_3625 + _T_3626; // @[Bitwise.scala 48:55:@3651.4]
  assign _GEN_578 = {{1'd0}, _T_3624}; // @[Bitwise.scala 48:55:@3652.4]
  assign _T_3640 = _GEN_578 + _T_3639; // @[Bitwise.scala 48:55:@3652.4]
  assign _GEN_579 = {{1'd0}, _T_3638}; // @[Bitwise.scala 48:55:@3653.4]
  assign _T_3641 = _GEN_579 + _T_3640; // @[Bitwise.scala 48:55:@3653.4]
  assign _GEN_580 = {{1'd0}, _T_3637}; // @[Bitwise.scala 48:55:@3654.4]
  assign _T_3642 = _GEN_580 + _T_3641; // @[Bitwise.scala 48:55:@3654.4]
  assign _T_3643 = _T_3634 + _T_3642; // @[Bitwise.scala 48:55:@3655.4]
  assign _T_3707 = _T_2230[18:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3720.4]
  assign _T_3708 = _T_3707[0]; // @[Bitwise.scala 50:65:@3721.4]
  assign _T_3709 = _T_3707[1]; // @[Bitwise.scala 50:65:@3722.4]
  assign _T_3710 = _T_3707[2]; // @[Bitwise.scala 50:65:@3723.4]
  assign _T_3711 = _T_3707[3]; // @[Bitwise.scala 50:65:@3724.4]
  assign _T_3712 = _T_3707[4]; // @[Bitwise.scala 50:65:@3725.4]
  assign _T_3713 = _T_3707[5]; // @[Bitwise.scala 50:65:@3726.4]
  assign _T_3714 = _T_3707[6]; // @[Bitwise.scala 50:65:@3727.4]
  assign _T_3715 = _T_3707[7]; // @[Bitwise.scala 50:65:@3728.4]
  assign _T_3716 = _T_3707[8]; // @[Bitwise.scala 50:65:@3729.4]
  assign _T_3717 = _T_3707[9]; // @[Bitwise.scala 50:65:@3730.4]
  assign _T_3718 = _T_3707[10]; // @[Bitwise.scala 50:65:@3731.4]
  assign _T_3719 = _T_3707[11]; // @[Bitwise.scala 50:65:@3732.4]
  assign _T_3720 = _T_3707[12]; // @[Bitwise.scala 50:65:@3733.4]
  assign _T_3721 = _T_3707[13]; // @[Bitwise.scala 50:65:@3734.4]
  assign _T_3722 = _T_3707[14]; // @[Bitwise.scala 50:65:@3735.4]
  assign _T_3723 = _T_3707[15]; // @[Bitwise.scala 50:65:@3736.4]
  assign _T_3724 = _T_3707[16]; // @[Bitwise.scala 50:65:@3737.4]
  assign _T_3725 = _T_3707[17]; // @[Bitwise.scala 50:65:@3738.4]
  assign _T_3726 = _T_3707[18]; // @[Bitwise.scala 50:65:@3739.4]
  assign _T_3727 = _T_3708 + _T_3709; // @[Bitwise.scala 48:55:@3740.4]
  assign _T_3728 = _T_3710 + _T_3711; // @[Bitwise.scala 48:55:@3741.4]
  assign _T_3729 = _T_3727 + _T_3728; // @[Bitwise.scala 48:55:@3742.4]
  assign _T_3730 = _T_3712 + _T_3713; // @[Bitwise.scala 48:55:@3743.4]
  assign _T_3731 = _T_3715 + _T_3716; // @[Bitwise.scala 48:55:@3744.4]
  assign _GEN_581 = {{1'd0}, _T_3714}; // @[Bitwise.scala 48:55:@3745.4]
  assign _T_3732 = _GEN_581 + _T_3731; // @[Bitwise.scala 48:55:@3745.4]
  assign _GEN_582 = {{1'd0}, _T_3730}; // @[Bitwise.scala 48:55:@3746.4]
  assign _T_3733 = _GEN_582 + _T_3732; // @[Bitwise.scala 48:55:@3746.4]
  assign _GEN_583 = {{1'd0}, _T_3729}; // @[Bitwise.scala 48:55:@3747.4]
  assign _T_3734 = _GEN_583 + _T_3733; // @[Bitwise.scala 48:55:@3747.4]
  assign _T_3735 = _T_3717 + _T_3718; // @[Bitwise.scala 48:55:@3748.4]
  assign _T_3736 = _T_3720 + _T_3721; // @[Bitwise.scala 48:55:@3749.4]
  assign _GEN_584 = {{1'd0}, _T_3719}; // @[Bitwise.scala 48:55:@3750.4]
  assign _T_3737 = _GEN_584 + _T_3736; // @[Bitwise.scala 48:55:@3750.4]
  assign _GEN_585 = {{1'd0}, _T_3735}; // @[Bitwise.scala 48:55:@3751.4]
  assign _T_3738 = _GEN_585 + _T_3737; // @[Bitwise.scala 48:55:@3751.4]
  assign _T_3739 = _T_3722 + _T_3723; // @[Bitwise.scala 48:55:@3752.4]
  assign _T_3740 = _T_3725 + _T_3726; // @[Bitwise.scala 48:55:@3753.4]
  assign _GEN_586 = {{1'd0}, _T_3724}; // @[Bitwise.scala 48:55:@3754.4]
  assign _T_3741 = _GEN_586 + _T_3740; // @[Bitwise.scala 48:55:@3754.4]
  assign _GEN_587 = {{1'd0}, _T_3739}; // @[Bitwise.scala 48:55:@3755.4]
  assign _T_3742 = _GEN_587 + _T_3741; // @[Bitwise.scala 48:55:@3755.4]
  assign _T_3743 = _T_3738 + _T_3742; // @[Bitwise.scala 48:55:@3756.4]
  assign _T_3744 = _T_3734 + _T_3743; // @[Bitwise.scala 48:55:@3757.4]
  assign _T_3808 = _T_2230[19:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3822.4]
  assign _T_3809 = _T_3808[0]; // @[Bitwise.scala 50:65:@3823.4]
  assign _T_3810 = _T_3808[1]; // @[Bitwise.scala 50:65:@3824.4]
  assign _T_3811 = _T_3808[2]; // @[Bitwise.scala 50:65:@3825.4]
  assign _T_3812 = _T_3808[3]; // @[Bitwise.scala 50:65:@3826.4]
  assign _T_3813 = _T_3808[4]; // @[Bitwise.scala 50:65:@3827.4]
  assign _T_3814 = _T_3808[5]; // @[Bitwise.scala 50:65:@3828.4]
  assign _T_3815 = _T_3808[6]; // @[Bitwise.scala 50:65:@3829.4]
  assign _T_3816 = _T_3808[7]; // @[Bitwise.scala 50:65:@3830.4]
  assign _T_3817 = _T_3808[8]; // @[Bitwise.scala 50:65:@3831.4]
  assign _T_3818 = _T_3808[9]; // @[Bitwise.scala 50:65:@3832.4]
  assign _T_3819 = _T_3808[10]; // @[Bitwise.scala 50:65:@3833.4]
  assign _T_3820 = _T_3808[11]; // @[Bitwise.scala 50:65:@3834.4]
  assign _T_3821 = _T_3808[12]; // @[Bitwise.scala 50:65:@3835.4]
  assign _T_3822 = _T_3808[13]; // @[Bitwise.scala 50:65:@3836.4]
  assign _T_3823 = _T_3808[14]; // @[Bitwise.scala 50:65:@3837.4]
  assign _T_3824 = _T_3808[15]; // @[Bitwise.scala 50:65:@3838.4]
  assign _T_3825 = _T_3808[16]; // @[Bitwise.scala 50:65:@3839.4]
  assign _T_3826 = _T_3808[17]; // @[Bitwise.scala 50:65:@3840.4]
  assign _T_3827 = _T_3808[18]; // @[Bitwise.scala 50:65:@3841.4]
  assign _T_3828 = _T_3808[19]; // @[Bitwise.scala 50:65:@3842.4]
  assign _T_3829 = _T_3809 + _T_3810; // @[Bitwise.scala 48:55:@3843.4]
  assign _T_3830 = _T_3812 + _T_3813; // @[Bitwise.scala 48:55:@3844.4]
  assign _GEN_588 = {{1'd0}, _T_3811}; // @[Bitwise.scala 48:55:@3845.4]
  assign _T_3831 = _GEN_588 + _T_3830; // @[Bitwise.scala 48:55:@3845.4]
  assign _GEN_589 = {{1'd0}, _T_3829}; // @[Bitwise.scala 48:55:@3846.4]
  assign _T_3832 = _GEN_589 + _T_3831; // @[Bitwise.scala 48:55:@3846.4]
  assign _T_3833 = _T_3814 + _T_3815; // @[Bitwise.scala 48:55:@3847.4]
  assign _T_3834 = _T_3817 + _T_3818; // @[Bitwise.scala 48:55:@3848.4]
  assign _GEN_590 = {{1'd0}, _T_3816}; // @[Bitwise.scala 48:55:@3849.4]
  assign _T_3835 = _GEN_590 + _T_3834; // @[Bitwise.scala 48:55:@3849.4]
  assign _GEN_591 = {{1'd0}, _T_3833}; // @[Bitwise.scala 48:55:@3850.4]
  assign _T_3836 = _GEN_591 + _T_3835; // @[Bitwise.scala 48:55:@3850.4]
  assign _T_3837 = _T_3832 + _T_3836; // @[Bitwise.scala 48:55:@3851.4]
  assign _T_3838 = _T_3819 + _T_3820; // @[Bitwise.scala 48:55:@3852.4]
  assign _T_3839 = _T_3822 + _T_3823; // @[Bitwise.scala 48:55:@3853.4]
  assign _GEN_592 = {{1'd0}, _T_3821}; // @[Bitwise.scala 48:55:@3854.4]
  assign _T_3840 = _GEN_592 + _T_3839; // @[Bitwise.scala 48:55:@3854.4]
  assign _GEN_593 = {{1'd0}, _T_3838}; // @[Bitwise.scala 48:55:@3855.4]
  assign _T_3841 = _GEN_593 + _T_3840; // @[Bitwise.scala 48:55:@3855.4]
  assign _T_3842 = _T_3824 + _T_3825; // @[Bitwise.scala 48:55:@3856.4]
  assign _T_3843 = _T_3827 + _T_3828; // @[Bitwise.scala 48:55:@3857.4]
  assign _GEN_594 = {{1'd0}, _T_3826}; // @[Bitwise.scala 48:55:@3858.4]
  assign _T_3844 = _GEN_594 + _T_3843; // @[Bitwise.scala 48:55:@3858.4]
  assign _GEN_595 = {{1'd0}, _T_3842}; // @[Bitwise.scala 48:55:@3859.4]
  assign _T_3845 = _GEN_595 + _T_3844; // @[Bitwise.scala 48:55:@3859.4]
  assign _T_3846 = _T_3841 + _T_3845; // @[Bitwise.scala 48:55:@3860.4]
  assign _T_3847 = _T_3837 + _T_3846; // @[Bitwise.scala 48:55:@3861.4]
  assign _T_3911 = _T_2230[20:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3926.4]
  assign _T_3912 = _T_3911[0]; // @[Bitwise.scala 50:65:@3927.4]
  assign _T_3913 = _T_3911[1]; // @[Bitwise.scala 50:65:@3928.4]
  assign _T_3914 = _T_3911[2]; // @[Bitwise.scala 50:65:@3929.4]
  assign _T_3915 = _T_3911[3]; // @[Bitwise.scala 50:65:@3930.4]
  assign _T_3916 = _T_3911[4]; // @[Bitwise.scala 50:65:@3931.4]
  assign _T_3917 = _T_3911[5]; // @[Bitwise.scala 50:65:@3932.4]
  assign _T_3918 = _T_3911[6]; // @[Bitwise.scala 50:65:@3933.4]
  assign _T_3919 = _T_3911[7]; // @[Bitwise.scala 50:65:@3934.4]
  assign _T_3920 = _T_3911[8]; // @[Bitwise.scala 50:65:@3935.4]
  assign _T_3921 = _T_3911[9]; // @[Bitwise.scala 50:65:@3936.4]
  assign _T_3922 = _T_3911[10]; // @[Bitwise.scala 50:65:@3937.4]
  assign _T_3923 = _T_3911[11]; // @[Bitwise.scala 50:65:@3938.4]
  assign _T_3924 = _T_3911[12]; // @[Bitwise.scala 50:65:@3939.4]
  assign _T_3925 = _T_3911[13]; // @[Bitwise.scala 50:65:@3940.4]
  assign _T_3926 = _T_3911[14]; // @[Bitwise.scala 50:65:@3941.4]
  assign _T_3927 = _T_3911[15]; // @[Bitwise.scala 50:65:@3942.4]
  assign _T_3928 = _T_3911[16]; // @[Bitwise.scala 50:65:@3943.4]
  assign _T_3929 = _T_3911[17]; // @[Bitwise.scala 50:65:@3944.4]
  assign _T_3930 = _T_3911[18]; // @[Bitwise.scala 50:65:@3945.4]
  assign _T_3931 = _T_3911[19]; // @[Bitwise.scala 50:65:@3946.4]
  assign _T_3932 = _T_3911[20]; // @[Bitwise.scala 50:65:@3947.4]
  assign _T_3933 = _T_3912 + _T_3913; // @[Bitwise.scala 48:55:@3948.4]
  assign _T_3934 = _T_3915 + _T_3916; // @[Bitwise.scala 48:55:@3949.4]
  assign _GEN_596 = {{1'd0}, _T_3914}; // @[Bitwise.scala 48:55:@3950.4]
  assign _T_3935 = _GEN_596 + _T_3934; // @[Bitwise.scala 48:55:@3950.4]
  assign _GEN_597 = {{1'd0}, _T_3933}; // @[Bitwise.scala 48:55:@3951.4]
  assign _T_3936 = _GEN_597 + _T_3935; // @[Bitwise.scala 48:55:@3951.4]
  assign _T_3937 = _T_3917 + _T_3918; // @[Bitwise.scala 48:55:@3952.4]
  assign _T_3938 = _T_3920 + _T_3921; // @[Bitwise.scala 48:55:@3953.4]
  assign _GEN_598 = {{1'd0}, _T_3919}; // @[Bitwise.scala 48:55:@3954.4]
  assign _T_3939 = _GEN_598 + _T_3938; // @[Bitwise.scala 48:55:@3954.4]
  assign _GEN_599 = {{1'd0}, _T_3937}; // @[Bitwise.scala 48:55:@3955.4]
  assign _T_3940 = _GEN_599 + _T_3939; // @[Bitwise.scala 48:55:@3955.4]
  assign _T_3941 = _T_3936 + _T_3940; // @[Bitwise.scala 48:55:@3956.4]
  assign _T_3942 = _T_3922 + _T_3923; // @[Bitwise.scala 48:55:@3957.4]
  assign _T_3943 = _T_3925 + _T_3926; // @[Bitwise.scala 48:55:@3958.4]
  assign _GEN_600 = {{1'd0}, _T_3924}; // @[Bitwise.scala 48:55:@3959.4]
  assign _T_3944 = _GEN_600 + _T_3943; // @[Bitwise.scala 48:55:@3959.4]
  assign _GEN_601 = {{1'd0}, _T_3942}; // @[Bitwise.scala 48:55:@3960.4]
  assign _T_3945 = _GEN_601 + _T_3944; // @[Bitwise.scala 48:55:@3960.4]
  assign _T_3946 = _T_3928 + _T_3929; // @[Bitwise.scala 48:55:@3961.4]
  assign _GEN_602 = {{1'd0}, _T_3927}; // @[Bitwise.scala 48:55:@3962.4]
  assign _T_3947 = _GEN_602 + _T_3946; // @[Bitwise.scala 48:55:@3962.4]
  assign _T_3948 = _T_3931 + _T_3932; // @[Bitwise.scala 48:55:@3963.4]
  assign _GEN_603 = {{1'd0}, _T_3930}; // @[Bitwise.scala 48:55:@3964.4]
  assign _T_3949 = _GEN_603 + _T_3948; // @[Bitwise.scala 48:55:@3964.4]
  assign _T_3950 = _T_3947 + _T_3949; // @[Bitwise.scala 48:55:@3965.4]
  assign _T_3951 = _T_3945 + _T_3950; // @[Bitwise.scala 48:55:@3966.4]
  assign _T_3952 = _T_3941 + _T_3951; // @[Bitwise.scala 48:55:@3967.4]
  assign _T_4016 = _T_2230[21:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4032.4]
  assign _T_4017 = _T_4016[0]; // @[Bitwise.scala 50:65:@4033.4]
  assign _T_4018 = _T_4016[1]; // @[Bitwise.scala 50:65:@4034.4]
  assign _T_4019 = _T_4016[2]; // @[Bitwise.scala 50:65:@4035.4]
  assign _T_4020 = _T_4016[3]; // @[Bitwise.scala 50:65:@4036.4]
  assign _T_4021 = _T_4016[4]; // @[Bitwise.scala 50:65:@4037.4]
  assign _T_4022 = _T_4016[5]; // @[Bitwise.scala 50:65:@4038.4]
  assign _T_4023 = _T_4016[6]; // @[Bitwise.scala 50:65:@4039.4]
  assign _T_4024 = _T_4016[7]; // @[Bitwise.scala 50:65:@4040.4]
  assign _T_4025 = _T_4016[8]; // @[Bitwise.scala 50:65:@4041.4]
  assign _T_4026 = _T_4016[9]; // @[Bitwise.scala 50:65:@4042.4]
  assign _T_4027 = _T_4016[10]; // @[Bitwise.scala 50:65:@4043.4]
  assign _T_4028 = _T_4016[11]; // @[Bitwise.scala 50:65:@4044.4]
  assign _T_4029 = _T_4016[12]; // @[Bitwise.scala 50:65:@4045.4]
  assign _T_4030 = _T_4016[13]; // @[Bitwise.scala 50:65:@4046.4]
  assign _T_4031 = _T_4016[14]; // @[Bitwise.scala 50:65:@4047.4]
  assign _T_4032 = _T_4016[15]; // @[Bitwise.scala 50:65:@4048.4]
  assign _T_4033 = _T_4016[16]; // @[Bitwise.scala 50:65:@4049.4]
  assign _T_4034 = _T_4016[17]; // @[Bitwise.scala 50:65:@4050.4]
  assign _T_4035 = _T_4016[18]; // @[Bitwise.scala 50:65:@4051.4]
  assign _T_4036 = _T_4016[19]; // @[Bitwise.scala 50:65:@4052.4]
  assign _T_4037 = _T_4016[20]; // @[Bitwise.scala 50:65:@4053.4]
  assign _T_4038 = _T_4016[21]; // @[Bitwise.scala 50:65:@4054.4]
  assign _T_4039 = _T_4017 + _T_4018; // @[Bitwise.scala 48:55:@4055.4]
  assign _T_4040 = _T_4020 + _T_4021; // @[Bitwise.scala 48:55:@4056.4]
  assign _GEN_604 = {{1'd0}, _T_4019}; // @[Bitwise.scala 48:55:@4057.4]
  assign _T_4041 = _GEN_604 + _T_4040; // @[Bitwise.scala 48:55:@4057.4]
  assign _GEN_605 = {{1'd0}, _T_4039}; // @[Bitwise.scala 48:55:@4058.4]
  assign _T_4042 = _GEN_605 + _T_4041; // @[Bitwise.scala 48:55:@4058.4]
  assign _T_4043 = _T_4023 + _T_4024; // @[Bitwise.scala 48:55:@4059.4]
  assign _GEN_606 = {{1'd0}, _T_4022}; // @[Bitwise.scala 48:55:@4060.4]
  assign _T_4044 = _GEN_606 + _T_4043; // @[Bitwise.scala 48:55:@4060.4]
  assign _T_4045 = _T_4026 + _T_4027; // @[Bitwise.scala 48:55:@4061.4]
  assign _GEN_607 = {{1'd0}, _T_4025}; // @[Bitwise.scala 48:55:@4062.4]
  assign _T_4046 = _GEN_607 + _T_4045; // @[Bitwise.scala 48:55:@4062.4]
  assign _T_4047 = _T_4044 + _T_4046; // @[Bitwise.scala 48:55:@4063.4]
  assign _T_4048 = _T_4042 + _T_4047; // @[Bitwise.scala 48:55:@4064.4]
  assign _T_4049 = _T_4028 + _T_4029; // @[Bitwise.scala 48:55:@4065.4]
  assign _T_4050 = _T_4031 + _T_4032; // @[Bitwise.scala 48:55:@4066.4]
  assign _GEN_608 = {{1'd0}, _T_4030}; // @[Bitwise.scala 48:55:@4067.4]
  assign _T_4051 = _GEN_608 + _T_4050; // @[Bitwise.scala 48:55:@4067.4]
  assign _GEN_609 = {{1'd0}, _T_4049}; // @[Bitwise.scala 48:55:@4068.4]
  assign _T_4052 = _GEN_609 + _T_4051; // @[Bitwise.scala 48:55:@4068.4]
  assign _T_4053 = _T_4034 + _T_4035; // @[Bitwise.scala 48:55:@4069.4]
  assign _GEN_610 = {{1'd0}, _T_4033}; // @[Bitwise.scala 48:55:@4070.4]
  assign _T_4054 = _GEN_610 + _T_4053; // @[Bitwise.scala 48:55:@4070.4]
  assign _T_4055 = _T_4037 + _T_4038; // @[Bitwise.scala 48:55:@4071.4]
  assign _GEN_611 = {{1'd0}, _T_4036}; // @[Bitwise.scala 48:55:@4072.4]
  assign _T_4056 = _GEN_611 + _T_4055; // @[Bitwise.scala 48:55:@4072.4]
  assign _T_4057 = _T_4054 + _T_4056; // @[Bitwise.scala 48:55:@4073.4]
  assign _T_4058 = _T_4052 + _T_4057; // @[Bitwise.scala 48:55:@4074.4]
  assign _T_4059 = _T_4048 + _T_4058; // @[Bitwise.scala 48:55:@4075.4]
  assign _T_4123 = _T_2230[22:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4140.4]
  assign _T_4124 = _T_4123[0]; // @[Bitwise.scala 50:65:@4141.4]
  assign _T_4125 = _T_4123[1]; // @[Bitwise.scala 50:65:@4142.4]
  assign _T_4126 = _T_4123[2]; // @[Bitwise.scala 50:65:@4143.4]
  assign _T_4127 = _T_4123[3]; // @[Bitwise.scala 50:65:@4144.4]
  assign _T_4128 = _T_4123[4]; // @[Bitwise.scala 50:65:@4145.4]
  assign _T_4129 = _T_4123[5]; // @[Bitwise.scala 50:65:@4146.4]
  assign _T_4130 = _T_4123[6]; // @[Bitwise.scala 50:65:@4147.4]
  assign _T_4131 = _T_4123[7]; // @[Bitwise.scala 50:65:@4148.4]
  assign _T_4132 = _T_4123[8]; // @[Bitwise.scala 50:65:@4149.4]
  assign _T_4133 = _T_4123[9]; // @[Bitwise.scala 50:65:@4150.4]
  assign _T_4134 = _T_4123[10]; // @[Bitwise.scala 50:65:@4151.4]
  assign _T_4135 = _T_4123[11]; // @[Bitwise.scala 50:65:@4152.4]
  assign _T_4136 = _T_4123[12]; // @[Bitwise.scala 50:65:@4153.4]
  assign _T_4137 = _T_4123[13]; // @[Bitwise.scala 50:65:@4154.4]
  assign _T_4138 = _T_4123[14]; // @[Bitwise.scala 50:65:@4155.4]
  assign _T_4139 = _T_4123[15]; // @[Bitwise.scala 50:65:@4156.4]
  assign _T_4140 = _T_4123[16]; // @[Bitwise.scala 50:65:@4157.4]
  assign _T_4141 = _T_4123[17]; // @[Bitwise.scala 50:65:@4158.4]
  assign _T_4142 = _T_4123[18]; // @[Bitwise.scala 50:65:@4159.4]
  assign _T_4143 = _T_4123[19]; // @[Bitwise.scala 50:65:@4160.4]
  assign _T_4144 = _T_4123[20]; // @[Bitwise.scala 50:65:@4161.4]
  assign _T_4145 = _T_4123[21]; // @[Bitwise.scala 50:65:@4162.4]
  assign _T_4146 = _T_4123[22]; // @[Bitwise.scala 50:65:@4163.4]
  assign _T_4147 = _T_4124 + _T_4125; // @[Bitwise.scala 48:55:@4164.4]
  assign _T_4148 = _T_4127 + _T_4128; // @[Bitwise.scala 48:55:@4165.4]
  assign _GEN_612 = {{1'd0}, _T_4126}; // @[Bitwise.scala 48:55:@4166.4]
  assign _T_4149 = _GEN_612 + _T_4148; // @[Bitwise.scala 48:55:@4166.4]
  assign _GEN_613 = {{1'd0}, _T_4147}; // @[Bitwise.scala 48:55:@4167.4]
  assign _T_4150 = _GEN_613 + _T_4149; // @[Bitwise.scala 48:55:@4167.4]
  assign _T_4151 = _T_4130 + _T_4131; // @[Bitwise.scala 48:55:@4168.4]
  assign _GEN_614 = {{1'd0}, _T_4129}; // @[Bitwise.scala 48:55:@4169.4]
  assign _T_4152 = _GEN_614 + _T_4151; // @[Bitwise.scala 48:55:@4169.4]
  assign _T_4153 = _T_4133 + _T_4134; // @[Bitwise.scala 48:55:@4170.4]
  assign _GEN_615 = {{1'd0}, _T_4132}; // @[Bitwise.scala 48:55:@4171.4]
  assign _T_4154 = _GEN_615 + _T_4153; // @[Bitwise.scala 48:55:@4171.4]
  assign _T_4155 = _T_4152 + _T_4154; // @[Bitwise.scala 48:55:@4172.4]
  assign _T_4156 = _T_4150 + _T_4155; // @[Bitwise.scala 48:55:@4173.4]
  assign _T_4157 = _T_4136 + _T_4137; // @[Bitwise.scala 48:55:@4174.4]
  assign _GEN_616 = {{1'd0}, _T_4135}; // @[Bitwise.scala 48:55:@4175.4]
  assign _T_4158 = _GEN_616 + _T_4157; // @[Bitwise.scala 48:55:@4175.4]
  assign _T_4159 = _T_4139 + _T_4140; // @[Bitwise.scala 48:55:@4176.4]
  assign _GEN_617 = {{1'd0}, _T_4138}; // @[Bitwise.scala 48:55:@4177.4]
  assign _T_4160 = _GEN_617 + _T_4159; // @[Bitwise.scala 48:55:@4177.4]
  assign _T_4161 = _T_4158 + _T_4160; // @[Bitwise.scala 48:55:@4178.4]
  assign _T_4162 = _T_4142 + _T_4143; // @[Bitwise.scala 48:55:@4179.4]
  assign _GEN_618 = {{1'd0}, _T_4141}; // @[Bitwise.scala 48:55:@4180.4]
  assign _T_4163 = _GEN_618 + _T_4162; // @[Bitwise.scala 48:55:@4180.4]
  assign _T_4164 = _T_4145 + _T_4146; // @[Bitwise.scala 48:55:@4181.4]
  assign _GEN_619 = {{1'd0}, _T_4144}; // @[Bitwise.scala 48:55:@4182.4]
  assign _T_4165 = _GEN_619 + _T_4164; // @[Bitwise.scala 48:55:@4182.4]
  assign _T_4166 = _T_4163 + _T_4165; // @[Bitwise.scala 48:55:@4183.4]
  assign _T_4167 = _T_4161 + _T_4166; // @[Bitwise.scala 48:55:@4184.4]
  assign _T_4168 = _T_4156 + _T_4167; // @[Bitwise.scala 48:55:@4185.4]
  assign _T_4232 = _T_2230[23:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4250.4]
  assign _T_4233 = _T_4232[0]; // @[Bitwise.scala 50:65:@4251.4]
  assign _T_4234 = _T_4232[1]; // @[Bitwise.scala 50:65:@4252.4]
  assign _T_4235 = _T_4232[2]; // @[Bitwise.scala 50:65:@4253.4]
  assign _T_4236 = _T_4232[3]; // @[Bitwise.scala 50:65:@4254.4]
  assign _T_4237 = _T_4232[4]; // @[Bitwise.scala 50:65:@4255.4]
  assign _T_4238 = _T_4232[5]; // @[Bitwise.scala 50:65:@4256.4]
  assign _T_4239 = _T_4232[6]; // @[Bitwise.scala 50:65:@4257.4]
  assign _T_4240 = _T_4232[7]; // @[Bitwise.scala 50:65:@4258.4]
  assign _T_4241 = _T_4232[8]; // @[Bitwise.scala 50:65:@4259.4]
  assign _T_4242 = _T_4232[9]; // @[Bitwise.scala 50:65:@4260.4]
  assign _T_4243 = _T_4232[10]; // @[Bitwise.scala 50:65:@4261.4]
  assign _T_4244 = _T_4232[11]; // @[Bitwise.scala 50:65:@4262.4]
  assign _T_4245 = _T_4232[12]; // @[Bitwise.scala 50:65:@4263.4]
  assign _T_4246 = _T_4232[13]; // @[Bitwise.scala 50:65:@4264.4]
  assign _T_4247 = _T_4232[14]; // @[Bitwise.scala 50:65:@4265.4]
  assign _T_4248 = _T_4232[15]; // @[Bitwise.scala 50:65:@4266.4]
  assign _T_4249 = _T_4232[16]; // @[Bitwise.scala 50:65:@4267.4]
  assign _T_4250 = _T_4232[17]; // @[Bitwise.scala 50:65:@4268.4]
  assign _T_4251 = _T_4232[18]; // @[Bitwise.scala 50:65:@4269.4]
  assign _T_4252 = _T_4232[19]; // @[Bitwise.scala 50:65:@4270.4]
  assign _T_4253 = _T_4232[20]; // @[Bitwise.scala 50:65:@4271.4]
  assign _T_4254 = _T_4232[21]; // @[Bitwise.scala 50:65:@4272.4]
  assign _T_4255 = _T_4232[22]; // @[Bitwise.scala 50:65:@4273.4]
  assign _T_4256 = _T_4232[23]; // @[Bitwise.scala 50:65:@4274.4]
  assign _T_4257 = _T_4234 + _T_4235; // @[Bitwise.scala 48:55:@4275.4]
  assign _GEN_620 = {{1'd0}, _T_4233}; // @[Bitwise.scala 48:55:@4276.4]
  assign _T_4258 = _GEN_620 + _T_4257; // @[Bitwise.scala 48:55:@4276.4]
  assign _T_4259 = _T_4237 + _T_4238; // @[Bitwise.scala 48:55:@4277.4]
  assign _GEN_621 = {{1'd0}, _T_4236}; // @[Bitwise.scala 48:55:@4278.4]
  assign _T_4260 = _GEN_621 + _T_4259; // @[Bitwise.scala 48:55:@4278.4]
  assign _T_4261 = _T_4258 + _T_4260; // @[Bitwise.scala 48:55:@4279.4]
  assign _T_4262 = _T_4240 + _T_4241; // @[Bitwise.scala 48:55:@4280.4]
  assign _GEN_622 = {{1'd0}, _T_4239}; // @[Bitwise.scala 48:55:@4281.4]
  assign _T_4263 = _GEN_622 + _T_4262; // @[Bitwise.scala 48:55:@4281.4]
  assign _T_4264 = _T_4243 + _T_4244; // @[Bitwise.scala 48:55:@4282.4]
  assign _GEN_623 = {{1'd0}, _T_4242}; // @[Bitwise.scala 48:55:@4283.4]
  assign _T_4265 = _GEN_623 + _T_4264; // @[Bitwise.scala 48:55:@4283.4]
  assign _T_4266 = _T_4263 + _T_4265; // @[Bitwise.scala 48:55:@4284.4]
  assign _T_4267 = _T_4261 + _T_4266; // @[Bitwise.scala 48:55:@4285.4]
  assign _T_4268 = _T_4246 + _T_4247; // @[Bitwise.scala 48:55:@4286.4]
  assign _GEN_624 = {{1'd0}, _T_4245}; // @[Bitwise.scala 48:55:@4287.4]
  assign _T_4269 = _GEN_624 + _T_4268; // @[Bitwise.scala 48:55:@4287.4]
  assign _T_4270 = _T_4249 + _T_4250; // @[Bitwise.scala 48:55:@4288.4]
  assign _GEN_625 = {{1'd0}, _T_4248}; // @[Bitwise.scala 48:55:@4289.4]
  assign _T_4271 = _GEN_625 + _T_4270; // @[Bitwise.scala 48:55:@4289.4]
  assign _T_4272 = _T_4269 + _T_4271; // @[Bitwise.scala 48:55:@4290.4]
  assign _T_4273 = _T_4252 + _T_4253; // @[Bitwise.scala 48:55:@4291.4]
  assign _GEN_626 = {{1'd0}, _T_4251}; // @[Bitwise.scala 48:55:@4292.4]
  assign _T_4274 = _GEN_626 + _T_4273; // @[Bitwise.scala 48:55:@4292.4]
  assign _T_4275 = _T_4255 + _T_4256; // @[Bitwise.scala 48:55:@4293.4]
  assign _GEN_627 = {{1'd0}, _T_4254}; // @[Bitwise.scala 48:55:@4294.4]
  assign _T_4276 = _GEN_627 + _T_4275; // @[Bitwise.scala 48:55:@4294.4]
  assign _T_4277 = _T_4274 + _T_4276; // @[Bitwise.scala 48:55:@4295.4]
  assign _T_4278 = _T_4272 + _T_4277; // @[Bitwise.scala 48:55:@4296.4]
  assign _T_4279 = _T_4267 + _T_4278; // @[Bitwise.scala 48:55:@4297.4]
  assign _T_4343 = _T_2230[24:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4362.4]
  assign _T_4344 = _T_4343[0]; // @[Bitwise.scala 50:65:@4363.4]
  assign _T_4345 = _T_4343[1]; // @[Bitwise.scala 50:65:@4364.4]
  assign _T_4346 = _T_4343[2]; // @[Bitwise.scala 50:65:@4365.4]
  assign _T_4347 = _T_4343[3]; // @[Bitwise.scala 50:65:@4366.4]
  assign _T_4348 = _T_4343[4]; // @[Bitwise.scala 50:65:@4367.4]
  assign _T_4349 = _T_4343[5]; // @[Bitwise.scala 50:65:@4368.4]
  assign _T_4350 = _T_4343[6]; // @[Bitwise.scala 50:65:@4369.4]
  assign _T_4351 = _T_4343[7]; // @[Bitwise.scala 50:65:@4370.4]
  assign _T_4352 = _T_4343[8]; // @[Bitwise.scala 50:65:@4371.4]
  assign _T_4353 = _T_4343[9]; // @[Bitwise.scala 50:65:@4372.4]
  assign _T_4354 = _T_4343[10]; // @[Bitwise.scala 50:65:@4373.4]
  assign _T_4355 = _T_4343[11]; // @[Bitwise.scala 50:65:@4374.4]
  assign _T_4356 = _T_4343[12]; // @[Bitwise.scala 50:65:@4375.4]
  assign _T_4357 = _T_4343[13]; // @[Bitwise.scala 50:65:@4376.4]
  assign _T_4358 = _T_4343[14]; // @[Bitwise.scala 50:65:@4377.4]
  assign _T_4359 = _T_4343[15]; // @[Bitwise.scala 50:65:@4378.4]
  assign _T_4360 = _T_4343[16]; // @[Bitwise.scala 50:65:@4379.4]
  assign _T_4361 = _T_4343[17]; // @[Bitwise.scala 50:65:@4380.4]
  assign _T_4362 = _T_4343[18]; // @[Bitwise.scala 50:65:@4381.4]
  assign _T_4363 = _T_4343[19]; // @[Bitwise.scala 50:65:@4382.4]
  assign _T_4364 = _T_4343[20]; // @[Bitwise.scala 50:65:@4383.4]
  assign _T_4365 = _T_4343[21]; // @[Bitwise.scala 50:65:@4384.4]
  assign _T_4366 = _T_4343[22]; // @[Bitwise.scala 50:65:@4385.4]
  assign _T_4367 = _T_4343[23]; // @[Bitwise.scala 50:65:@4386.4]
  assign _T_4368 = _T_4343[24]; // @[Bitwise.scala 50:65:@4387.4]
  assign _T_4369 = _T_4345 + _T_4346; // @[Bitwise.scala 48:55:@4388.4]
  assign _GEN_628 = {{1'd0}, _T_4344}; // @[Bitwise.scala 48:55:@4389.4]
  assign _T_4370 = _GEN_628 + _T_4369; // @[Bitwise.scala 48:55:@4389.4]
  assign _T_4371 = _T_4348 + _T_4349; // @[Bitwise.scala 48:55:@4390.4]
  assign _GEN_629 = {{1'd0}, _T_4347}; // @[Bitwise.scala 48:55:@4391.4]
  assign _T_4372 = _GEN_629 + _T_4371; // @[Bitwise.scala 48:55:@4391.4]
  assign _T_4373 = _T_4370 + _T_4372; // @[Bitwise.scala 48:55:@4392.4]
  assign _T_4374 = _T_4351 + _T_4352; // @[Bitwise.scala 48:55:@4393.4]
  assign _GEN_630 = {{1'd0}, _T_4350}; // @[Bitwise.scala 48:55:@4394.4]
  assign _T_4375 = _GEN_630 + _T_4374; // @[Bitwise.scala 48:55:@4394.4]
  assign _T_4376 = _T_4354 + _T_4355; // @[Bitwise.scala 48:55:@4395.4]
  assign _GEN_631 = {{1'd0}, _T_4353}; // @[Bitwise.scala 48:55:@4396.4]
  assign _T_4377 = _GEN_631 + _T_4376; // @[Bitwise.scala 48:55:@4396.4]
  assign _T_4378 = _T_4375 + _T_4377; // @[Bitwise.scala 48:55:@4397.4]
  assign _T_4379 = _T_4373 + _T_4378; // @[Bitwise.scala 48:55:@4398.4]
  assign _T_4380 = _T_4357 + _T_4358; // @[Bitwise.scala 48:55:@4399.4]
  assign _GEN_632 = {{1'd0}, _T_4356}; // @[Bitwise.scala 48:55:@4400.4]
  assign _T_4381 = _GEN_632 + _T_4380; // @[Bitwise.scala 48:55:@4400.4]
  assign _T_4382 = _T_4360 + _T_4361; // @[Bitwise.scala 48:55:@4401.4]
  assign _GEN_633 = {{1'd0}, _T_4359}; // @[Bitwise.scala 48:55:@4402.4]
  assign _T_4383 = _GEN_633 + _T_4382; // @[Bitwise.scala 48:55:@4402.4]
  assign _T_4384 = _T_4381 + _T_4383; // @[Bitwise.scala 48:55:@4403.4]
  assign _T_4385 = _T_4363 + _T_4364; // @[Bitwise.scala 48:55:@4404.4]
  assign _GEN_634 = {{1'd0}, _T_4362}; // @[Bitwise.scala 48:55:@4405.4]
  assign _T_4386 = _GEN_634 + _T_4385; // @[Bitwise.scala 48:55:@4405.4]
  assign _T_4387 = _T_4365 + _T_4366; // @[Bitwise.scala 48:55:@4406.4]
  assign _T_4388 = _T_4367 + _T_4368; // @[Bitwise.scala 48:55:@4407.4]
  assign _T_4389 = _T_4387 + _T_4388; // @[Bitwise.scala 48:55:@4408.4]
  assign _T_4390 = _T_4386 + _T_4389; // @[Bitwise.scala 48:55:@4409.4]
  assign _T_4391 = _T_4384 + _T_4390; // @[Bitwise.scala 48:55:@4410.4]
  assign _T_4392 = _T_4379 + _T_4391; // @[Bitwise.scala 48:55:@4411.4]
  assign _T_4456 = _T_2230[25:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4476.4]
  assign _T_4457 = _T_4456[0]; // @[Bitwise.scala 50:65:@4477.4]
  assign _T_4458 = _T_4456[1]; // @[Bitwise.scala 50:65:@4478.4]
  assign _T_4459 = _T_4456[2]; // @[Bitwise.scala 50:65:@4479.4]
  assign _T_4460 = _T_4456[3]; // @[Bitwise.scala 50:65:@4480.4]
  assign _T_4461 = _T_4456[4]; // @[Bitwise.scala 50:65:@4481.4]
  assign _T_4462 = _T_4456[5]; // @[Bitwise.scala 50:65:@4482.4]
  assign _T_4463 = _T_4456[6]; // @[Bitwise.scala 50:65:@4483.4]
  assign _T_4464 = _T_4456[7]; // @[Bitwise.scala 50:65:@4484.4]
  assign _T_4465 = _T_4456[8]; // @[Bitwise.scala 50:65:@4485.4]
  assign _T_4466 = _T_4456[9]; // @[Bitwise.scala 50:65:@4486.4]
  assign _T_4467 = _T_4456[10]; // @[Bitwise.scala 50:65:@4487.4]
  assign _T_4468 = _T_4456[11]; // @[Bitwise.scala 50:65:@4488.4]
  assign _T_4469 = _T_4456[12]; // @[Bitwise.scala 50:65:@4489.4]
  assign _T_4470 = _T_4456[13]; // @[Bitwise.scala 50:65:@4490.4]
  assign _T_4471 = _T_4456[14]; // @[Bitwise.scala 50:65:@4491.4]
  assign _T_4472 = _T_4456[15]; // @[Bitwise.scala 50:65:@4492.4]
  assign _T_4473 = _T_4456[16]; // @[Bitwise.scala 50:65:@4493.4]
  assign _T_4474 = _T_4456[17]; // @[Bitwise.scala 50:65:@4494.4]
  assign _T_4475 = _T_4456[18]; // @[Bitwise.scala 50:65:@4495.4]
  assign _T_4476 = _T_4456[19]; // @[Bitwise.scala 50:65:@4496.4]
  assign _T_4477 = _T_4456[20]; // @[Bitwise.scala 50:65:@4497.4]
  assign _T_4478 = _T_4456[21]; // @[Bitwise.scala 50:65:@4498.4]
  assign _T_4479 = _T_4456[22]; // @[Bitwise.scala 50:65:@4499.4]
  assign _T_4480 = _T_4456[23]; // @[Bitwise.scala 50:65:@4500.4]
  assign _T_4481 = _T_4456[24]; // @[Bitwise.scala 50:65:@4501.4]
  assign _T_4482 = _T_4456[25]; // @[Bitwise.scala 50:65:@4502.4]
  assign _T_4483 = _T_4458 + _T_4459; // @[Bitwise.scala 48:55:@4503.4]
  assign _GEN_635 = {{1'd0}, _T_4457}; // @[Bitwise.scala 48:55:@4504.4]
  assign _T_4484 = _GEN_635 + _T_4483; // @[Bitwise.scala 48:55:@4504.4]
  assign _T_4485 = _T_4461 + _T_4462; // @[Bitwise.scala 48:55:@4505.4]
  assign _GEN_636 = {{1'd0}, _T_4460}; // @[Bitwise.scala 48:55:@4506.4]
  assign _T_4486 = _GEN_636 + _T_4485; // @[Bitwise.scala 48:55:@4506.4]
  assign _T_4487 = _T_4484 + _T_4486; // @[Bitwise.scala 48:55:@4507.4]
  assign _T_4488 = _T_4464 + _T_4465; // @[Bitwise.scala 48:55:@4508.4]
  assign _GEN_637 = {{1'd0}, _T_4463}; // @[Bitwise.scala 48:55:@4509.4]
  assign _T_4489 = _GEN_637 + _T_4488; // @[Bitwise.scala 48:55:@4509.4]
  assign _T_4490 = _T_4466 + _T_4467; // @[Bitwise.scala 48:55:@4510.4]
  assign _T_4491 = _T_4468 + _T_4469; // @[Bitwise.scala 48:55:@4511.4]
  assign _T_4492 = _T_4490 + _T_4491; // @[Bitwise.scala 48:55:@4512.4]
  assign _T_4493 = _T_4489 + _T_4492; // @[Bitwise.scala 48:55:@4513.4]
  assign _T_4494 = _T_4487 + _T_4493; // @[Bitwise.scala 48:55:@4514.4]
  assign _T_4495 = _T_4471 + _T_4472; // @[Bitwise.scala 48:55:@4515.4]
  assign _GEN_638 = {{1'd0}, _T_4470}; // @[Bitwise.scala 48:55:@4516.4]
  assign _T_4496 = _GEN_638 + _T_4495; // @[Bitwise.scala 48:55:@4516.4]
  assign _T_4497 = _T_4474 + _T_4475; // @[Bitwise.scala 48:55:@4517.4]
  assign _GEN_639 = {{1'd0}, _T_4473}; // @[Bitwise.scala 48:55:@4518.4]
  assign _T_4498 = _GEN_639 + _T_4497; // @[Bitwise.scala 48:55:@4518.4]
  assign _T_4499 = _T_4496 + _T_4498; // @[Bitwise.scala 48:55:@4519.4]
  assign _T_4500 = _T_4477 + _T_4478; // @[Bitwise.scala 48:55:@4520.4]
  assign _GEN_640 = {{1'd0}, _T_4476}; // @[Bitwise.scala 48:55:@4521.4]
  assign _T_4501 = _GEN_640 + _T_4500; // @[Bitwise.scala 48:55:@4521.4]
  assign _T_4502 = _T_4479 + _T_4480; // @[Bitwise.scala 48:55:@4522.4]
  assign _T_4503 = _T_4481 + _T_4482; // @[Bitwise.scala 48:55:@4523.4]
  assign _T_4504 = _T_4502 + _T_4503; // @[Bitwise.scala 48:55:@4524.4]
  assign _T_4505 = _T_4501 + _T_4504; // @[Bitwise.scala 48:55:@4525.4]
  assign _T_4506 = _T_4499 + _T_4505; // @[Bitwise.scala 48:55:@4526.4]
  assign _T_4507 = _T_4494 + _T_4506; // @[Bitwise.scala 48:55:@4527.4]
  assign _T_4571 = _T_2230[26:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4592.4]
  assign _T_4572 = _T_4571[0]; // @[Bitwise.scala 50:65:@4593.4]
  assign _T_4573 = _T_4571[1]; // @[Bitwise.scala 50:65:@4594.4]
  assign _T_4574 = _T_4571[2]; // @[Bitwise.scala 50:65:@4595.4]
  assign _T_4575 = _T_4571[3]; // @[Bitwise.scala 50:65:@4596.4]
  assign _T_4576 = _T_4571[4]; // @[Bitwise.scala 50:65:@4597.4]
  assign _T_4577 = _T_4571[5]; // @[Bitwise.scala 50:65:@4598.4]
  assign _T_4578 = _T_4571[6]; // @[Bitwise.scala 50:65:@4599.4]
  assign _T_4579 = _T_4571[7]; // @[Bitwise.scala 50:65:@4600.4]
  assign _T_4580 = _T_4571[8]; // @[Bitwise.scala 50:65:@4601.4]
  assign _T_4581 = _T_4571[9]; // @[Bitwise.scala 50:65:@4602.4]
  assign _T_4582 = _T_4571[10]; // @[Bitwise.scala 50:65:@4603.4]
  assign _T_4583 = _T_4571[11]; // @[Bitwise.scala 50:65:@4604.4]
  assign _T_4584 = _T_4571[12]; // @[Bitwise.scala 50:65:@4605.4]
  assign _T_4585 = _T_4571[13]; // @[Bitwise.scala 50:65:@4606.4]
  assign _T_4586 = _T_4571[14]; // @[Bitwise.scala 50:65:@4607.4]
  assign _T_4587 = _T_4571[15]; // @[Bitwise.scala 50:65:@4608.4]
  assign _T_4588 = _T_4571[16]; // @[Bitwise.scala 50:65:@4609.4]
  assign _T_4589 = _T_4571[17]; // @[Bitwise.scala 50:65:@4610.4]
  assign _T_4590 = _T_4571[18]; // @[Bitwise.scala 50:65:@4611.4]
  assign _T_4591 = _T_4571[19]; // @[Bitwise.scala 50:65:@4612.4]
  assign _T_4592 = _T_4571[20]; // @[Bitwise.scala 50:65:@4613.4]
  assign _T_4593 = _T_4571[21]; // @[Bitwise.scala 50:65:@4614.4]
  assign _T_4594 = _T_4571[22]; // @[Bitwise.scala 50:65:@4615.4]
  assign _T_4595 = _T_4571[23]; // @[Bitwise.scala 50:65:@4616.4]
  assign _T_4596 = _T_4571[24]; // @[Bitwise.scala 50:65:@4617.4]
  assign _T_4597 = _T_4571[25]; // @[Bitwise.scala 50:65:@4618.4]
  assign _T_4598 = _T_4571[26]; // @[Bitwise.scala 50:65:@4619.4]
  assign _T_4599 = _T_4573 + _T_4574; // @[Bitwise.scala 48:55:@4620.4]
  assign _GEN_641 = {{1'd0}, _T_4572}; // @[Bitwise.scala 48:55:@4621.4]
  assign _T_4600 = _GEN_641 + _T_4599; // @[Bitwise.scala 48:55:@4621.4]
  assign _T_4601 = _T_4576 + _T_4577; // @[Bitwise.scala 48:55:@4622.4]
  assign _GEN_642 = {{1'd0}, _T_4575}; // @[Bitwise.scala 48:55:@4623.4]
  assign _T_4602 = _GEN_642 + _T_4601; // @[Bitwise.scala 48:55:@4623.4]
  assign _T_4603 = _T_4600 + _T_4602; // @[Bitwise.scala 48:55:@4624.4]
  assign _T_4604 = _T_4579 + _T_4580; // @[Bitwise.scala 48:55:@4625.4]
  assign _GEN_643 = {{1'd0}, _T_4578}; // @[Bitwise.scala 48:55:@4626.4]
  assign _T_4605 = _GEN_643 + _T_4604; // @[Bitwise.scala 48:55:@4626.4]
  assign _T_4606 = _T_4581 + _T_4582; // @[Bitwise.scala 48:55:@4627.4]
  assign _T_4607 = _T_4583 + _T_4584; // @[Bitwise.scala 48:55:@4628.4]
  assign _T_4608 = _T_4606 + _T_4607; // @[Bitwise.scala 48:55:@4629.4]
  assign _T_4609 = _T_4605 + _T_4608; // @[Bitwise.scala 48:55:@4630.4]
  assign _T_4610 = _T_4603 + _T_4609; // @[Bitwise.scala 48:55:@4631.4]
  assign _T_4611 = _T_4586 + _T_4587; // @[Bitwise.scala 48:55:@4632.4]
  assign _GEN_644 = {{1'd0}, _T_4585}; // @[Bitwise.scala 48:55:@4633.4]
  assign _T_4612 = _GEN_644 + _T_4611; // @[Bitwise.scala 48:55:@4633.4]
  assign _T_4613 = _T_4588 + _T_4589; // @[Bitwise.scala 48:55:@4634.4]
  assign _T_4614 = _T_4590 + _T_4591; // @[Bitwise.scala 48:55:@4635.4]
  assign _T_4615 = _T_4613 + _T_4614; // @[Bitwise.scala 48:55:@4636.4]
  assign _T_4616 = _T_4612 + _T_4615; // @[Bitwise.scala 48:55:@4637.4]
  assign _T_4617 = _T_4593 + _T_4594; // @[Bitwise.scala 48:55:@4638.4]
  assign _GEN_645 = {{1'd0}, _T_4592}; // @[Bitwise.scala 48:55:@4639.4]
  assign _T_4618 = _GEN_645 + _T_4617; // @[Bitwise.scala 48:55:@4639.4]
  assign _T_4619 = _T_4595 + _T_4596; // @[Bitwise.scala 48:55:@4640.4]
  assign _T_4620 = _T_4597 + _T_4598; // @[Bitwise.scala 48:55:@4641.4]
  assign _T_4621 = _T_4619 + _T_4620; // @[Bitwise.scala 48:55:@4642.4]
  assign _T_4622 = _T_4618 + _T_4621; // @[Bitwise.scala 48:55:@4643.4]
  assign _T_4623 = _T_4616 + _T_4622; // @[Bitwise.scala 48:55:@4644.4]
  assign _T_4624 = _T_4610 + _T_4623; // @[Bitwise.scala 48:55:@4645.4]
  assign _T_4688 = _T_2230[27:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4710.4]
  assign _T_4689 = _T_4688[0]; // @[Bitwise.scala 50:65:@4711.4]
  assign _T_4690 = _T_4688[1]; // @[Bitwise.scala 50:65:@4712.4]
  assign _T_4691 = _T_4688[2]; // @[Bitwise.scala 50:65:@4713.4]
  assign _T_4692 = _T_4688[3]; // @[Bitwise.scala 50:65:@4714.4]
  assign _T_4693 = _T_4688[4]; // @[Bitwise.scala 50:65:@4715.4]
  assign _T_4694 = _T_4688[5]; // @[Bitwise.scala 50:65:@4716.4]
  assign _T_4695 = _T_4688[6]; // @[Bitwise.scala 50:65:@4717.4]
  assign _T_4696 = _T_4688[7]; // @[Bitwise.scala 50:65:@4718.4]
  assign _T_4697 = _T_4688[8]; // @[Bitwise.scala 50:65:@4719.4]
  assign _T_4698 = _T_4688[9]; // @[Bitwise.scala 50:65:@4720.4]
  assign _T_4699 = _T_4688[10]; // @[Bitwise.scala 50:65:@4721.4]
  assign _T_4700 = _T_4688[11]; // @[Bitwise.scala 50:65:@4722.4]
  assign _T_4701 = _T_4688[12]; // @[Bitwise.scala 50:65:@4723.4]
  assign _T_4702 = _T_4688[13]; // @[Bitwise.scala 50:65:@4724.4]
  assign _T_4703 = _T_4688[14]; // @[Bitwise.scala 50:65:@4725.4]
  assign _T_4704 = _T_4688[15]; // @[Bitwise.scala 50:65:@4726.4]
  assign _T_4705 = _T_4688[16]; // @[Bitwise.scala 50:65:@4727.4]
  assign _T_4706 = _T_4688[17]; // @[Bitwise.scala 50:65:@4728.4]
  assign _T_4707 = _T_4688[18]; // @[Bitwise.scala 50:65:@4729.4]
  assign _T_4708 = _T_4688[19]; // @[Bitwise.scala 50:65:@4730.4]
  assign _T_4709 = _T_4688[20]; // @[Bitwise.scala 50:65:@4731.4]
  assign _T_4710 = _T_4688[21]; // @[Bitwise.scala 50:65:@4732.4]
  assign _T_4711 = _T_4688[22]; // @[Bitwise.scala 50:65:@4733.4]
  assign _T_4712 = _T_4688[23]; // @[Bitwise.scala 50:65:@4734.4]
  assign _T_4713 = _T_4688[24]; // @[Bitwise.scala 50:65:@4735.4]
  assign _T_4714 = _T_4688[25]; // @[Bitwise.scala 50:65:@4736.4]
  assign _T_4715 = _T_4688[26]; // @[Bitwise.scala 50:65:@4737.4]
  assign _T_4716 = _T_4688[27]; // @[Bitwise.scala 50:65:@4738.4]
  assign _T_4717 = _T_4690 + _T_4691; // @[Bitwise.scala 48:55:@4739.4]
  assign _GEN_646 = {{1'd0}, _T_4689}; // @[Bitwise.scala 48:55:@4740.4]
  assign _T_4718 = _GEN_646 + _T_4717; // @[Bitwise.scala 48:55:@4740.4]
  assign _T_4719 = _T_4692 + _T_4693; // @[Bitwise.scala 48:55:@4741.4]
  assign _T_4720 = _T_4694 + _T_4695; // @[Bitwise.scala 48:55:@4742.4]
  assign _T_4721 = _T_4719 + _T_4720; // @[Bitwise.scala 48:55:@4743.4]
  assign _T_4722 = _T_4718 + _T_4721; // @[Bitwise.scala 48:55:@4744.4]
  assign _T_4723 = _T_4697 + _T_4698; // @[Bitwise.scala 48:55:@4745.4]
  assign _GEN_647 = {{1'd0}, _T_4696}; // @[Bitwise.scala 48:55:@4746.4]
  assign _T_4724 = _GEN_647 + _T_4723; // @[Bitwise.scala 48:55:@4746.4]
  assign _T_4725 = _T_4699 + _T_4700; // @[Bitwise.scala 48:55:@4747.4]
  assign _T_4726 = _T_4701 + _T_4702; // @[Bitwise.scala 48:55:@4748.4]
  assign _T_4727 = _T_4725 + _T_4726; // @[Bitwise.scala 48:55:@4749.4]
  assign _T_4728 = _T_4724 + _T_4727; // @[Bitwise.scala 48:55:@4750.4]
  assign _T_4729 = _T_4722 + _T_4728; // @[Bitwise.scala 48:55:@4751.4]
  assign _T_4730 = _T_4704 + _T_4705; // @[Bitwise.scala 48:55:@4752.4]
  assign _GEN_648 = {{1'd0}, _T_4703}; // @[Bitwise.scala 48:55:@4753.4]
  assign _T_4731 = _GEN_648 + _T_4730; // @[Bitwise.scala 48:55:@4753.4]
  assign _T_4732 = _T_4706 + _T_4707; // @[Bitwise.scala 48:55:@4754.4]
  assign _T_4733 = _T_4708 + _T_4709; // @[Bitwise.scala 48:55:@4755.4]
  assign _T_4734 = _T_4732 + _T_4733; // @[Bitwise.scala 48:55:@4756.4]
  assign _T_4735 = _T_4731 + _T_4734; // @[Bitwise.scala 48:55:@4757.4]
  assign _T_4736 = _T_4711 + _T_4712; // @[Bitwise.scala 48:55:@4758.4]
  assign _GEN_649 = {{1'd0}, _T_4710}; // @[Bitwise.scala 48:55:@4759.4]
  assign _T_4737 = _GEN_649 + _T_4736; // @[Bitwise.scala 48:55:@4759.4]
  assign _T_4738 = _T_4713 + _T_4714; // @[Bitwise.scala 48:55:@4760.4]
  assign _T_4739 = _T_4715 + _T_4716; // @[Bitwise.scala 48:55:@4761.4]
  assign _T_4740 = _T_4738 + _T_4739; // @[Bitwise.scala 48:55:@4762.4]
  assign _T_4741 = _T_4737 + _T_4740; // @[Bitwise.scala 48:55:@4763.4]
  assign _T_4742 = _T_4735 + _T_4741; // @[Bitwise.scala 48:55:@4764.4]
  assign _T_4743 = _T_4729 + _T_4742; // @[Bitwise.scala 48:55:@4765.4]
  assign _T_4807 = _T_2230[28:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4830.4]
  assign _T_4808 = _T_4807[0]; // @[Bitwise.scala 50:65:@4831.4]
  assign _T_4809 = _T_4807[1]; // @[Bitwise.scala 50:65:@4832.4]
  assign _T_4810 = _T_4807[2]; // @[Bitwise.scala 50:65:@4833.4]
  assign _T_4811 = _T_4807[3]; // @[Bitwise.scala 50:65:@4834.4]
  assign _T_4812 = _T_4807[4]; // @[Bitwise.scala 50:65:@4835.4]
  assign _T_4813 = _T_4807[5]; // @[Bitwise.scala 50:65:@4836.4]
  assign _T_4814 = _T_4807[6]; // @[Bitwise.scala 50:65:@4837.4]
  assign _T_4815 = _T_4807[7]; // @[Bitwise.scala 50:65:@4838.4]
  assign _T_4816 = _T_4807[8]; // @[Bitwise.scala 50:65:@4839.4]
  assign _T_4817 = _T_4807[9]; // @[Bitwise.scala 50:65:@4840.4]
  assign _T_4818 = _T_4807[10]; // @[Bitwise.scala 50:65:@4841.4]
  assign _T_4819 = _T_4807[11]; // @[Bitwise.scala 50:65:@4842.4]
  assign _T_4820 = _T_4807[12]; // @[Bitwise.scala 50:65:@4843.4]
  assign _T_4821 = _T_4807[13]; // @[Bitwise.scala 50:65:@4844.4]
  assign _T_4822 = _T_4807[14]; // @[Bitwise.scala 50:65:@4845.4]
  assign _T_4823 = _T_4807[15]; // @[Bitwise.scala 50:65:@4846.4]
  assign _T_4824 = _T_4807[16]; // @[Bitwise.scala 50:65:@4847.4]
  assign _T_4825 = _T_4807[17]; // @[Bitwise.scala 50:65:@4848.4]
  assign _T_4826 = _T_4807[18]; // @[Bitwise.scala 50:65:@4849.4]
  assign _T_4827 = _T_4807[19]; // @[Bitwise.scala 50:65:@4850.4]
  assign _T_4828 = _T_4807[20]; // @[Bitwise.scala 50:65:@4851.4]
  assign _T_4829 = _T_4807[21]; // @[Bitwise.scala 50:65:@4852.4]
  assign _T_4830 = _T_4807[22]; // @[Bitwise.scala 50:65:@4853.4]
  assign _T_4831 = _T_4807[23]; // @[Bitwise.scala 50:65:@4854.4]
  assign _T_4832 = _T_4807[24]; // @[Bitwise.scala 50:65:@4855.4]
  assign _T_4833 = _T_4807[25]; // @[Bitwise.scala 50:65:@4856.4]
  assign _T_4834 = _T_4807[26]; // @[Bitwise.scala 50:65:@4857.4]
  assign _T_4835 = _T_4807[27]; // @[Bitwise.scala 50:65:@4858.4]
  assign _T_4836 = _T_4807[28]; // @[Bitwise.scala 50:65:@4859.4]
  assign _T_4837 = _T_4809 + _T_4810; // @[Bitwise.scala 48:55:@4860.4]
  assign _GEN_650 = {{1'd0}, _T_4808}; // @[Bitwise.scala 48:55:@4861.4]
  assign _T_4838 = _GEN_650 + _T_4837; // @[Bitwise.scala 48:55:@4861.4]
  assign _T_4839 = _T_4811 + _T_4812; // @[Bitwise.scala 48:55:@4862.4]
  assign _T_4840 = _T_4813 + _T_4814; // @[Bitwise.scala 48:55:@4863.4]
  assign _T_4841 = _T_4839 + _T_4840; // @[Bitwise.scala 48:55:@4864.4]
  assign _T_4842 = _T_4838 + _T_4841; // @[Bitwise.scala 48:55:@4865.4]
  assign _T_4843 = _T_4816 + _T_4817; // @[Bitwise.scala 48:55:@4866.4]
  assign _GEN_651 = {{1'd0}, _T_4815}; // @[Bitwise.scala 48:55:@4867.4]
  assign _T_4844 = _GEN_651 + _T_4843; // @[Bitwise.scala 48:55:@4867.4]
  assign _T_4845 = _T_4818 + _T_4819; // @[Bitwise.scala 48:55:@4868.4]
  assign _T_4846 = _T_4820 + _T_4821; // @[Bitwise.scala 48:55:@4869.4]
  assign _T_4847 = _T_4845 + _T_4846; // @[Bitwise.scala 48:55:@4870.4]
  assign _T_4848 = _T_4844 + _T_4847; // @[Bitwise.scala 48:55:@4871.4]
  assign _T_4849 = _T_4842 + _T_4848; // @[Bitwise.scala 48:55:@4872.4]
  assign _T_4850 = _T_4823 + _T_4824; // @[Bitwise.scala 48:55:@4873.4]
  assign _GEN_652 = {{1'd0}, _T_4822}; // @[Bitwise.scala 48:55:@4874.4]
  assign _T_4851 = _GEN_652 + _T_4850; // @[Bitwise.scala 48:55:@4874.4]
  assign _T_4852 = _T_4825 + _T_4826; // @[Bitwise.scala 48:55:@4875.4]
  assign _T_4853 = _T_4827 + _T_4828; // @[Bitwise.scala 48:55:@4876.4]
  assign _T_4854 = _T_4852 + _T_4853; // @[Bitwise.scala 48:55:@4877.4]
  assign _T_4855 = _T_4851 + _T_4854; // @[Bitwise.scala 48:55:@4878.4]
  assign _T_4856 = _T_4829 + _T_4830; // @[Bitwise.scala 48:55:@4879.4]
  assign _T_4857 = _T_4831 + _T_4832; // @[Bitwise.scala 48:55:@4880.4]
  assign _T_4858 = _T_4856 + _T_4857; // @[Bitwise.scala 48:55:@4881.4]
  assign _T_4859 = _T_4833 + _T_4834; // @[Bitwise.scala 48:55:@4882.4]
  assign _T_4860 = _T_4835 + _T_4836; // @[Bitwise.scala 48:55:@4883.4]
  assign _T_4861 = _T_4859 + _T_4860; // @[Bitwise.scala 48:55:@4884.4]
  assign _T_4862 = _T_4858 + _T_4861; // @[Bitwise.scala 48:55:@4885.4]
  assign _T_4863 = _T_4855 + _T_4862; // @[Bitwise.scala 48:55:@4886.4]
  assign _T_4864 = _T_4849 + _T_4863; // @[Bitwise.scala 48:55:@4887.4]
  assign _T_4928 = _T_2230[29:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4952.4]
  assign _T_4929 = _T_4928[0]; // @[Bitwise.scala 50:65:@4953.4]
  assign _T_4930 = _T_4928[1]; // @[Bitwise.scala 50:65:@4954.4]
  assign _T_4931 = _T_4928[2]; // @[Bitwise.scala 50:65:@4955.4]
  assign _T_4932 = _T_4928[3]; // @[Bitwise.scala 50:65:@4956.4]
  assign _T_4933 = _T_4928[4]; // @[Bitwise.scala 50:65:@4957.4]
  assign _T_4934 = _T_4928[5]; // @[Bitwise.scala 50:65:@4958.4]
  assign _T_4935 = _T_4928[6]; // @[Bitwise.scala 50:65:@4959.4]
  assign _T_4936 = _T_4928[7]; // @[Bitwise.scala 50:65:@4960.4]
  assign _T_4937 = _T_4928[8]; // @[Bitwise.scala 50:65:@4961.4]
  assign _T_4938 = _T_4928[9]; // @[Bitwise.scala 50:65:@4962.4]
  assign _T_4939 = _T_4928[10]; // @[Bitwise.scala 50:65:@4963.4]
  assign _T_4940 = _T_4928[11]; // @[Bitwise.scala 50:65:@4964.4]
  assign _T_4941 = _T_4928[12]; // @[Bitwise.scala 50:65:@4965.4]
  assign _T_4942 = _T_4928[13]; // @[Bitwise.scala 50:65:@4966.4]
  assign _T_4943 = _T_4928[14]; // @[Bitwise.scala 50:65:@4967.4]
  assign _T_4944 = _T_4928[15]; // @[Bitwise.scala 50:65:@4968.4]
  assign _T_4945 = _T_4928[16]; // @[Bitwise.scala 50:65:@4969.4]
  assign _T_4946 = _T_4928[17]; // @[Bitwise.scala 50:65:@4970.4]
  assign _T_4947 = _T_4928[18]; // @[Bitwise.scala 50:65:@4971.4]
  assign _T_4948 = _T_4928[19]; // @[Bitwise.scala 50:65:@4972.4]
  assign _T_4949 = _T_4928[20]; // @[Bitwise.scala 50:65:@4973.4]
  assign _T_4950 = _T_4928[21]; // @[Bitwise.scala 50:65:@4974.4]
  assign _T_4951 = _T_4928[22]; // @[Bitwise.scala 50:65:@4975.4]
  assign _T_4952 = _T_4928[23]; // @[Bitwise.scala 50:65:@4976.4]
  assign _T_4953 = _T_4928[24]; // @[Bitwise.scala 50:65:@4977.4]
  assign _T_4954 = _T_4928[25]; // @[Bitwise.scala 50:65:@4978.4]
  assign _T_4955 = _T_4928[26]; // @[Bitwise.scala 50:65:@4979.4]
  assign _T_4956 = _T_4928[27]; // @[Bitwise.scala 50:65:@4980.4]
  assign _T_4957 = _T_4928[28]; // @[Bitwise.scala 50:65:@4981.4]
  assign _T_4958 = _T_4928[29]; // @[Bitwise.scala 50:65:@4982.4]
  assign _T_4959 = _T_4930 + _T_4931; // @[Bitwise.scala 48:55:@4983.4]
  assign _GEN_653 = {{1'd0}, _T_4929}; // @[Bitwise.scala 48:55:@4984.4]
  assign _T_4960 = _GEN_653 + _T_4959; // @[Bitwise.scala 48:55:@4984.4]
  assign _T_4961 = _T_4932 + _T_4933; // @[Bitwise.scala 48:55:@4985.4]
  assign _T_4962 = _T_4934 + _T_4935; // @[Bitwise.scala 48:55:@4986.4]
  assign _T_4963 = _T_4961 + _T_4962; // @[Bitwise.scala 48:55:@4987.4]
  assign _T_4964 = _T_4960 + _T_4963; // @[Bitwise.scala 48:55:@4988.4]
  assign _T_4965 = _T_4936 + _T_4937; // @[Bitwise.scala 48:55:@4989.4]
  assign _T_4966 = _T_4938 + _T_4939; // @[Bitwise.scala 48:55:@4990.4]
  assign _T_4967 = _T_4965 + _T_4966; // @[Bitwise.scala 48:55:@4991.4]
  assign _T_4968 = _T_4940 + _T_4941; // @[Bitwise.scala 48:55:@4992.4]
  assign _T_4969 = _T_4942 + _T_4943; // @[Bitwise.scala 48:55:@4993.4]
  assign _T_4970 = _T_4968 + _T_4969; // @[Bitwise.scala 48:55:@4994.4]
  assign _T_4971 = _T_4967 + _T_4970; // @[Bitwise.scala 48:55:@4995.4]
  assign _T_4972 = _T_4964 + _T_4971; // @[Bitwise.scala 48:55:@4996.4]
  assign _T_4973 = _T_4945 + _T_4946; // @[Bitwise.scala 48:55:@4997.4]
  assign _GEN_654 = {{1'd0}, _T_4944}; // @[Bitwise.scala 48:55:@4998.4]
  assign _T_4974 = _GEN_654 + _T_4973; // @[Bitwise.scala 48:55:@4998.4]
  assign _T_4975 = _T_4947 + _T_4948; // @[Bitwise.scala 48:55:@4999.4]
  assign _T_4976 = _T_4949 + _T_4950; // @[Bitwise.scala 48:55:@5000.4]
  assign _T_4977 = _T_4975 + _T_4976; // @[Bitwise.scala 48:55:@5001.4]
  assign _T_4978 = _T_4974 + _T_4977; // @[Bitwise.scala 48:55:@5002.4]
  assign _T_4979 = _T_4951 + _T_4952; // @[Bitwise.scala 48:55:@5003.4]
  assign _T_4980 = _T_4953 + _T_4954; // @[Bitwise.scala 48:55:@5004.4]
  assign _T_4981 = _T_4979 + _T_4980; // @[Bitwise.scala 48:55:@5005.4]
  assign _T_4982 = _T_4955 + _T_4956; // @[Bitwise.scala 48:55:@5006.4]
  assign _T_4983 = _T_4957 + _T_4958; // @[Bitwise.scala 48:55:@5007.4]
  assign _T_4984 = _T_4982 + _T_4983; // @[Bitwise.scala 48:55:@5008.4]
  assign _T_4985 = _T_4981 + _T_4984; // @[Bitwise.scala 48:55:@5009.4]
  assign _T_4986 = _T_4978 + _T_4985; // @[Bitwise.scala 48:55:@5010.4]
  assign _T_4987 = _T_4972 + _T_4986; // @[Bitwise.scala 48:55:@5011.4]
  assign _T_5051 = _T_2230[30:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5076.4]
  assign _T_5052 = _T_5051[0]; // @[Bitwise.scala 50:65:@5077.4]
  assign _T_5053 = _T_5051[1]; // @[Bitwise.scala 50:65:@5078.4]
  assign _T_5054 = _T_5051[2]; // @[Bitwise.scala 50:65:@5079.4]
  assign _T_5055 = _T_5051[3]; // @[Bitwise.scala 50:65:@5080.4]
  assign _T_5056 = _T_5051[4]; // @[Bitwise.scala 50:65:@5081.4]
  assign _T_5057 = _T_5051[5]; // @[Bitwise.scala 50:65:@5082.4]
  assign _T_5058 = _T_5051[6]; // @[Bitwise.scala 50:65:@5083.4]
  assign _T_5059 = _T_5051[7]; // @[Bitwise.scala 50:65:@5084.4]
  assign _T_5060 = _T_5051[8]; // @[Bitwise.scala 50:65:@5085.4]
  assign _T_5061 = _T_5051[9]; // @[Bitwise.scala 50:65:@5086.4]
  assign _T_5062 = _T_5051[10]; // @[Bitwise.scala 50:65:@5087.4]
  assign _T_5063 = _T_5051[11]; // @[Bitwise.scala 50:65:@5088.4]
  assign _T_5064 = _T_5051[12]; // @[Bitwise.scala 50:65:@5089.4]
  assign _T_5065 = _T_5051[13]; // @[Bitwise.scala 50:65:@5090.4]
  assign _T_5066 = _T_5051[14]; // @[Bitwise.scala 50:65:@5091.4]
  assign _T_5067 = _T_5051[15]; // @[Bitwise.scala 50:65:@5092.4]
  assign _T_5068 = _T_5051[16]; // @[Bitwise.scala 50:65:@5093.4]
  assign _T_5069 = _T_5051[17]; // @[Bitwise.scala 50:65:@5094.4]
  assign _T_5070 = _T_5051[18]; // @[Bitwise.scala 50:65:@5095.4]
  assign _T_5071 = _T_5051[19]; // @[Bitwise.scala 50:65:@5096.4]
  assign _T_5072 = _T_5051[20]; // @[Bitwise.scala 50:65:@5097.4]
  assign _T_5073 = _T_5051[21]; // @[Bitwise.scala 50:65:@5098.4]
  assign _T_5074 = _T_5051[22]; // @[Bitwise.scala 50:65:@5099.4]
  assign _T_5075 = _T_5051[23]; // @[Bitwise.scala 50:65:@5100.4]
  assign _T_5076 = _T_5051[24]; // @[Bitwise.scala 50:65:@5101.4]
  assign _T_5077 = _T_5051[25]; // @[Bitwise.scala 50:65:@5102.4]
  assign _T_5078 = _T_5051[26]; // @[Bitwise.scala 50:65:@5103.4]
  assign _T_5079 = _T_5051[27]; // @[Bitwise.scala 50:65:@5104.4]
  assign _T_5080 = _T_5051[28]; // @[Bitwise.scala 50:65:@5105.4]
  assign _T_5081 = _T_5051[29]; // @[Bitwise.scala 50:65:@5106.4]
  assign _T_5082 = _T_5051[30]; // @[Bitwise.scala 50:65:@5107.4]
  assign _T_5083 = _T_5053 + _T_5054; // @[Bitwise.scala 48:55:@5108.4]
  assign _GEN_655 = {{1'd0}, _T_5052}; // @[Bitwise.scala 48:55:@5109.4]
  assign _T_5084 = _GEN_655 + _T_5083; // @[Bitwise.scala 48:55:@5109.4]
  assign _T_5085 = _T_5055 + _T_5056; // @[Bitwise.scala 48:55:@5110.4]
  assign _T_5086 = _T_5057 + _T_5058; // @[Bitwise.scala 48:55:@5111.4]
  assign _T_5087 = _T_5085 + _T_5086; // @[Bitwise.scala 48:55:@5112.4]
  assign _T_5088 = _T_5084 + _T_5087; // @[Bitwise.scala 48:55:@5113.4]
  assign _T_5089 = _T_5059 + _T_5060; // @[Bitwise.scala 48:55:@5114.4]
  assign _T_5090 = _T_5061 + _T_5062; // @[Bitwise.scala 48:55:@5115.4]
  assign _T_5091 = _T_5089 + _T_5090; // @[Bitwise.scala 48:55:@5116.4]
  assign _T_5092 = _T_5063 + _T_5064; // @[Bitwise.scala 48:55:@5117.4]
  assign _T_5093 = _T_5065 + _T_5066; // @[Bitwise.scala 48:55:@5118.4]
  assign _T_5094 = _T_5092 + _T_5093; // @[Bitwise.scala 48:55:@5119.4]
  assign _T_5095 = _T_5091 + _T_5094; // @[Bitwise.scala 48:55:@5120.4]
  assign _T_5096 = _T_5088 + _T_5095; // @[Bitwise.scala 48:55:@5121.4]
  assign _T_5097 = _T_5067 + _T_5068; // @[Bitwise.scala 48:55:@5122.4]
  assign _T_5098 = _T_5069 + _T_5070; // @[Bitwise.scala 48:55:@5123.4]
  assign _T_5099 = _T_5097 + _T_5098; // @[Bitwise.scala 48:55:@5124.4]
  assign _T_5100 = _T_5071 + _T_5072; // @[Bitwise.scala 48:55:@5125.4]
  assign _T_5101 = _T_5073 + _T_5074; // @[Bitwise.scala 48:55:@5126.4]
  assign _T_5102 = _T_5100 + _T_5101; // @[Bitwise.scala 48:55:@5127.4]
  assign _T_5103 = _T_5099 + _T_5102; // @[Bitwise.scala 48:55:@5128.4]
  assign _T_5104 = _T_5075 + _T_5076; // @[Bitwise.scala 48:55:@5129.4]
  assign _T_5105 = _T_5077 + _T_5078; // @[Bitwise.scala 48:55:@5130.4]
  assign _T_5106 = _T_5104 + _T_5105; // @[Bitwise.scala 48:55:@5131.4]
  assign _T_5107 = _T_5079 + _T_5080; // @[Bitwise.scala 48:55:@5132.4]
  assign _T_5108 = _T_5081 + _T_5082; // @[Bitwise.scala 48:55:@5133.4]
  assign _T_5109 = _T_5107 + _T_5108; // @[Bitwise.scala 48:55:@5134.4]
  assign _T_5110 = _T_5106 + _T_5109; // @[Bitwise.scala 48:55:@5135.4]
  assign _T_5111 = _T_5103 + _T_5110; // @[Bitwise.scala 48:55:@5136.4]
  assign _T_5112 = _T_5096 + _T_5111; // @[Bitwise.scala 48:55:@5137.4]
  assign _T_5176 = _T_2230[31:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5202.4]
  assign _T_5177 = _T_5176[0]; // @[Bitwise.scala 50:65:@5203.4]
  assign _T_5178 = _T_5176[1]; // @[Bitwise.scala 50:65:@5204.4]
  assign _T_5179 = _T_5176[2]; // @[Bitwise.scala 50:65:@5205.4]
  assign _T_5180 = _T_5176[3]; // @[Bitwise.scala 50:65:@5206.4]
  assign _T_5181 = _T_5176[4]; // @[Bitwise.scala 50:65:@5207.4]
  assign _T_5182 = _T_5176[5]; // @[Bitwise.scala 50:65:@5208.4]
  assign _T_5183 = _T_5176[6]; // @[Bitwise.scala 50:65:@5209.4]
  assign _T_5184 = _T_5176[7]; // @[Bitwise.scala 50:65:@5210.4]
  assign _T_5185 = _T_5176[8]; // @[Bitwise.scala 50:65:@5211.4]
  assign _T_5186 = _T_5176[9]; // @[Bitwise.scala 50:65:@5212.4]
  assign _T_5187 = _T_5176[10]; // @[Bitwise.scala 50:65:@5213.4]
  assign _T_5188 = _T_5176[11]; // @[Bitwise.scala 50:65:@5214.4]
  assign _T_5189 = _T_5176[12]; // @[Bitwise.scala 50:65:@5215.4]
  assign _T_5190 = _T_5176[13]; // @[Bitwise.scala 50:65:@5216.4]
  assign _T_5191 = _T_5176[14]; // @[Bitwise.scala 50:65:@5217.4]
  assign _T_5192 = _T_5176[15]; // @[Bitwise.scala 50:65:@5218.4]
  assign _T_5193 = _T_5176[16]; // @[Bitwise.scala 50:65:@5219.4]
  assign _T_5194 = _T_5176[17]; // @[Bitwise.scala 50:65:@5220.4]
  assign _T_5195 = _T_5176[18]; // @[Bitwise.scala 50:65:@5221.4]
  assign _T_5196 = _T_5176[19]; // @[Bitwise.scala 50:65:@5222.4]
  assign _T_5197 = _T_5176[20]; // @[Bitwise.scala 50:65:@5223.4]
  assign _T_5198 = _T_5176[21]; // @[Bitwise.scala 50:65:@5224.4]
  assign _T_5199 = _T_5176[22]; // @[Bitwise.scala 50:65:@5225.4]
  assign _T_5200 = _T_5176[23]; // @[Bitwise.scala 50:65:@5226.4]
  assign _T_5201 = _T_5176[24]; // @[Bitwise.scala 50:65:@5227.4]
  assign _T_5202 = _T_5176[25]; // @[Bitwise.scala 50:65:@5228.4]
  assign _T_5203 = _T_5176[26]; // @[Bitwise.scala 50:65:@5229.4]
  assign _T_5204 = _T_5176[27]; // @[Bitwise.scala 50:65:@5230.4]
  assign _T_5205 = _T_5176[28]; // @[Bitwise.scala 50:65:@5231.4]
  assign _T_5206 = _T_5176[29]; // @[Bitwise.scala 50:65:@5232.4]
  assign _T_5207 = _T_5176[30]; // @[Bitwise.scala 50:65:@5233.4]
  assign _T_5208 = _T_5176[31]; // @[Bitwise.scala 50:65:@5234.4]
  assign _T_5209 = _T_5177 + _T_5178; // @[Bitwise.scala 48:55:@5235.4]
  assign _T_5210 = _T_5179 + _T_5180; // @[Bitwise.scala 48:55:@5236.4]
  assign _T_5211 = _T_5209 + _T_5210; // @[Bitwise.scala 48:55:@5237.4]
  assign _T_5212 = _T_5181 + _T_5182; // @[Bitwise.scala 48:55:@5238.4]
  assign _T_5213 = _T_5183 + _T_5184; // @[Bitwise.scala 48:55:@5239.4]
  assign _T_5214 = _T_5212 + _T_5213; // @[Bitwise.scala 48:55:@5240.4]
  assign _T_5215 = _T_5211 + _T_5214; // @[Bitwise.scala 48:55:@5241.4]
  assign _T_5216 = _T_5185 + _T_5186; // @[Bitwise.scala 48:55:@5242.4]
  assign _T_5217 = _T_5187 + _T_5188; // @[Bitwise.scala 48:55:@5243.4]
  assign _T_5218 = _T_5216 + _T_5217; // @[Bitwise.scala 48:55:@5244.4]
  assign _T_5219 = _T_5189 + _T_5190; // @[Bitwise.scala 48:55:@5245.4]
  assign _T_5220 = _T_5191 + _T_5192; // @[Bitwise.scala 48:55:@5246.4]
  assign _T_5221 = _T_5219 + _T_5220; // @[Bitwise.scala 48:55:@5247.4]
  assign _T_5222 = _T_5218 + _T_5221; // @[Bitwise.scala 48:55:@5248.4]
  assign _T_5223 = _T_5215 + _T_5222; // @[Bitwise.scala 48:55:@5249.4]
  assign _T_5224 = _T_5193 + _T_5194; // @[Bitwise.scala 48:55:@5250.4]
  assign _T_5225 = _T_5195 + _T_5196; // @[Bitwise.scala 48:55:@5251.4]
  assign _T_5226 = _T_5224 + _T_5225; // @[Bitwise.scala 48:55:@5252.4]
  assign _T_5227 = _T_5197 + _T_5198; // @[Bitwise.scala 48:55:@5253.4]
  assign _T_5228 = _T_5199 + _T_5200; // @[Bitwise.scala 48:55:@5254.4]
  assign _T_5229 = _T_5227 + _T_5228; // @[Bitwise.scala 48:55:@5255.4]
  assign _T_5230 = _T_5226 + _T_5229; // @[Bitwise.scala 48:55:@5256.4]
  assign _T_5231 = _T_5201 + _T_5202; // @[Bitwise.scala 48:55:@5257.4]
  assign _T_5232 = _T_5203 + _T_5204; // @[Bitwise.scala 48:55:@5258.4]
  assign _T_5233 = _T_5231 + _T_5232; // @[Bitwise.scala 48:55:@5259.4]
  assign _T_5234 = _T_5205 + _T_5206; // @[Bitwise.scala 48:55:@5260.4]
  assign _T_5235 = _T_5207 + _T_5208; // @[Bitwise.scala 48:55:@5261.4]
  assign _T_5236 = _T_5234 + _T_5235; // @[Bitwise.scala 48:55:@5262.4]
  assign _T_5237 = _T_5233 + _T_5236; // @[Bitwise.scala 48:55:@5263.4]
  assign _T_5238 = _T_5230 + _T_5237; // @[Bitwise.scala 48:55:@5264.4]
  assign _T_5239 = _T_5223 + _T_5238; // @[Bitwise.scala 48:55:@5265.4]
  assign _T_5303 = _T_2230[32:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5330.4]
  assign _T_5304 = _T_5303[0]; // @[Bitwise.scala 50:65:@5331.4]
  assign _T_5305 = _T_5303[1]; // @[Bitwise.scala 50:65:@5332.4]
  assign _T_5306 = _T_5303[2]; // @[Bitwise.scala 50:65:@5333.4]
  assign _T_5307 = _T_5303[3]; // @[Bitwise.scala 50:65:@5334.4]
  assign _T_5308 = _T_5303[4]; // @[Bitwise.scala 50:65:@5335.4]
  assign _T_5309 = _T_5303[5]; // @[Bitwise.scala 50:65:@5336.4]
  assign _T_5310 = _T_5303[6]; // @[Bitwise.scala 50:65:@5337.4]
  assign _T_5311 = _T_5303[7]; // @[Bitwise.scala 50:65:@5338.4]
  assign _T_5312 = _T_5303[8]; // @[Bitwise.scala 50:65:@5339.4]
  assign _T_5313 = _T_5303[9]; // @[Bitwise.scala 50:65:@5340.4]
  assign _T_5314 = _T_5303[10]; // @[Bitwise.scala 50:65:@5341.4]
  assign _T_5315 = _T_5303[11]; // @[Bitwise.scala 50:65:@5342.4]
  assign _T_5316 = _T_5303[12]; // @[Bitwise.scala 50:65:@5343.4]
  assign _T_5317 = _T_5303[13]; // @[Bitwise.scala 50:65:@5344.4]
  assign _T_5318 = _T_5303[14]; // @[Bitwise.scala 50:65:@5345.4]
  assign _T_5319 = _T_5303[15]; // @[Bitwise.scala 50:65:@5346.4]
  assign _T_5320 = _T_5303[16]; // @[Bitwise.scala 50:65:@5347.4]
  assign _T_5321 = _T_5303[17]; // @[Bitwise.scala 50:65:@5348.4]
  assign _T_5322 = _T_5303[18]; // @[Bitwise.scala 50:65:@5349.4]
  assign _T_5323 = _T_5303[19]; // @[Bitwise.scala 50:65:@5350.4]
  assign _T_5324 = _T_5303[20]; // @[Bitwise.scala 50:65:@5351.4]
  assign _T_5325 = _T_5303[21]; // @[Bitwise.scala 50:65:@5352.4]
  assign _T_5326 = _T_5303[22]; // @[Bitwise.scala 50:65:@5353.4]
  assign _T_5327 = _T_5303[23]; // @[Bitwise.scala 50:65:@5354.4]
  assign _T_5328 = _T_5303[24]; // @[Bitwise.scala 50:65:@5355.4]
  assign _T_5329 = _T_5303[25]; // @[Bitwise.scala 50:65:@5356.4]
  assign _T_5330 = _T_5303[26]; // @[Bitwise.scala 50:65:@5357.4]
  assign _T_5331 = _T_5303[27]; // @[Bitwise.scala 50:65:@5358.4]
  assign _T_5332 = _T_5303[28]; // @[Bitwise.scala 50:65:@5359.4]
  assign _T_5333 = _T_5303[29]; // @[Bitwise.scala 50:65:@5360.4]
  assign _T_5334 = _T_5303[30]; // @[Bitwise.scala 50:65:@5361.4]
  assign _T_5335 = _T_5303[31]; // @[Bitwise.scala 50:65:@5362.4]
  assign _T_5336 = _T_5303[32]; // @[Bitwise.scala 50:65:@5363.4]
  assign _T_5337 = _T_5304 + _T_5305; // @[Bitwise.scala 48:55:@5364.4]
  assign _T_5338 = _T_5306 + _T_5307; // @[Bitwise.scala 48:55:@5365.4]
  assign _T_5339 = _T_5337 + _T_5338; // @[Bitwise.scala 48:55:@5366.4]
  assign _T_5340 = _T_5308 + _T_5309; // @[Bitwise.scala 48:55:@5367.4]
  assign _T_5341 = _T_5310 + _T_5311; // @[Bitwise.scala 48:55:@5368.4]
  assign _T_5342 = _T_5340 + _T_5341; // @[Bitwise.scala 48:55:@5369.4]
  assign _T_5343 = _T_5339 + _T_5342; // @[Bitwise.scala 48:55:@5370.4]
  assign _T_5344 = _T_5312 + _T_5313; // @[Bitwise.scala 48:55:@5371.4]
  assign _T_5345 = _T_5314 + _T_5315; // @[Bitwise.scala 48:55:@5372.4]
  assign _T_5346 = _T_5344 + _T_5345; // @[Bitwise.scala 48:55:@5373.4]
  assign _T_5347 = _T_5316 + _T_5317; // @[Bitwise.scala 48:55:@5374.4]
  assign _T_5348 = _T_5318 + _T_5319; // @[Bitwise.scala 48:55:@5375.4]
  assign _T_5349 = _T_5347 + _T_5348; // @[Bitwise.scala 48:55:@5376.4]
  assign _T_5350 = _T_5346 + _T_5349; // @[Bitwise.scala 48:55:@5377.4]
  assign _T_5351 = _T_5343 + _T_5350; // @[Bitwise.scala 48:55:@5378.4]
  assign _T_5352 = _T_5320 + _T_5321; // @[Bitwise.scala 48:55:@5379.4]
  assign _T_5353 = _T_5322 + _T_5323; // @[Bitwise.scala 48:55:@5380.4]
  assign _T_5354 = _T_5352 + _T_5353; // @[Bitwise.scala 48:55:@5381.4]
  assign _T_5355 = _T_5324 + _T_5325; // @[Bitwise.scala 48:55:@5382.4]
  assign _T_5356 = _T_5326 + _T_5327; // @[Bitwise.scala 48:55:@5383.4]
  assign _T_5357 = _T_5355 + _T_5356; // @[Bitwise.scala 48:55:@5384.4]
  assign _T_5358 = _T_5354 + _T_5357; // @[Bitwise.scala 48:55:@5385.4]
  assign _T_5359 = _T_5328 + _T_5329; // @[Bitwise.scala 48:55:@5386.4]
  assign _T_5360 = _T_5330 + _T_5331; // @[Bitwise.scala 48:55:@5387.4]
  assign _T_5361 = _T_5359 + _T_5360; // @[Bitwise.scala 48:55:@5388.4]
  assign _T_5362 = _T_5332 + _T_5333; // @[Bitwise.scala 48:55:@5389.4]
  assign _T_5363 = _T_5335 + _T_5336; // @[Bitwise.scala 48:55:@5390.4]
  assign _GEN_656 = {{1'd0}, _T_5334}; // @[Bitwise.scala 48:55:@5391.4]
  assign _T_5364 = _GEN_656 + _T_5363; // @[Bitwise.scala 48:55:@5391.4]
  assign _GEN_657 = {{1'd0}, _T_5362}; // @[Bitwise.scala 48:55:@5392.4]
  assign _T_5365 = _GEN_657 + _T_5364; // @[Bitwise.scala 48:55:@5392.4]
  assign _GEN_658 = {{1'd0}, _T_5361}; // @[Bitwise.scala 48:55:@5393.4]
  assign _T_5366 = _GEN_658 + _T_5365; // @[Bitwise.scala 48:55:@5393.4]
  assign _GEN_659 = {{1'd0}, _T_5358}; // @[Bitwise.scala 48:55:@5394.4]
  assign _T_5367 = _GEN_659 + _T_5366; // @[Bitwise.scala 48:55:@5394.4]
  assign _GEN_660 = {{1'd0}, _T_5351}; // @[Bitwise.scala 48:55:@5395.4]
  assign _T_5368 = _GEN_660 + _T_5367; // @[Bitwise.scala 48:55:@5395.4]
  assign _T_5432 = _T_2230[33:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5460.4]
  assign _T_5433 = _T_5432[0]; // @[Bitwise.scala 50:65:@5461.4]
  assign _T_5434 = _T_5432[1]; // @[Bitwise.scala 50:65:@5462.4]
  assign _T_5435 = _T_5432[2]; // @[Bitwise.scala 50:65:@5463.4]
  assign _T_5436 = _T_5432[3]; // @[Bitwise.scala 50:65:@5464.4]
  assign _T_5437 = _T_5432[4]; // @[Bitwise.scala 50:65:@5465.4]
  assign _T_5438 = _T_5432[5]; // @[Bitwise.scala 50:65:@5466.4]
  assign _T_5439 = _T_5432[6]; // @[Bitwise.scala 50:65:@5467.4]
  assign _T_5440 = _T_5432[7]; // @[Bitwise.scala 50:65:@5468.4]
  assign _T_5441 = _T_5432[8]; // @[Bitwise.scala 50:65:@5469.4]
  assign _T_5442 = _T_5432[9]; // @[Bitwise.scala 50:65:@5470.4]
  assign _T_5443 = _T_5432[10]; // @[Bitwise.scala 50:65:@5471.4]
  assign _T_5444 = _T_5432[11]; // @[Bitwise.scala 50:65:@5472.4]
  assign _T_5445 = _T_5432[12]; // @[Bitwise.scala 50:65:@5473.4]
  assign _T_5446 = _T_5432[13]; // @[Bitwise.scala 50:65:@5474.4]
  assign _T_5447 = _T_5432[14]; // @[Bitwise.scala 50:65:@5475.4]
  assign _T_5448 = _T_5432[15]; // @[Bitwise.scala 50:65:@5476.4]
  assign _T_5449 = _T_5432[16]; // @[Bitwise.scala 50:65:@5477.4]
  assign _T_5450 = _T_5432[17]; // @[Bitwise.scala 50:65:@5478.4]
  assign _T_5451 = _T_5432[18]; // @[Bitwise.scala 50:65:@5479.4]
  assign _T_5452 = _T_5432[19]; // @[Bitwise.scala 50:65:@5480.4]
  assign _T_5453 = _T_5432[20]; // @[Bitwise.scala 50:65:@5481.4]
  assign _T_5454 = _T_5432[21]; // @[Bitwise.scala 50:65:@5482.4]
  assign _T_5455 = _T_5432[22]; // @[Bitwise.scala 50:65:@5483.4]
  assign _T_5456 = _T_5432[23]; // @[Bitwise.scala 50:65:@5484.4]
  assign _T_5457 = _T_5432[24]; // @[Bitwise.scala 50:65:@5485.4]
  assign _T_5458 = _T_5432[25]; // @[Bitwise.scala 50:65:@5486.4]
  assign _T_5459 = _T_5432[26]; // @[Bitwise.scala 50:65:@5487.4]
  assign _T_5460 = _T_5432[27]; // @[Bitwise.scala 50:65:@5488.4]
  assign _T_5461 = _T_5432[28]; // @[Bitwise.scala 50:65:@5489.4]
  assign _T_5462 = _T_5432[29]; // @[Bitwise.scala 50:65:@5490.4]
  assign _T_5463 = _T_5432[30]; // @[Bitwise.scala 50:65:@5491.4]
  assign _T_5464 = _T_5432[31]; // @[Bitwise.scala 50:65:@5492.4]
  assign _T_5465 = _T_5432[32]; // @[Bitwise.scala 50:65:@5493.4]
  assign _T_5466 = _T_5432[33]; // @[Bitwise.scala 50:65:@5494.4]
  assign _T_5467 = _T_5433 + _T_5434; // @[Bitwise.scala 48:55:@5495.4]
  assign _T_5468 = _T_5435 + _T_5436; // @[Bitwise.scala 48:55:@5496.4]
  assign _T_5469 = _T_5467 + _T_5468; // @[Bitwise.scala 48:55:@5497.4]
  assign _T_5470 = _T_5437 + _T_5438; // @[Bitwise.scala 48:55:@5498.4]
  assign _T_5471 = _T_5439 + _T_5440; // @[Bitwise.scala 48:55:@5499.4]
  assign _T_5472 = _T_5470 + _T_5471; // @[Bitwise.scala 48:55:@5500.4]
  assign _T_5473 = _T_5469 + _T_5472; // @[Bitwise.scala 48:55:@5501.4]
  assign _T_5474 = _T_5441 + _T_5442; // @[Bitwise.scala 48:55:@5502.4]
  assign _T_5475 = _T_5443 + _T_5444; // @[Bitwise.scala 48:55:@5503.4]
  assign _T_5476 = _T_5474 + _T_5475; // @[Bitwise.scala 48:55:@5504.4]
  assign _T_5477 = _T_5445 + _T_5446; // @[Bitwise.scala 48:55:@5505.4]
  assign _T_5478 = _T_5448 + _T_5449; // @[Bitwise.scala 48:55:@5506.4]
  assign _GEN_661 = {{1'd0}, _T_5447}; // @[Bitwise.scala 48:55:@5507.4]
  assign _T_5479 = _GEN_661 + _T_5478; // @[Bitwise.scala 48:55:@5507.4]
  assign _GEN_662 = {{1'd0}, _T_5477}; // @[Bitwise.scala 48:55:@5508.4]
  assign _T_5480 = _GEN_662 + _T_5479; // @[Bitwise.scala 48:55:@5508.4]
  assign _GEN_663 = {{1'd0}, _T_5476}; // @[Bitwise.scala 48:55:@5509.4]
  assign _T_5481 = _GEN_663 + _T_5480; // @[Bitwise.scala 48:55:@5509.4]
  assign _GEN_664 = {{1'd0}, _T_5473}; // @[Bitwise.scala 48:55:@5510.4]
  assign _T_5482 = _GEN_664 + _T_5481; // @[Bitwise.scala 48:55:@5510.4]
  assign _T_5483 = _T_5450 + _T_5451; // @[Bitwise.scala 48:55:@5511.4]
  assign _T_5484 = _T_5452 + _T_5453; // @[Bitwise.scala 48:55:@5512.4]
  assign _T_5485 = _T_5483 + _T_5484; // @[Bitwise.scala 48:55:@5513.4]
  assign _T_5486 = _T_5454 + _T_5455; // @[Bitwise.scala 48:55:@5514.4]
  assign _T_5487 = _T_5456 + _T_5457; // @[Bitwise.scala 48:55:@5515.4]
  assign _T_5488 = _T_5486 + _T_5487; // @[Bitwise.scala 48:55:@5516.4]
  assign _T_5489 = _T_5485 + _T_5488; // @[Bitwise.scala 48:55:@5517.4]
  assign _T_5490 = _T_5458 + _T_5459; // @[Bitwise.scala 48:55:@5518.4]
  assign _T_5491 = _T_5460 + _T_5461; // @[Bitwise.scala 48:55:@5519.4]
  assign _T_5492 = _T_5490 + _T_5491; // @[Bitwise.scala 48:55:@5520.4]
  assign _T_5493 = _T_5462 + _T_5463; // @[Bitwise.scala 48:55:@5521.4]
  assign _T_5494 = _T_5465 + _T_5466; // @[Bitwise.scala 48:55:@5522.4]
  assign _GEN_665 = {{1'd0}, _T_5464}; // @[Bitwise.scala 48:55:@5523.4]
  assign _T_5495 = _GEN_665 + _T_5494; // @[Bitwise.scala 48:55:@5523.4]
  assign _GEN_666 = {{1'd0}, _T_5493}; // @[Bitwise.scala 48:55:@5524.4]
  assign _T_5496 = _GEN_666 + _T_5495; // @[Bitwise.scala 48:55:@5524.4]
  assign _GEN_667 = {{1'd0}, _T_5492}; // @[Bitwise.scala 48:55:@5525.4]
  assign _T_5497 = _GEN_667 + _T_5496; // @[Bitwise.scala 48:55:@5525.4]
  assign _GEN_668 = {{1'd0}, _T_5489}; // @[Bitwise.scala 48:55:@5526.4]
  assign _T_5498 = _GEN_668 + _T_5497; // @[Bitwise.scala 48:55:@5526.4]
  assign _T_5499 = _T_5482 + _T_5498; // @[Bitwise.scala 48:55:@5527.4]
  assign _T_5563 = _T_2230[34:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5592.4]
  assign _T_5564 = _T_5563[0]; // @[Bitwise.scala 50:65:@5593.4]
  assign _T_5565 = _T_5563[1]; // @[Bitwise.scala 50:65:@5594.4]
  assign _T_5566 = _T_5563[2]; // @[Bitwise.scala 50:65:@5595.4]
  assign _T_5567 = _T_5563[3]; // @[Bitwise.scala 50:65:@5596.4]
  assign _T_5568 = _T_5563[4]; // @[Bitwise.scala 50:65:@5597.4]
  assign _T_5569 = _T_5563[5]; // @[Bitwise.scala 50:65:@5598.4]
  assign _T_5570 = _T_5563[6]; // @[Bitwise.scala 50:65:@5599.4]
  assign _T_5571 = _T_5563[7]; // @[Bitwise.scala 50:65:@5600.4]
  assign _T_5572 = _T_5563[8]; // @[Bitwise.scala 50:65:@5601.4]
  assign _T_5573 = _T_5563[9]; // @[Bitwise.scala 50:65:@5602.4]
  assign _T_5574 = _T_5563[10]; // @[Bitwise.scala 50:65:@5603.4]
  assign _T_5575 = _T_5563[11]; // @[Bitwise.scala 50:65:@5604.4]
  assign _T_5576 = _T_5563[12]; // @[Bitwise.scala 50:65:@5605.4]
  assign _T_5577 = _T_5563[13]; // @[Bitwise.scala 50:65:@5606.4]
  assign _T_5578 = _T_5563[14]; // @[Bitwise.scala 50:65:@5607.4]
  assign _T_5579 = _T_5563[15]; // @[Bitwise.scala 50:65:@5608.4]
  assign _T_5580 = _T_5563[16]; // @[Bitwise.scala 50:65:@5609.4]
  assign _T_5581 = _T_5563[17]; // @[Bitwise.scala 50:65:@5610.4]
  assign _T_5582 = _T_5563[18]; // @[Bitwise.scala 50:65:@5611.4]
  assign _T_5583 = _T_5563[19]; // @[Bitwise.scala 50:65:@5612.4]
  assign _T_5584 = _T_5563[20]; // @[Bitwise.scala 50:65:@5613.4]
  assign _T_5585 = _T_5563[21]; // @[Bitwise.scala 50:65:@5614.4]
  assign _T_5586 = _T_5563[22]; // @[Bitwise.scala 50:65:@5615.4]
  assign _T_5587 = _T_5563[23]; // @[Bitwise.scala 50:65:@5616.4]
  assign _T_5588 = _T_5563[24]; // @[Bitwise.scala 50:65:@5617.4]
  assign _T_5589 = _T_5563[25]; // @[Bitwise.scala 50:65:@5618.4]
  assign _T_5590 = _T_5563[26]; // @[Bitwise.scala 50:65:@5619.4]
  assign _T_5591 = _T_5563[27]; // @[Bitwise.scala 50:65:@5620.4]
  assign _T_5592 = _T_5563[28]; // @[Bitwise.scala 50:65:@5621.4]
  assign _T_5593 = _T_5563[29]; // @[Bitwise.scala 50:65:@5622.4]
  assign _T_5594 = _T_5563[30]; // @[Bitwise.scala 50:65:@5623.4]
  assign _T_5595 = _T_5563[31]; // @[Bitwise.scala 50:65:@5624.4]
  assign _T_5596 = _T_5563[32]; // @[Bitwise.scala 50:65:@5625.4]
  assign _T_5597 = _T_5563[33]; // @[Bitwise.scala 50:65:@5626.4]
  assign _T_5598 = _T_5563[34]; // @[Bitwise.scala 50:65:@5627.4]
  assign _T_5599 = _T_5564 + _T_5565; // @[Bitwise.scala 48:55:@5628.4]
  assign _T_5600 = _T_5566 + _T_5567; // @[Bitwise.scala 48:55:@5629.4]
  assign _T_5601 = _T_5599 + _T_5600; // @[Bitwise.scala 48:55:@5630.4]
  assign _T_5602 = _T_5568 + _T_5569; // @[Bitwise.scala 48:55:@5631.4]
  assign _T_5603 = _T_5570 + _T_5571; // @[Bitwise.scala 48:55:@5632.4]
  assign _T_5604 = _T_5602 + _T_5603; // @[Bitwise.scala 48:55:@5633.4]
  assign _T_5605 = _T_5601 + _T_5604; // @[Bitwise.scala 48:55:@5634.4]
  assign _T_5606 = _T_5572 + _T_5573; // @[Bitwise.scala 48:55:@5635.4]
  assign _T_5607 = _T_5574 + _T_5575; // @[Bitwise.scala 48:55:@5636.4]
  assign _T_5608 = _T_5606 + _T_5607; // @[Bitwise.scala 48:55:@5637.4]
  assign _T_5609 = _T_5576 + _T_5577; // @[Bitwise.scala 48:55:@5638.4]
  assign _T_5610 = _T_5579 + _T_5580; // @[Bitwise.scala 48:55:@5639.4]
  assign _GEN_669 = {{1'd0}, _T_5578}; // @[Bitwise.scala 48:55:@5640.4]
  assign _T_5611 = _GEN_669 + _T_5610; // @[Bitwise.scala 48:55:@5640.4]
  assign _GEN_670 = {{1'd0}, _T_5609}; // @[Bitwise.scala 48:55:@5641.4]
  assign _T_5612 = _GEN_670 + _T_5611; // @[Bitwise.scala 48:55:@5641.4]
  assign _GEN_671 = {{1'd0}, _T_5608}; // @[Bitwise.scala 48:55:@5642.4]
  assign _T_5613 = _GEN_671 + _T_5612; // @[Bitwise.scala 48:55:@5642.4]
  assign _GEN_672 = {{1'd0}, _T_5605}; // @[Bitwise.scala 48:55:@5643.4]
  assign _T_5614 = _GEN_672 + _T_5613; // @[Bitwise.scala 48:55:@5643.4]
  assign _T_5615 = _T_5581 + _T_5582; // @[Bitwise.scala 48:55:@5644.4]
  assign _T_5616 = _T_5583 + _T_5584; // @[Bitwise.scala 48:55:@5645.4]
  assign _T_5617 = _T_5615 + _T_5616; // @[Bitwise.scala 48:55:@5646.4]
  assign _T_5618 = _T_5585 + _T_5586; // @[Bitwise.scala 48:55:@5647.4]
  assign _T_5619 = _T_5588 + _T_5589; // @[Bitwise.scala 48:55:@5648.4]
  assign _GEN_673 = {{1'd0}, _T_5587}; // @[Bitwise.scala 48:55:@5649.4]
  assign _T_5620 = _GEN_673 + _T_5619; // @[Bitwise.scala 48:55:@5649.4]
  assign _GEN_674 = {{1'd0}, _T_5618}; // @[Bitwise.scala 48:55:@5650.4]
  assign _T_5621 = _GEN_674 + _T_5620; // @[Bitwise.scala 48:55:@5650.4]
  assign _GEN_675 = {{1'd0}, _T_5617}; // @[Bitwise.scala 48:55:@5651.4]
  assign _T_5622 = _GEN_675 + _T_5621; // @[Bitwise.scala 48:55:@5651.4]
  assign _T_5623 = _T_5590 + _T_5591; // @[Bitwise.scala 48:55:@5652.4]
  assign _T_5624 = _T_5592 + _T_5593; // @[Bitwise.scala 48:55:@5653.4]
  assign _T_5625 = _T_5623 + _T_5624; // @[Bitwise.scala 48:55:@5654.4]
  assign _T_5626 = _T_5594 + _T_5595; // @[Bitwise.scala 48:55:@5655.4]
  assign _T_5627 = _T_5597 + _T_5598; // @[Bitwise.scala 48:55:@5656.4]
  assign _GEN_676 = {{1'd0}, _T_5596}; // @[Bitwise.scala 48:55:@5657.4]
  assign _T_5628 = _GEN_676 + _T_5627; // @[Bitwise.scala 48:55:@5657.4]
  assign _GEN_677 = {{1'd0}, _T_5626}; // @[Bitwise.scala 48:55:@5658.4]
  assign _T_5629 = _GEN_677 + _T_5628; // @[Bitwise.scala 48:55:@5658.4]
  assign _GEN_678 = {{1'd0}, _T_5625}; // @[Bitwise.scala 48:55:@5659.4]
  assign _T_5630 = _GEN_678 + _T_5629; // @[Bitwise.scala 48:55:@5659.4]
  assign _T_5631 = _T_5622 + _T_5630; // @[Bitwise.scala 48:55:@5660.4]
  assign _T_5632 = _T_5614 + _T_5631; // @[Bitwise.scala 48:55:@5661.4]
  assign _T_5696 = _T_2230[35:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5726.4]
  assign _T_5697 = _T_5696[0]; // @[Bitwise.scala 50:65:@5727.4]
  assign _T_5698 = _T_5696[1]; // @[Bitwise.scala 50:65:@5728.4]
  assign _T_5699 = _T_5696[2]; // @[Bitwise.scala 50:65:@5729.4]
  assign _T_5700 = _T_5696[3]; // @[Bitwise.scala 50:65:@5730.4]
  assign _T_5701 = _T_5696[4]; // @[Bitwise.scala 50:65:@5731.4]
  assign _T_5702 = _T_5696[5]; // @[Bitwise.scala 50:65:@5732.4]
  assign _T_5703 = _T_5696[6]; // @[Bitwise.scala 50:65:@5733.4]
  assign _T_5704 = _T_5696[7]; // @[Bitwise.scala 50:65:@5734.4]
  assign _T_5705 = _T_5696[8]; // @[Bitwise.scala 50:65:@5735.4]
  assign _T_5706 = _T_5696[9]; // @[Bitwise.scala 50:65:@5736.4]
  assign _T_5707 = _T_5696[10]; // @[Bitwise.scala 50:65:@5737.4]
  assign _T_5708 = _T_5696[11]; // @[Bitwise.scala 50:65:@5738.4]
  assign _T_5709 = _T_5696[12]; // @[Bitwise.scala 50:65:@5739.4]
  assign _T_5710 = _T_5696[13]; // @[Bitwise.scala 50:65:@5740.4]
  assign _T_5711 = _T_5696[14]; // @[Bitwise.scala 50:65:@5741.4]
  assign _T_5712 = _T_5696[15]; // @[Bitwise.scala 50:65:@5742.4]
  assign _T_5713 = _T_5696[16]; // @[Bitwise.scala 50:65:@5743.4]
  assign _T_5714 = _T_5696[17]; // @[Bitwise.scala 50:65:@5744.4]
  assign _T_5715 = _T_5696[18]; // @[Bitwise.scala 50:65:@5745.4]
  assign _T_5716 = _T_5696[19]; // @[Bitwise.scala 50:65:@5746.4]
  assign _T_5717 = _T_5696[20]; // @[Bitwise.scala 50:65:@5747.4]
  assign _T_5718 = _T_5696[21]; // @[Bitwise.scala 50:65:@5748.4]
  assign _T_5719 = _T_5696[22]; // @[Bitwise.scala 50:65:@5749.4]
  assign _T_5720 = _T_5696[23]; // @[Bitwise.scala 50:65:@5750.4]
  assign _T_5721 = _T_5696[24]; // @[Bitwise.scala 50:65:@5751.4]
  assign _T_5722 = _T_5696[25]; // @[Bitwise.scala 50:65:@5752.4]
  assign _T_5723 = _T_5696[26]; // @[Bitwise.scala 50:65:@5753.4]
  assign _T_5724 = _T_5696[27]; // @[Bitwise.scala 50:65:@5754.4]
  assign _T_5725 = _T_5696[28]; // @[Bitwise.scala 50:65:@5755.4]
  assign _T_5726 = _T_5696[29]; // @[Bitwise.scala 50:65:@5756.4]
  assign _T_5727 = _T_5696[30]; // @[Bitwise.scala 50:65:@5757.4]
  assign _T_5728 = _T_5696[31]; // @[Bitwise.scala 50:65:@5758.4]
  assign _T_5729 = _T_5696[32]; // @[Bitwise.scala 50:65:@5759.4]
  assign _T_5730 = _T_5696[33]; // @[Bitwise.scala 50:65:@5760.4]
  assign _T_5731 = _T_5696[34]; // @[Bitwise.scala 50:65:@5761.4]
  assign _T_5732 = _T_5696[35]; // @[Bitwise.scala 50:65:@5762.4]
  assign _T_5733 = _T_5697 + _T_5698; // @[Bitwise.scala 48:55:@5763.4]
  assign _T_5734 = _T_5699 + _T_5700; // @[Bitwise.scala 48:55:@5764.4]
  assign _T_5735 = _T_5733 + _T_5734; // @[Bitwise.scala 48:55:@5765.4]
  assign _T_5736 = _T_5701 + _T_5702; // @[Bitwise.scala 48:55:@5766.4]
  assign _T_5737 = _T_5704 + _T_5705; // @[Bitwise.scala 48:55:@5767.4]
  assign _GEN_679 = {{1'd0}, _T_5703}; // @[Bitwise.scala 48:55:@5768.4]
  assign _T_5738 = _GEN_679 + _T_5737; // @[Bitwise.scala 48:55:@5768.4]
  assign _GEN_680 = {{1'd0}, _T_5736}; // @[Bitwise.scala 48:55:@5769.4]
  assign _T_5739 = _GEN_680 + _T_5738; // @[Bitwise.scala 48:55:@5769.4]
  assign _GEN_681 = {{1'd0}, _T_5735}; // @[Bitwise.scala 48:55:@5770.4]
  assign _T_5740 = _GEN_681 + _T_5739; // @[Bitwise.scala 48:55:@5770.4]
  assign _T_5741 = _T_5706 + _T_5707; // @[Bitwise.scala 48:55:@5771.4]
  assign _T_5742 = _T_5708 + _T_5709; // @[Bitwise.scala 48:55:@5772.4]
  assign _T_5743 = _T_5741 + _T_5742; // @[Bitwise.scala 48:55:@5773.4]
  assign _T_5744 = _T_5710 + _T_5711; // @[Bitwise.scala 48:55:@5774.4]
  assign _T_5745 = _T_5713 + _T_5714; // @[Bitwise.scala 48:55:@5775.4]
  assign _GEN_682 = {{1'd0}, _T_5712}; // @[Bitwise.scala 48:55:@5776.4]
  assign _T_5746 = _GEN_682 + _T_5745; // @[Bitwise.scala 48:55:@5776.4]
  assign _GEN_683 = {{1'd0}, _T_5744}; // @[Bitwise.scala 48:55:@5777.4]
  assign _T_5747 = _GEN_683 + _T_5746; // @[Bitwise.scala 48:55:@5777.4]
  assign _GEN_684 = {{1'd0}, _T_5743}; // @[Bitwise.scala 48:55:@5778.4]
  assign _T_5748 = _GEN_684 + _T_5747; // @[Bitwise.scala 48:55:@5778.4]
  assign _T_5749 = _T_5740 + _T_5748; // @[Bitwise.scala 48:55:@5779.4]
  assign _T_5750 = _T_5715 + _T_5716; // @[Bitwise.scala 48:55:@5780.4]
  assign _T_5751 = _T_5717 + _T_5718; // @[Bitwise.scala 48:55:@5781.4]
  assign _T_5752 = _T_5750 + _T_5751; // @[Bitwise.scala 48:55:@5782.4]
  assign _T_5753 = _T_5719 + _T_5720; // @[Bitwise.scala 48:55:@5783.4]
  assign _T_5754 = _T_5722 + _T_5723; // @[Bitwise.scala 48:55:@5784.4]
  assign _GEN_685 = {{1'd0}, _T_5721}; // @[Bitwise.scala 48:55:@5785.4]
  assign _T_5755 = _GEN_685 + _T_5754; // @[Bitwise.scala 48:55:@5785.4]
  assign _GEN_686 = {{1'd0}, _T_5753}; // @[Bitwise.scala 48:55:@5786.4]
  assign _T_5756 = _GEN_686 + _T_5755; // @[Bitwise.scala 48:55:@5786.4]
  assign _GEN_687 = {{1'd0}, _T_5752}; // @[Bitwise.scala 48:55:@5787.4]
  assign _T_5757 = _GEN_687 + _T_5756; // @[Bitwise.scala 48:55:@5787.4]
  assign _T_5758 = _T_5724 + _T_5725; // @[Bitwise.scala 48:55:@5788.4]
  assign _T_5759 = _T_5726 + _T_5727; // @[Bitwise.scala 48:55:@5789.4]
  assign _T_5760 = _T_5758 + _T_5759; // @[Bitwise.scala 48:55:@5790.4]
  assign _T_5761 = _T_5728 + _T_5729; // @[Bitwise.scala 48:55:@5791.4]
  assign _T_5762 = _T_5731 + _T_5732; // @[Bitwise.scala 48:55:@5792.4]
  assign _GEN_688 = {{1'd0}, _T_5730}; // @[Bitwise.scala 48:55:@5793.4]
  assign _T_5763 = _GEN_688 + _T_5762; // @[Bitwise.scala 48:55:@5793.4]
  assign _GEN_689 = {{1'd0}, _T_5761}; // @[Bitwise.scala 48:55:@5794.4]
  assign _T_5764 = _GEN_689 + _T_5763; // @[Bitwise.scala 48:55:@5794.4]
  assign _GEN_690 = {{1'd0}, _T_5760}; // @[Bitwise.scala 48:55:@5795.4]
  assign _T_5765 = _GEN_690 + _T_5764; // @[Bitwise.scala 48:55:@5795.4]
  assign _T_5766 = _T_5757 + _T_5765; // @[Bitwise.scala 48:55:@5796.4]
  assign _T_5767 = _T_5749 + _T_5766; // @[Bitwise.scala 48:55:@5797.4]
  assign _T_5831 = _T_2230[36:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5862.4]
  assign _T_5832 = _T_5831[0]; // @[Bitwise.scala 50:65:@5863.4]
  assign _T_5833 = _T_5831[1]; // @[Bitwise.scala 50:65:@5864.4]
  assign _T_5834 = _T_5831[2]; // @[Bitwise.scala 50:65:@5865.4]
  assign _T_5835 = _T_5831[3]; // @[Bitwise.scala 50:65:@5866.4]
  assign _T_5836 = _T_5831[4]; // @[Bitwise.scala 50:65:@5867.4]
  assign _T_5837 = _T_5831[5]; // @[Bitwise.scala 50:65:@5868.4]
  assign _T_5838 = _T_5831[6]; // @[Bitwise.scala 50:65:@5869.4]
  assign _T_5839 = _T_5831[7]; // @[Bitwise.scala 50:65:@5870.4]
  assign _T_5840 = _T_5831[8]; // @[Bitwise.scala 50:65:@5871.4]
  assign _T_5841 = _T_5831[9]; // @[Bitwise.scala 50:65:@5872.4]
  assign _T_5842 = _T_5831[10]; // @[Bitwise.scala 50:65:@5873.4]
  assign _T_5843 = _T_5831[11]; // @[Bitwise.scala 50:65:@5874.4]
  assign _T_5844 = _T_5831[12]; // @[Bitwise.scala 50:65:@5875.4]
  assign _T_5845 = _T_5831[13]; // @[Bitwise.scala 50:65:@5876.4]
  assign _T_5846 = _T_5831[14]; // @[Bitwise.scala 50:65:@5877.4]
  assign _T_5847 = _T_5831[15]; // @[Bitwise.scala 50:65:@5878.4]
  assign _T_5848 = _T_5831[16]; // @[Bitwise.scala 50:65:@5879.4]
  assign _T_5849 = _T_5831[17]; // @[Bitwise.scala 50:65:@5880.4]
  assign _T_5850 = _T_5831[18]; // @[Bitwise.scala 50:65:@5881.4]
  assign _T_5851 = _T_5831[19]; // @[Bitwise.scala 50:65:@5882.4]
  assign _T_5852 = _T_5831[20]; // @[Bitwise.scala 50:65:@5883.4]
  assign _T_5853 = _T_5831[21]; // @[Bitwise.scala 50:65:@5884.4]
  assign _T_5854 = _T_5831[22]; // @[Bitwise.scala 50:65:@5885.4]
  assign _T_5855 = _T_5831[23]; // @[Bitwise.scala 50:65:@5886.4]
  assign _T_5856 = _T_5831[24]; // @[Bitwise.scala 50:65:@5887.4]
  assign _T_5857 = _T_5831[25]; // @[Bitwise.scala 50:65:@5888.4]
  assign _T_5858 = _T_5831[26]; // @[Bitwise.scala 50:65:@5889.4]
  assign _T_5859 = _T_5831[27]; // @[Bitwise.scala 50:65:@5890.4]
  assign _T_5860 = _T_5831[28]; // @[Bitwise.scala 50:65:@5891.4]
  assign _T_5861 = _T_5831[29]; // @[Bitwise.scala 50:65:@5892.4]
  assign _T_5862 = _T_5831[30]; // @[Bitwise.scala 50:65:@5893.4]
  assign _T_5863 = _T_5831[31]; // @[Bitwise.scala 50:65:@5894.4]
  assign _T_5864 = _T_5831[32]; // @[Bitwise.scala 50:65:@5895.4]
  assign _T_5865 = _T_5831[33]; // @[Bitwise.scala 50:65:@5896.4]
  assign _T_5866 = _T_5831[34]; // @[Bitwise.scala 50:65:@5897.4]
  assign _T_5867 = _T_5831[35]; // @[Bitwise.scala 50:65:@5898.4]
  assign _T_5868 = _T_5831[36]; // @[Bitwise.scala 50:65:@5899.4]
  assign _T_5869 = _T_5832 + _T_5833; // @[Bitwise.scala 48:55:@5900.4]
  assign _T_5870 = _T_5834 + _T_5835; // @[Bitwise.scala 48:55:@5901.4]
  assign _T_5871 = _T_5869 + _T_5870; // @[Bitwise.scala 48:55:@5902.4]
  assign _T_5872 = _T_5836 + _T_5837; // @[Bitwise.scala 48:55:@5903.4]
  assign _T_5873 = _T_5839 + _T_5840; // @[Bitwise.scala 48:55:@5904.4]
  assign _GEN_691 = {{1'd0}, _T_5838}; // @[Bitwise.scala 48:55:@5905.4]
  assign _T_5874 = _GEN_691 + _T_5873; // @[Bitwise.scala 48:55:@5905.4]
  assign _GEN_692 = {{1'd0}, _T_5872}; // @[Bitwise.scala 48:55:@5906.4]
  assign _T_5875 = _GEN_692 + _T_5874; // @[Bitwise.scala 48:55:@5906.4]
  assign _GEN_693 = {{1'd0}, _T_5871}; // @[Bitwise.scala 48:55:@5907.4]
  assign _T_5876 = _GEN_693 + _T_5875; // @[Bitwise.scala 48:55:@5907.4]
  assign _T_5877 = _T_5841 + _T_5842; // @[Bitwise.scala 48:55:@5908.4]
  assign _T_5878 = _T_5843 + _T_5844; // @[Bitwise.scala 48:55:@5909.4]
  assign _T_5879 = _T_5877 + _T_5878; // @[Bitwise.scala 48:55:@5910.4]
  assign _T_5880 = _T_5845 + _T_5846; // @[Bitwise.scala 48:55:@5911.4]
  assign _T_5881 = _T_5848 + _T_5849; // @[Bitwise.scala 48:55:@5912.4]
  assign _GEN_694 = {{1'd0}, _T_5847}; // @[Bitwise.scala 48:55:@5913.4]
  assign _T_5882 = _GEN_694 + _T_5881; // @[Bitwise.scala 48:55:@5913.4]
  assign _GEN_695 = {{1'd0}, _T_5880}; // @[Bitwise.scala 48:55:@5914.4]
  assign _T_5883 = _GEN_695 + _T_5882; // @[Bitwise.scala 48:55:@5914.4]
  assign _GEN_696 = {{1'd0}, _T_5879}; // @[Bitwise.scala 48:55:@5915.4]
  assign _T_5884 = _GEN_696 + _T_5883; // @[Bitwise.scala 48:55:@5915.4]
  assign _T_5885 = _T_5876 + _T_5884; // @[Bitwise.scala 48:55:@5916.4]
  assign _T_5886 = _T_5850 + _T_5851; // @[Bitwise.scala 48:55:@5917.4]
  assign _T_5887 = _T_5852 + _T_5853; // @[Bitwise.scala 48:55:@5918.4]
  assign _T_5888 = _T_5886 + _T_5887; // @[Bitwise.scala 48:55:@5919.4]
  assign _T_5889 = _T_5854 + _T_5855; // @[Bitwise.scala 48:55:@5920.4]
  assign _T_5890 = _T_5857 + _T_5858; // @[Bitwise.scala 48:55:@5921.4]
  assign _GEN_697 = {{1'd0}, _T_5856}; // @[Bitwise.scala 48:55:@5922.4]
  assign _T_5891 = _GEN_697 + _T_5890; // @[Bitwise.scala 48:55:@5922.4]
  assign _GEN_698 = {{1'd0}, _T_5889}; // @[Bitwise.scala 48:55:@5923.4]
  assign _T_5892 = _GEN_698 + _T_5891; // @[Bitwise.scala 48:55:@5923.4]
  assign _GEN_699 = {{1'd0}, _T_5888}; // @[Bitwise.scala 48:55:@5924.4]
  assign _T_5893 = _GEN_699 + _T_5892; // @[Bitwise.scala 48:55:@5924.4]
  assign _T_5894 = _T_5859 + _T_5860; // @[Bitwise.scala 48:55:@5925.4]
  assign _T_5895 = _T_5862 + _T_5863; // @[Bitwise.scala 48:55:@5926.4]
  assign _GEN_700 = {{1'd0}, _T_5861}; // @[Bitwise.scala 48:55:@5927.4]
  assign _T_5896 = _GEN_700 + _T_5895; // @[Bitwise.scala 48:55:@5927.4]
  assign _GEN_701 = {{1'd0}, _T_5894}; // @[Bitwise.scala 48:55:@5928.4]
  assign _T_5897 = _GEN_701 + _T_5896; // @[Bitwise.scala 48:55:@5928.4]
  assign _T_5898 = _T_5864 + _T_5865; // @[Bitwise.scala 48:55:@5929.4]
  assign _T_5899 = _T_5867 + _T_5868; // @[Bitwise.scala 48:55:@5930.4]
  assign _GEN_702 = {{1'd0}, _T_5866}; // @[Bitwise.scala 48:55:@5931.4]
  assign _T_5900 = _GEN_702 + _T_5899; // @[Bitwise.scala 48:55:@5931.4]
  assign _GEN_703 = {{1'd0}, _T_5898}; // @[Bitwise.scala 48:55:@5932.4]
  assign _T_5901 = _GEN_703 + _T_5900; // @[Bitwise.scala 48:55:@5932.4]
  assign _T_5902 = _T_5897 + _T_5901; // @[Bitwise.scala 48:55:@5933.4]
  assign _T_5903 = _T_5893 + _T_5902; // @[Bitwise.scala 48:55:@5934.4]
  assign _T_5904 = _T_5885 + _T_5903; // @[Bitwise.scala 48:55:@5935.4]
  assign _T_5968 = _T_2230[37:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6000.4]
  assign _T_5969 = _T_5968[0]; // @[Bitwise.scala 50:65:@6001.4]
  assign _T_5970 = _T_5968[1]; // @[Bitwise.scala 50:65:@6002.4]
  assign _T_5971 = _T_5968[2]; // @[Bitwise.scala 50:65:@6003.4]
  assign _T_5972 = _T_5968[3]; // @[Bitwise.scala 50:65:@6004.4]
  assign _T_5973 = _T_5968[4]; // @[Bitwise.scala 50:65:@6005.4]
  assign _T_5974 = _T_5968[5]; // @[Bitwise.scala 50:65:@6006.4]
  assign _T_5975 = _T_5968[6]; // @[Bitwise.scala 50:65:@6007.4]
  assign _T_5976 = _T_5968[7]; // @[Bitwise.scala 50:65:@6008.4]
  assign _T_5977 = _T_5968[8]; // @[Bitwise.scala 50:65:@6009.4]
  assign _T_5978 = _T_5968[9]; // @[Bitwise.scala 50:65:@6010.4]
  assign _T_5979 = _T_5968[10]; // @[Bitwise.scala 50:65:@6011.4]
  assign _T_5980 = _T_5968[11]; // @[Bitwise.scala 50:65:@6012.4]
  assign _T_5981 = _T_5968[12]; // @[Bitwise.scala 50:65:@6013.4]
  assign _T_5982 = _T_5968[13]; // @[Bitwise.scala 50:65:@6014.4]
  assign _T_5983 = _T_5968[14]; // @[Bitwise.scala 50:65:@6015.4]
  assign _T_5984 = _T_5968[15]; // @[Bitwise.scala 50:65:@6016.4]
  assign _T_5985 = _T_5968[16]; // @[Bitwise.scala 50:65:@6017.4]
  assign _T_5986 = _T_5968[17]; // @[Bitwise.scala 50:65:@6018.4]
  assign _T_5987 = _T_5968[18]; // @[Bitwise.scala 50:65:@6019.4]
  assign _T_5988 = _T_5968[19]; // @[Bitwise.scala 50:65:@6020.4]
  assign _T_5989 = _T_5968[20]; // @[Bitwise.scala 50:65:@6021.4]
  assign _T_5990 = _T_5968[21]; // @[Bitwise.scala 50:65:@6022.4]
  assign _T_5991 = _T_5968[22]; // @[Bitwise.scala 50:65:@6023.4]
  assign _T_5992 = _T_5968[23]; // @[Bitwise.scala 50:65:@6024.4]
  assign _T_5993 = _T_5968[24]; // @[Bitwise.scala 50:65:@6025.4]
  assign _T_5994 = _T_5968[25]; // @[Bitwise.scala 50:65:@6026.4]
  assign _T_5995 = _T_5968[26]; // @[Bitwise.scala 50:65:@6027.4]
  assign _T_5996 = _T_5968[27]; // @[Bitwise.scala 50:65:@6028.4]
  assign _T_5997 = _T_5968[28]; // @[Bitwise.scala 50:65:@6029.4]
  assign _T_5998 = _T_5968[29]; // @[Bitwise.scala 50:65:@6030.4]
  assign _T_5999 = _T_5968[30]; // @[Bitwise.scala 50:65:@6031.4]
  assign _T_6000 = _T_5968[31]; // @[Bitwise.scala 50:65:@6032.4]
  assign _T_6001 = _T_5968[32]; // @[Bitwise.scala 50:65:@6033.4]
  assign _T_6002 = _T_5968[33]; // @[Bitwise.scala 50:65:@6034.4]
  assign _T_6003 = _T_5968[34]; // @[Bitwise.scala 50:65:@6035.4]
  assign _T_6004 = _T_5968[35]; // @[Bitwise.scala 50:65:@6036.4]
  assign _T_6005 = _T_5968[36]; // @[Bitwise.scala 50:65:@6037.4]
  assign _T_6006 = _T_5968[37]; // @[Bitwise.scala 50:65:@6038.4]
  assign _T_6007 = _T_5969 + _T_5970; // @[Bitwise.scala 48:55:@6039.4]
  assign _T_6008 = _T_5971 + _T_5972; // @[Bitwise.scala 48:55:@6040.4]
  assign _T_6009 = _T_6007 + _T_6008; // @[Bitwise.scala 48:55:@6041.4]
  assign _T_6010 = _T_5973 + _T_5974; // @[Bitwise.scala 48:55:@6042.4]
  assign _T_6011 = _T_5976 + _T_5977; // @[Bitwise.scala 48:55:@6043.4]
  assign _GEN_704 = {{1'd0}, _T_5975}; // @[Bitwise.scala 48:55:@6044.4]
  assign _T_6012 = _GEN_704 + _T_6011; // @[Bitwise.scala 48:55:@6044.4]
  assign _GEN_705 = {{1'd0}, _T_6010}; // @[Bitwise.scala 48:55:@6045.4]
  assign _T_6013 = _GEN_705 + _T_6012; // @[Bitwise.scala 48:55:@6045.4]
  assign _GEN_706 = {{1'd0}, _T_6009}; // @[Bitwise.scala 48:55:@6046.4]
  assign _T_6014 = _GEN_706 + _T_6013; // @[Bitwise.scala 48:55:@6046.4]
  assign _T_6015 = _T_5978 + _T_5979; // @[Bitwise.scala 48:55:@6047.4]
  assign _T_6016 = _T_5981 + _T_5982; // @[Bitwise.scala 48:55:@6048.4]
  assign _GEN_707 = {{1'd0}, _T_5980}; // @[Bitwise.scala 48:55:@6049.4]
  assign _T_6017 = _GEN_707 + _T_6016; // @[Bitwise.scala 48:55:@6049.4]
  assign _GEN_708 = {{1'd0}, _T_6015}; // @[Bitwise.scala 48:55:@6050.4]
  assign _T_6018 = _GEN_708 + _T_6017; // @[Bitwise.scala 48:55:@6050.4]
  assign _T_6019 = _T_5983 + _T_5984; // @[Bitwise.scala 48:55:@6051.4]
  assign _T_6020 = _T_5986 + _T_5987; // @[Bitwise.scala 48:55:@6052.4]
  assign _GEN_709 = {{1'd0}, _T_5985}; // @[Bitwise.scala 48:55:@6053.4]
  assign _T_6021 = _GEN_709 + _T_6020; // @[Bitwise.scala 48:55:@6053.4]
  assign _GEN_710 = {{1'd0}, _T_6019}; // @[Bitwise.scala 48:55:@6054.4]
  assign _T_6022 = _GEN_710 + _T_6021; // @[Bitwise.scala 48:55:@6054.4]
  assign _T_6023 = _T_6018 + _T_6022; // @[Bitwise.scala 48:55:@6055.4]
  assign _T_6024 = _T_6014 + _T_6023; // @[Bitwise.scala 48:55:@6056.4]
  assign _T_6025 = _T_5988 + _T_5989; // @[Bitwise.scala 48:55:@6057.4]
  assign _T_6026 = _T_5990 + _T_5991; // @[Bitwise.scala 48:55:@6058.4]
  assign _T_6027 = _T_6025 + _T_6026; // @[Bitwise.scala 48:55:@6059.4]
  assign _T_6028 = _T_5992 + _T_5993; // @[Bitwise.scala 48:55:@6060.4]
  assign _T_6029 = _T_5995 + _T_5996; // @[Bitwise.scala 48:55:@6061.4]
  assign _GEN_711 = {{1'd0}, _T_5994}; // @[Bitwise.scala 48:55:@6062.4]
  assign _T_6030 = _GEN_711 + _T_6029; // @[Bitwise.scala 48:55:@6062.4]
  assign _GEN_712 = {{1'd0}, _T_6028}; // @[Bitwise.scala 48:55:@6063.4]
  assign _T_6031 = _GEN_712 + _T_6030; // @[Bitwise.scala 48:55:@6063.4]
  assign _GEN_713 = {{1'd0}, _T_6027}; // @[Bitwise.scala 48:55:@6064.4]
  assign _T_6032 = _GEN_713 + _T_6031; // @[Bitwise.scala 48:55:@6064.4]
  assign _T_6033 = _T_5997 + _T_5998; // @[Bitwise.scala 48:55:@6065.4]
  assign _T_6034 = _T_6000 + _T_6001; // @[Bitwise.scala 48:55:@6066.4]
  assign _GEN_714 = {{1'd0}, _T_5999}; // @[Bitwise.scala 48:55:@6067.4]
  assign _T_6035 = _GEN_714 + _T_6034; // @[Bitwise.scala 48:55:@6067.4]
  assign _GEN_715 = {{1'd0}, _T_6033}; // @[Bitwise.scala 48:55:@6068.4]
  assign _T_6036 = _GEN_715 + _T_6035; // @[Bitwise.scala 48:55:@6068.4]
  assign _T_6037 = _T_6002 + _T_6003; // @[Bitwise.scala 48:55:@6069.4]
  assign _T_6038 = _T_6005 + _T_6006; // @[Bitwise.scala 48:55:@6070.4]
  assign _GEN_716 = {{1'd0}, _T_6004}; // @[Bitwise.scala 48:55:@6071.4]
  assign _T_6039 = _GEN_716 + _T_6038; // @[Bitwise.scala 48:55:@6071.4]
  assign _GEN_717 = {{1'd0}, _T_6037}; // @[Bitwise.scala 48:55:@6072.4]
  assign _T_6040 = _GEN_717 + _T_6039; // @[Bitwise.scala 48:55:@6072.4]
  assign _T_6041 = _T_6036 + _T_6040; // @[Bitwise.scala 48:55:@6073.4]
  assign _T_6042 = _T_6032 + _T_6041; // @[Bitwise.scala 48:55:@6074.4]
  assign _T_6043 = _T_6024 + _T_6042; // @[Bitwise.scala 48:55:@6075.4]
  assign _T_6107 = _T_2230[38:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6140.4]
  assign _T_6108 = _T_6107[0]; // @[Bitwise.scala 50:65:@6141.4]
  assign _T_6109 = _T_6107[1]; // @[Bitwise.scala 50:65:@6142.4]
  assign _T_6110 = _T_6107[2]; // @[Bitwise.scala 50:65:@6143.4]
  assign _T_6111 = _T_6107[3]; // @[Bitwise.scala 50:65:@6144.4]
  assign _T_6112 = _T_6107[4]; // @[Bitwise.scala 50:65:@6145.4]
  assign _T_6113 = _T_6107[5]; // @[Bitwise.scala 50:65:@6146.4]
  assign _T_6114 = _T_6107[6]; // @[Bitwise.scala 50:65:@6147.4]
  assign _T_6115 = _T_6107[7]; // @[Bitwise.scala 50:65:@6148.4]
  assign _T_6116 = _T_6107[8]; // @[Bitwise.scala 50:65:@6149.4]
  assign _T_6117 = _T_6107[9]; // @[Bitwise.scala 50:65:@6150.4]
  assign _T_6118 = _T_6107[10]; // @[Bitwise.scala 50:65:@6151.4]
  assign _T_6119 = _T_6107[11]; // @[Bitwise.scala 50:65:@6152.4]
  assign _T_6120 = _T_6107[12]; // @[Bitwise.scala 50:65:@6153.4]
  assign _T_6121 = _T_6107[13]; // @[Bitwise.scala 50:65:@6154.4]
  assign _T_6122 = _T_6107[14]; // @[Bitwise.scala 50:65:@6155.4]
  assign _T_6123 = _T_6107[15]; // @[Bitwise.scala 50:65:@6156.4]
  assign _T_6124 = _T_6107[16]; // @[Bitwise.scala 50:65:@6157.4]
  assign _T_6125 = _T_6107[17]; // @[Bitwise.scala 50:65:@6158.4]
  assign _T_6126 = _T_6107[18]; // @[Bitwise.scala 50:65:@6159.4]
  assign _T_6127 = _T_6107[19]; // @[Bitwise.scala 50:65:@6160.4]
  assign _T_6128 = _T_6107[20]; // @[Bitwise.scala 50:65:@6161.4]
  assign _T_6129 = _T_6107[21]; // @[Bitwise.scala 50:65:@6162.4]
  assign _T_6130 = _T_6107[22]; // @[Bitwise.scala 50:65:@6163.4]
  assign _T_6131 = _T_6107[23]; // @[Bitwise.scala 50:65:@6164.4]
  assign _T_6132 = _T_6107[24]; // @[Bitwise.scala 50:65:@6165.4]
  assign _T_6133 = _T_6107[25]; // @[Bitwise.scala 50:65:@6166.4]
  assign _T_6134 = _T_6107[26]; // @[Bitwise.scala 50:65:@6167.4]
  assign _T_6135 = _T_6107[27]; // @[Bitwise.scala 50:65:@6168.4]
  assign _T_6136 = _T_6107[28]; // @[Bitwise.scala 50:65:@6169.4]
  assign _T_6137 = _T_6107[29]; // @[Bitwise.scala 50:65:@6170.4]
  assign _T_6138 = _T_6107[30]; // @[Bitwise.scala 50:65:@6171.4]
  assign _T_6139 = _T_6107[31]; // @[Bitwise.scala 50:65:@6172.4]
  assign _T_6140 = _T_6107[32]; // @[Bitwise.scala 50:65:@6173.4]
  assign _T_6141 = _T_6107[33]; // @[Bitwise.scala 50:65:@6174.4]
  assign _T_6142 = _T_6107[34]; // @[Bitwise.scala 50:65:@6175.4]
  assign _T_6143 = _T_6107[35]; // @[Bitwise.scala 50:65:@6176.4]
  assign _T_6144 = _T_6107[36]; // @[Bitwise.scala 50:65:@6177.4]
  assign _T_6145 = _T_6107[37]; // @[Bitwise.scala 50:65:@6178.4]
  assign _T_6146 = _T_6107[38]; // @[Bitwise.scala 50:65:@6179.4]
  assign _T_6147 = _T_6108 + _T_6109; // @[Bitwise.scala 48:55:@6180.4]
  assign _T_6148 = _T_6110 + _T_6111; // @[Bitwise.scala 48:55:@6181.4]
  assign _T_6149 = _T_6147 + _T_6148; // @[Bitwise.scala 48:55:@6182.4]
  assign _T_6150 = _T_6112 + _T_6113; // @[Bitwise.scala 48:55:@6183.4]
  assign _T_6151 = _T_6115 + _T_6116; // @[Bitwise.scala 48:55:@6184.4]
  assign _GEN_718 = {{1'd0}, _T_6114}; // @[Bitwise.scala 48:55:@6185.4]
  assign _T_6152 = _GEN_718 + _T_6151; // @[Bitwise.scala 48:55:@6185.4]
  assign _GEN_719 = {{1'd0}, _T_6150}; // @[Bitwise.scala 48:55:@6186.4]
  assign _T_6153 = _GEN_719 + _T_6152; // @[Bitwise.scala 48:55:@6186.4]
  assign _GEN_720 = {{1'd0}, _T_6149}; // @[Bitwise.scala 48:55:@6187.4]
  assign _T_6154 = _GEN_720 + _T_6153; // @[Bitwise.scala 48:55:@6187.4]
  assign _T_6155 = _T_6117 + _T_6118; // @[Bitwise.scala 48:55:@6188.4]
  assign _T_6156 = _T_6120 + _T_6121; // @[Bitwise.scala 48:55:@6189.4]
  assign _GEN_721 = {{1'd0}, _T_6119}; // @[Bitwise.scala 48:55:@6190.4]
  assign _T_6157 = _GEN_721 + _T_6156; // @[Bitwise.scala 48:55:@6190.4]
  assign _GEN_722 = {{1'd0}, _T_6155}; // @[Bitwise.scala 48:55:@6191.4]
  assign _T_6158 = _GEN_722 + _T_6157; // @[Bitwise.scala 48:55:@6191.4]
  assign _T_6159 = _T_6122 + _T_6123; // @[Bitwise.scala 48:55:@6192.4]
  assign _T_6160 = _T_6125 + _T_6126; // @[Bitwise.scala 48:55:@6193.4]
  assign _GEN_723 = {{1'd0}, _T_6124}; // @[Bitwise.scala 48:55:@6194.4]
  assign _T_6161 = _GEN_723 + _T_6160; // @[Bitwise.scala 48:55:@6194.4]
  assign _GEN_724 = {{1'd0}, _T_6159}; // @[Bitwise.scala 48:55:@6195.4]
  assign _T_6162 = _GEN_724 + _T_6161; // @[Bitwise.scala 48:55:@6195.4]
  assign _T_6163 = _T_6158 + _T_6162; // @[Bitwise.scala 48:55:@6196.4]
  assign _T_6164 = _T_6154 + _T_6163; // @[Bitwise.scala 48:55:@6197.4]
  assign _T_6165 = _T_6127 + _T_6128; // @[Bitwise.scala 48:55:@6198.4]
  assign _T_6166 = _T_6130 + _T_6131; // @[Bitwise.scala 48:55:@6199.4]
  assign _GEN_725 = {{1'd0}, _T_6129}; // @[Bitwise.scala 48:55:@6200.4]
  assign _T_6167 = _GEN_725 + _T_6166; // @[Bitwise.scala 48:55:@6200.4]
  assign _GEN_726 = {{1'd0}, _T_6165}; // @[Bitwise.scala 48:55:@6201.4]
  assign _T_6168 = _GEN_726 + _T_6167; // @[Bitwise.scala 48:55:@6201.4]
  assign _T_6169 = _T_6132 + _T_6133; // @[Bitwise.scala 48:55:@6202.4]
  assign _T_6170 = _T_6135 + _T_6136; // @[Bitwise.scala 48:55:@6203.4]
  assign _GEN_727 = {{1'd0}, _T_6134}; // @[Bitwise.scala 48:55:@6204.4]
  assign _T_6171 = _GEN_727 + _T_6170; // @[Bitwise.scala 48:55:@6204.4]
  assign _GEN_728 = {{1'd0}, _T_6169}; // @[Bitwise.scala 48:55:@6205.4]
  assign _T_6172 = _GEN_728 + _T_6171; // @[Bitwise.scala 48:55:@6205.4]
  assign _T_6173 = _T_6168 + _T_6172; // @[Bitwise.scala 48:55:@6206.4]
  assign _T_6174 = _T_6137 + _T_6138; // @[Bitwise.scala 48:55:@6207.4]
  assign _T_6175 = _T_6140 + _T_6141; // @[Bitwise.scala 48:55:@6208.4]
  assign _GEN_729 = {{1'd0}, _T_6139}; // @[Bitwise.scala 48:55:@6209.4]
  assign _T_6176 = _GEN_729 + _T_6175; // @[Bitwise.scala 48:55:@6209.4]
  assign _GEN_730 = {{1'd0}, _T_6174}; // @[Bitwise.scala 48:55:@6210.4]
  assign _T_6177 = _GEN_730 + _T_6176; // @[Bitwise.scala 48:55:@6210.4]
  assign _T_6178 = _T_6142 + _T_6143; // @[Bitwise.scala 48:55:@6211.4]
  assign _T_6179 = _T_6145 + _T_6146; // @[Bitwise.scala 48:55:@6212.4]
  assign _GEN_731 = {{1'd0}, _T_6144}; // @[Bitwise.scala 48:55:@6213.4]
  assign _T_6180 = _GEN_731 + _T_6179; // @[Bitwise.scala 48:55:@6213.4]
  assign _GEN_732 = {{1'd0}, _T_6178}; // @[Bitwise.scala 48:55:@6214.4]
  assign _T_6181 = _GEN_732 + _T_6180; // @[Bitwise.scala 48:55:@6214.4]
  assign _T_6182 = _T_6177 + _T_6181; // @[Bitwise.scala 48:55:@6215.4]
  assign _T_6183 = _T_6173 + _T_6182; // @[Bitwise.scala 48:55:@6216.4]
  assign _T_6184 = _T_6164 + _T_6183; // @[Bitwise.scala 48:55:@6217.4]
  assign _T_6248 = _T_2230[39:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6282.4]
  assign _T_6249 = _T_6248[0]; // @[Bitwise.scala 50:65:@6283.4]
  assign _T_6250 = _T_6248[1]; // @[Bitwise.scala 50:65:@6284.4]
  assign _T_6251 = _T_6248[2]; // @[Bitwise.scala 50:65:@6285.4]
  assign _T_6252 = _T_6248[3]; // @[Bitwise.scala 50:65:@6286.4]
  assign _T_6253 = _T_6248[4]; // @[Bitwise.scala 50:65:@6287.4]
  assign _T_6254 = _T_6248[5]; // @[Bitwise.scala 50:65:@6288.4]
  assign _T_6255 = _T_6248[6]; // @[Bitwise.scala 50:65:@6289.4]
  assign _T_6256 = _T_6248[7]; // @[Bitwise.scala 50:65:@6290.4]
  assign _T_6257 = _T_6248[8]; // @[Bitwise.scala 50:65:@6291.4]
  assign _T_6258 = _T_6248[9]; // @[Bitwise.scala 50:65:@6292.4]
  assign _T_6259 = _T_6248[10]; // @[Bitwise.scala 50:65:@6293.4]
  assign _T_6260 = _T_6248[11]; // @[Bitwise.scala 50:65:@6294.4]
  assign _T_6261 = _T_6248[12]; // @[Bitwise.scala 50:65:@6295.4]
  assign _T_6262 = _T_6248[13]; // @[Bitwise.scala 50:65:@6296.4]
  assign _T_6263 = _T_6248[14]; // @[Bitwise.scala 50:65:@6297.4]
  assign _T_6264 = _T_6248[15]; // @[Bitwise.scala 50:65:@6298.4]
  assign _T_6265 = _T_6248[16]; // @[Bitwise.scala 50:65:@6299.4]
  assign _T_6266 = _T_6248[17]; // @[Bitwise.scala 50:65:@6300.4]
  assign _T_6267 = _T_6248[18]; // @[Bitwise.scala 50:65:@6301.4]
  assign _T_6268 = _T_6248[19]; // @[Bitwise.scala 50:65:@6302.4]
  assign _T_6269 = _T_6248[20]; // @[Bitwise.scala 50:65:@6303.4]
  assign _T_6270 = _T_6248[21]; // @[Bitwise.scala 50:65:@6304.4]
  assign _T_6271 = _T_6248[22]; // @[Bitwise.scala 50:65:@6305.4]
  assign _T_6272 = _T_6248[23]; // @[Bitwise.scala 50:65:@6306.4]
  assign _T_6273 = _T_6248[24]; // @[Bitwise.scala 50:65:@6307.4]
  assign _T_6274 = _T_6248[25]; // @[Bitwise.scala 50:65:@6308.4]
  assign _T_6275 = _T_6248[26]; // @[Bitwise.scala 50:65:@6309.4]
  assign _T_6276 = _T_6248[27]; // @[Bitwise.scala 50:65:@6310.4]
  assign _T_6277 = _T_6248[28]; // @[Bitwise.scala 50:65:@6311.4]
  assign _T_6278 = _T_6248[29]; // @[Bitwise.scala 50:65:@6312.4]
  assign _T_6279 = _T_6248[30]; // @[Bitwise.scala 50:65:@6313.4]
  assign _T_6280 = _T_6248[31]; // @[Bitwise.scala 50:65:@6314.4]
  assign _T_6281 = _T_6248[32]; // @[Bitwise.scala 50:65:@6315.4]
  assign _T_6282 = _T_6248[33]; // @[Bitwise.scala 50:65:@6316.4]
  assign _T_6283 = _T_6248[34]; // @[Bitwise.scala 50:65:@6317.4]
  assign _T_6284 = _T_6248[35]; // @[Bitwise.scala 50:65:@6318.4]
  assign _T_6285 = _T_6248[36]; // @[Bitwise.scala 50:65:@6319.4]
  assign _T_6286 = _T_6248[37]; // @[Bitwise.scala 50:65:@6320.4]
  assign _T_6287 = _T_6248[38]; // @[Bitwise.scala 50:65:@6321.4]
  assign _T_6288 = _T_6248[39]; // @[Bitwise.scala 50:65:@6322.4]
  assign _T_6289 = _T_6249 + _T_6250; // @[Bitwise.scala 48:55:@6323.4]
  assign _T_6290 = _T_6252 + _T_6253; // @[Bitwise.scala 48:55:@6324.4]
  assign _GEN_733 = {{1'd0}, _T_6251}; // @[Bitwise.scala 48:55:@6325.4]
  assign _T_6291 = _GEN_733 + _T_6290; // @[Bitwise.scala 48:55:@6325.4]
  assign _GEN_734 = {{1'd0}, _T_6289}; // @[Bitwise.scala 48:55:@6326.4]
  assign _T_6292 = _GEN_734 + _T_6291; // @[Bitwise.scala 48:55:@6326.4]
  assign _T_6293 = _T_6254 + _T_6255; // @[Bitwise.scala 48:55:@6327.4]
  assign _T_6294 = _T_6257 + _T_6258; // @[Bitwise.scala 48:55:@6328.4]
  assign _GEN_735 = {{1'd0}, _T_6256}; // @[Bitwise.scala 48:55:@6329.4]
  assign _T_6295 = _GEN_735 + _T_6294; // @[Bitwise.scala 48:55:@6329.4]
  assign _GEN_736 = {{1'd0}, _T_6293}; // @[Bitwise.scala 48:55:@6330.4]
  assign _T_6296 = _GEN_736 + _T_6295; // @[Bitwise.scala 48:55:@6330.4]
  assign _T_6297 = _T_6292 + _T_6296; // @[Bitwise.scala 48:55:@6331.4]
  assign _T_6298 = _T_6259 + _T_6260; // @[Bitwise.scala 48:55:@6332.4]
  assign _T_6299 = _T_6262 + _T_6263; // @[Bitwise.scala 48:55:@6333.4]
  assign _GEN_737 = {{1'd0}, _T_6261}; // @[Bitwise.scala 48:55:@6334.4]
  assign _T_6300 = _GEN_737 + _T_6299; // @[Bitwise.scala 48:55:@6334.4]
  assign _GEN_738 = {{1'd0}, _T_6298}; // @[Bitwise.scala 48:55:@6335.4]
  assign _T_6301 = _GEN_738 + _T_6300; // @[Bitwise.scala 48:55:@6335.4]
  assign _T_6302 = _T_6264 + _T_6265; // @[Bitwise.scala 48:55:@6336.4]
  assign _T_6303 = _T_6267 + _T_6268; // @[Bitwise.scala 48:55:@6337.4]
  assign _GEN_739 = {{1'd0}, _T_6266}; // @[Bitwise.scala 48:55:@6338.4]
  assign _T_6304 = _GEN_739 + _T_6303; // @[Bitwise.scala 48:55:@6338.4]
  assign _GEN_740 = {{1'd0}, _T_6302}; // @[Bitwise.scala 48:55:@6339.4]
  assign _T_6305 = _GEN_740 + _T_6304; // @[Bitwise.scala 48:55:@6339.4]
  assign _T_6306 = _T_6301 + _T_6305; // @[Bitwise.scala 48:55:@6340.4]
  assign _T_6307 = _T_6297 + _T_6306; // @[Bitwise.scala 48:55:@6341.4]
  assign _T_6308 = _T_6269 + _T_6270; // @[Bitwise.scala 48:55:@6342.4]
  assign _T_6309 = _T_6272 + _T_6273; // @[Bitwise.scala 48:55:@6343.4]
  assign _GEN_741 = {{1'd0}, _T_6271}; // @[Bitwise.scala 48:55:@6344.4]
  assign _T_6310 = _GEN_741 + _T_6309; // @[Bitwise.scala 48:55:@6344.4]
  assign _GEN_742 = {{1'd0}, _T_6308}; // @[Bitwise.scala 48:55:@6345.4]
  assign _T_6311 = _GEN_742 + _T_6310; // @[Bitwise.scala 48:55:@6345.4]
  assign _T_6312 = _T_6274 + _T_6275; // @[Bitwise.scala 48:55:@6346.4]
  assign _T_6313 = _T_6277 + _T_6278; // @[Bitwise.scala 48:55:@6347.4]
  assign _GEN_743 = {{1'd0}, _T_6276}; // @[Bitwise.scala 48:55:@6348.4]
  assign _T_6314 = _GEN_743 + _T_6313; // @[Bitwise.scala 48:55:@6348.4]
  assign _GEN_744 = {{1'd0}, _T_6312}; // @[Bitwise.scala 48:55:@6349.4]
  assign _T_6315 = _GEN_744 + _T_6314; // @[Bitwise.scala 48:55:@6349.4]
  assign _T_6316 = _T_6311 + _T_6315; // @[Bitwise.scala 48:55:@6350.4]
  assign _T_6317 = _T_6279 + _T_6280; // @[Bitwise.scala 48:55:@6351.4]
  assign _T_6318 = _T_6282 + _T_6283; // @[Bitwise.scala 48:55:@6352.4]
  assign _GEN_745 = {{1'd0}, _T_6281}; // @[Bitwise.scala 48:55:@6353.4]
  assign _T_6319 = _GEN_745 + _T_6318; // @[Bitwise.scala 48:55:@6353.4]
  assign _GEN_746 = {{1'd0}, _T_6317}; // @[Bitwise.scala 48:55:@6354.4]
  assign _T_6320 = _GEN_746 + _T_6319; // @[Bitwise.scala 48:55:@6354.4]
  assign _T_6321 = _T_6284 + _T_6285; // @[Bitwise.scala 48:55:@6355.4]
  assign _T_6322 = _T_6287 + _T_6288; // @[Bitwise.scala 48:55:@6356.4]
  assign _GEN_747 = {{1'd0}, _T_6286}; // @[Bitwise.scala 48:55:@6357.4]
  assign _T_6323 = _GEN_747 + _T_6322; // @[Bitwise.scala 48:55:@6357.4]
  assign _GEN_748 = {{1'd0}, _T_6321}; // @[Bitwise.scala 48:55:@6358.4]
  assign _T_6324 = _GEN_748 + _T_6323; // @[Bitwise.scala 48:55:@6358.4]
  assign _T_6325 = _T_6320 + _T_6324; // @[Bitwise.scala 48:55:@6359.4]
  assign _T_6326 = _T_6316 + _T_6325; // @[Bitwise.scala 48:55:@6360.4]
  assign _T_6327 = _T_6307 + _T_6326; // @[Bitwise.scala 48:55:@6361.4]
  assign _T_6391 = _T_2230[40:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6426.4]
  assign _T_6392 = _T_6391[0]; // @[Bitwise.scala 50:65:@6427.4]
  assign _T_6393 = _T_6391[1]; // @[Bitwise.scala 50:65:@6428.4]
  assign _T_6394 = _T_6391[2]; // @[Bitwise.scala 50:65:@6429.4]
  assign _T_6395 = _T_6391[3]; // @[Bitwise.scala 50:65:@6430.4]
  assign _T_6396 = _T_6391[4]; // @[Bitwise.scala 50:65:@6431.4]
  assign _T_6397 = _T_6391[5]; // @[Bitwise.scala 50:65:@6432.4]
  assign _T_6398 = _T_6391[6]; // @[Bitwise.scala 50:65:@6433.4]
  assign _T_6399 = _T_6391[7]; // @[Bitwise.scala 50:65:@6434.4]
  assign _T_6400 = _T_6391[8]; // @[Bitwise.scala 50:65:@6435.4]
  assign _T_6401 = _T_6391[9]; // @[Bitwise.scala 50:65:@6436.4]
  assign _T_6402 = _T_6391[10]; // @[Bitwise.scala 50:65:@6437.4]
  assign _T_6403 = _T_6391[11]; // @[Bitwise.scala 50:65:@6438.4]
  assign _T_6404 = _T_6391[12]; // @[Bitwise.scala 50:65:@6439.4]
  assign _T_6405 = _T_6391[13]; // @[Bitwise.scala 50:65:@6440.4]
  assign _T_6406 = _T_6391[14]; // @[Bitwise.scala 50:65:@6441.4]
  assign _T_6407 = _T_6391[15]; // @[Bitwise.scala 50:65:@6442.4]
  assign _T_6408 = _T_6391[16]; // @[Bitwise.scala 50:65:@6443.4]
  assign _T_6409 = _T_6391[17]; // @[Bitwise.scala 50:65:@6444.4]
  assign _T_6410 = _T_6391[18]; // @[Bitwise.scala 50:65:@6445.4]
  assign _T_6411 = _T_6391[19]; // @[Bitwise.scala 50:65:@6446.4]
  assign _T_6412 = _T_6391[20]; // @[Bitwise.scala 50:65:@6447.4]
  assign _T_6413 = _T_6391[21]; // @[Bitwise.scala 50:65:@6448.4]
  assign _T_6414 = _T_6391[22]; // @[Bitwise.scala 50:65:@6449.4]
  assign _T_6415 = _T_6391[23]; // @[Bitwise.scala 50:65:@6450.4]
  assign _T_6416 = _T_6391[24]; // @[Bitwise.scala 50:65:@6451.4]
  assign _T_6417 = _T_6391[25]; // @[Bitwise.scala 50:65:@6452.4]
  assign _T_6418 = _T_6391[26]; // @[Bitwise.scala 50:65:@6453.4]
  assign _T_6419 = _T_6391[27]; // @[Bitwise.scala 50:65:@6454.4]
  assign _T_6420 = _T_6391[28]; // @[Bitwise.scala 50:65:@6455.4]
  assign _T_6421 = _T_6391[29]; // @[Bitwise.scala 50:65:@6456.4]
  assign _T_6422 = _T_6391[30]; // @[Bitwise.scala 50:65:@6457.4]
  assign _T_6423 = _T_6391[31]; // @[Bitwise.scala 50:65:@6458.4]
  assign _T_6424 = _T_6391[32]; // @[Bitwise.scala 50:65:@6459.4]
  assign _T_6425 = _T_6391[33]; // @[Bitwise.scala 50:65:@6460.4]
  assign _T_6426 = _T_6391[34]; // @[Bitwise.scala 50:65:@6461.4]
  assign _T_6427 = _T_6391[35]; // @[Bitwise.scala 50:65:@6462.4]
  assign _T_6428 = _T_6391[36]; // @[Bitwise.scala 50:65:@6463.4]
  assign _T_6429 = _T_6391[37]; // @[Bitwise.scala 50:65:@6464.4]
  assign _T_6430 = _T_6391[38]; // @[Bitwise.scala 50:65:@6465.4]
  assign _T_6431 = _T_6391[39]; // @[Bitwise.scala 50:65:@6466.4]
  assign _T_6432 = _T_6391[40]; // @[Bitwise.scala 50:65:@6467.4]
  assign _T_6433 = _T_6392 + _T_6393; // @[Bitwise.scala 48:55:@6468.4]
  assign _T_6434 = _T_6395 + _T_6396; // @[Bitwise.scala 48:55:@6469.4]
  assign _GEN_749 = {{1'd0}, _T_6394}; // @[Bitwise.scala 48:55:@6470.4]
  assign _T_6435 = _GEN_749 + _T_6434; // @[Bitwise.scala 48:55:@6470.4]
  assign _GEN_750 = {{1'd0}, _T_6433}; // @[Bitwise.scala 48:55:@6471.4]
  assign _T_6436 = _GEN_750 + _T_6435; // @[Bitwise.scala 48:55:@6471.4]
  assign _T_6437 = _T_6397 + _T_6398; // @[Bitwise.scala 48:55:@6472.4]
  assign _T_6438 = _T_6400 + _T_6401; // @[Bitwise.scala 48:55:@6473.4]
  assign _GEN_751 = {{1'd0}, _T_6399}; // @[Bitwise.scala 48:55:@6474.4]
  assign _T_6439 = _GEN_751 + _T_6438; // @[Bitwise.scala 48:55:@6474.4]
  assign _GEN_752 = {{1'd0}, _T_6437}; // @[Bitwise.scala 48:55:@6475.4]
  assign _T_6440 = _GEN_752 + _T_6439; // @[Bitwise.scala 48:55:@6475.4]
  assign _T_6441 = _T_6436 + _T_6440; // @[Bitwise.scala 48:55:@6476.4]
  assign _T_6442 = _T_6402 + _T_6403; // @[Bitwise.scala 48:55:@6477.4]
  assign _T_6443 = _T_6405 + _T_6406; // @[Bitwise.scala 48:55:@6478.4]
  assign _GEN_753 = {{1'd0}, _T_6404}; // @[Bitwise.scala 48:55:@6479.4]
  assign _T_6444 = _GEN_753 + _T_6443; // @[Bitwise.scala 48:55:@6479.4]
  assign _GEN_754 = {{1'd0}, _T_6442}; // @[Bitwise.scala 48:55:@6480.4]
  assign _T_6445 = _GEN_754 + _T_6444; // @[Bitwise.scala 48:55:@6480.4]
  assign _T_6446 = _T_6407 + _T_6408; // @[Bitwise.scala 48:55:@6481.4]
  assign _T_6447 = _T_6410 + _T_6411; // @[Bitwise.scala 48:55:@6482.4]
  assign _GEN_755 = {{1'd0}, _T_6409}; // @[Bitwise.scala 48:55:@6483.4]
  assign _T_6448 = _GEN_755 + _T_6447; // @[Bitwise.scala 48:55:@6483.4]
  assign _GEN_756 = {{1'd0}, _T_6446}; // @[Bitwise.scala 48:55:@6484.4]
  assign _T_6449 = _GEN_756 + _T_6448; // @[Bitwise.scala 48:55:@6484.4]
  assign _T_6450 = _T_6445 + _T_6449; // @[Bitwise.scala 48:55:@6485.4]
  assign _T_6451 = _T_6441 + _T_6450; // @[Bitwise.scala 48:55:@6486.4]
  assign _T_6452 = _T_6412 + _T_6413; // @[Bitwise.scala 48:55:@6487.4]
  assign _T_6453 = _T_6415 + _T_6416; // @[Bitwise.scala 48:55:@6488.4]
  assign _GEN_757 = {{1'd0}, _T_6414}; // @[Bitwise.scala 48:55:@6489.4]
  assign _T_6454 = _GEN_757 + _T_6453; // @[Bitwise.scala 48:55:@6489.4]
  assign _GEN_758 = {{1'd0}, _T_6452}; // @[Bitwise.scala 48:55:@6490.4]
  assign _T_6455 = _GEN_758 + _T_6454; // @[Bitwise.scala 48:55:@6490.4]
  assign _T_6456 = _T_6417 + _T_6418; // @[Bitwise.scala 48:55:@6491.4]
  assign _T_6457 = _T_6420 + _T_6421; // @[Bitwise.scala 48:55:@6492.4]
  assign _GEN_759 = {{1'd0}, _T_6419}; // @[Bitwise.scala 48:55:@6493.4]
  assign _T_6458 = _GEN_759 + _T_6457; // @[Bitwise.scala 48:55:@6493.4]
  assign _GEN_760 = {{1'd0}, _T_6456}; // @[Bitwise.scala 48:55:@6494.4]
  assign _T_6459 = _GEN_760 + _T_6458; // @[Bitwise.scala 48:55:@6494.4]
  assign _T_6460 = _T_6455 + _T_6459; // @[Bitwise.scala 48:55:@6495.4]
  assign _T_6461 = _T_6422 + _T_6423; // @[Bitwise.scala 48:55:@6496.4]
  assign _T_6462 = _T_6425 + _T_6426; // @[Bitwise.scala 48:55:@6497.4]
  assign _GEN_761 = {{1'd0}, _T_6424}; // @[Bitwise.scala 48:55:@6498.4]
  assign _T_6463 = _GEN_761 + _T_6462; // @[Bitwise.scala 48:55:@6498.4]
  assign _GEN_762 = {{1'd0}, _T_6461}; // @[Bitwise.scala 48:55:@6499.4]
  assign _T_6464 = _GEN_762 + _T_6463; // @[Bitwise.scala 48:55:@6499.4]
  assign _T_6465 = _T_6428 + _T_6429; // @[Bitwise.scala 48:55:@6500.4]
  assign _GEN_763 = {{1'd0}, _T_6427}; // @[Bitwise.scala 48:55:@6501.4]
  assign _T_6466 = _GEN_763 + _T_6465; // @[Bitwise.scala 48:55:@6501.4]
  assign _T_6467 = _T_6431 + _T_6432; // @[Bitwise.scala 48:55:@6502.4]
  assign _GEN_764 = {{1'd0}, _T_6430}; // @[Bitwise.scala 48:55:@6503.4]
  assign _T_6468 = _GEN_764 + _T_6467; // @[Bitwise.scala 48:55:@6503.4]
  assign _T_6469 = _T_6466 + _T_6468; // @[Bitwise.scala 48:55:@6504.4]
  assign _T_6470 = _T_6464 + _T_6469; // @[Bitwise.scala 48:55:@6505.4]
  assign _T_6471 = _T_6460 + _T_6470; // @[Bitwise.scala 48:55:@6506.4]
  assign _T_6472 = _T_6451 + _T_6471; // @[Bitwise.scala 48:55:@6507.4]
  assign _T_6536 = _T_2230[41:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6572.4]
  assign _T_6537 = _T_6536[0]; // @[Bitwise.scala 50:65:@6573.4]
  assign _T_6538 = _T_6536[1]; // @[Bitwise.scala 50:65:@6574.4]
  assign _T_6539 = _T_6536[2]; // @[Bitwise.scala 50:65:@6575.4]
  assign _T_6540 = _T_6536[3]; // @[Bitwise.scala 50:65:@6576.4]
  assign _T_6541 = _T_6536[4]; // @[Bitwise.scala 50:65:@6577.4]
  assign _T_6542 = _T_6536[5]; // @[Bitwise.scala 50:65:@6578.4]
  assign _T_6543 = _T_6536[6]; // @[Bitwise.scala 50:65:@6579.4]
  assign _T_6544 = _T_6536[7]; // @[Bitwise.scala 50:65:@6580.4]
  assign _T_6545 = _T_6536[8]; // @[Bitwise.scala 50:65:@6581.4]
  assign _T_6546 = _T_6536[9]; // @[Bitwise.scala 50:65:@6582.4]
  assign _T_6547 = _T_6536[10]; // @[Bitwise.scala 50:65:@6583.4]
  assign _T_6548 = _T_6536[11]; // @[Bitwise.scala 50:65:@6584.4]
  assign _T_6549 = _T_6536[12]; // @[Bitwise.scala 50:65:@6585.4]
  assign _T_6550 = _T_6536[13]; // @[Bitwise.scala 50:65:@6586.4]
  assign _T_6551 = _T_6536[14]; // @[Bitwise.scala 50:65:@6587.4]
  assign _T_6552 = _T_6536[15]; // @[Bitwise.scala 50:65:@6588.4]
  assign _T_6553 = _T_6536[16]; // @[Bitwise.scala 50:65:@6589.4]
  assign _T_6554 = _T_6536[17]; // @[Bitwise.scala 50:65:@6590.4]
  assign _T_6555 = _T_6536[18]; // @[Bitwise.scala 50:65:@6591.4]
  assign _T_6556 = _T_6536[19]; // @[Bitwise.scala 50:65:@6592.4]
  assign _T_6557 = _T_6536[20]; // @[Bitwise.scala 50:65:@6593.4]
  assign _T_6558 = _T_6536[21]; // @[Bitwise.scala 50:65:@6594.4]
  assign _T_6559 = _T_6536[22]; // @[Bitwise.scala 50:65:@6595.4]
  assign _T_6560 = _T_6536[23]; // @[Bitwise.scala 50:65:@6596.4]
  assign _T_6561 = _T_6536[24]; // @[Bitwise.scala 50:65:@6597.4]
  assign _T_6562 = _T_6536[25]; // @[Bitwise.scala 50:65:@6598.4]
  assign _T_6563 = _T_6536[26]; // @[Bitwise.scala 50:65:@6599.4]
  assign _T_6564 = _T_6536[27]; // @[Bitwise.scala 50:65:@6600.4]
  assign _T_6565 = _T_6536[28]; // @[Bitwise.scala 50:65:@6601.4]
  assign _T_6566 = _T_6536[29]; // @[Bitwise.scala 50:65:@6602.4]
  assign _T_6567 = _T_6536[30]; // @[Bitwise.scala 50:65:@6603.4]
  assign _T_6568 = _T_6536[31]; // @[Bitwise.scala 50:65:@6604.4]
  assign _T_6569 = _T_6536[32]; // @[Bitwise.scala 50:65:@6605.4]
  assign _T_6570 = _T_6536[33]; // @[Bitwise.scala 50:65:@6606.4]
  assign _T_6571 = _T_6536[34]; // @[Bitwise.scala 50:65:@6607.4]
  assign _T_6572 = _T_6536[35]; // @[Bitwise.scala 50:65:@6608.4]
  assign _T_6573 = _T_6536[36]; // @[Bitwise.scala 50:65:@6609.4]
  assign _T_6574 = _T_6536[37]; // @[Bitwise.scala 50:65:@6610.4]
  assign _T_6575 = _T_6536[38]; // @[Bitwise.scala 50:65:@6611.4]
  assign _T_6576 = _T_6536[39]; // @[Bitwise.scala 50:65:@6612.4]
  assign _T_6577 = _T_6536[40]; // @[Bitwise.scala 50:65:@6613.4]
  assign _T_6578 = _T_6536[41]; // @[Bitwise.scala 50:65:@6614.4]
  assign _T_6579 = _T_6537 + _T_6538; // @[Bitwise.scala 48:55:@6615.4]
  assign _T_6580 = _T_6540 + _T_6541; // @[Bitwise.scala 48:55:@6616.4]
  assign _GEN_765 = {{1'd0}, _T_6539}; // @[Bitwise.scala 48:55:@6617.4]
  assign _T_6581 = _GEN_765 + _T_6580; // @[Bitwise.scala 48:55:@6617.4]
  assign _GEN_766 = {{1'd0}, _T_6579}; // @[Bitwise.scala 48:55:@6618.4]
  assign _T_6582 = _GEN_766 + _T_6581; // @[Bitwise.scala 48:55:@6618.4]
  assign _T_6583 = _T_6542 + _T_6543; // @[Bitwise.scala 48:55:@6619.4]
  assign _T_6584 = _T_6545 + _T_6546; // @[Bitwise.scala 48:55:@6620.4]
  assign _GEN_767 = {{1'd0}, _T_6544}; // @[Bitwise.scala 48:55:@6621.4]
  assign _T_6585 = _GEN_767 + _T_6584; // @[Bitwise.scala 48:55:@6621.4]
  assign _GEN_768 = {{1'd0}, _T_6583}; // @[Bitwise.scala 48:55:@6622.4]
  assign _T_6586 = _GEN_768 + _T_6585; // @[Bitwise.scala 48:55:@6622.4]
  assign _T_6587 = _T_6582 + _T_6586; // @[Bitwise.scala 48:55:@6623.4]
  assign _T_6588 = _T_6547 + _T_6548; // @[Bitwise.scala 48:55:@6624.4]
  assign _T_6589 = _T_6550 + _T_6551; // @[Bitwise.scala 48:55:@6625.4]
  assign _GEN_769 = {{1'd0}, _T_6549}; // @[Bitwise.scala 48:55:@6626.4]
  assign _T_6590 = _GEN_769 + _T_6589; // @[Bitwise.scala 48:55:@6626.4]
  assign _GEN_770 = {{1'd0}, _T_6588}; // @[Bitwise.scala 48:55:@6627.4]
  assign _T_6591 = _GEN_770 + _T_6590; // @[Bitwise.scala 48:55:@6627.4]
  assign _T_6592 = _T_6553 + _T_6554; // @[Bitwise.scala 48:55:@6628.4]
  assign _GEN_771 = {{1'd0}, _T_6552}; // @[Bitwise.scala 48:55:@6629.4]
  assign _T_6593 = _GEN_771 + _T_6592; // @[Bitwise.scala 48:55:@6629.4]
  assign _T_6594 = _T_6556 + _T_6557; // @[Bitwise.scala 48:55:@6630.4]
  assign _GEN_772 = {{1'd0}, _T_6555}; // @[Bitwise.scala 48:55:@6631.4]
  assign _T_6595 = _GEN_772 + _T_6594; // @[Bitwise.scala 48:55:@6631.4]
  assign _T_6596 = _T_6593 + _T_6595; // @[Bitwise.scala 48:55:@6632.4]
  assign _T_6597 = _T_6591 + _T_6596; // @[Bitwise.scala 48:55:@6633.4]
  assign _T_6598 = _T_6587 + _T_6597; // @[Bitwise.scala 48:55:@6634.4]
  assign _T_6599 = _T_6558 + _T_6559; // @[Bitwise.scala 48:55:@6635.4]
  assign _T_6600 = _T_6561 + _T_6562; // @[Bitwise.scala 48:55:@6636.4]
  assign _GEN_773 = {{1'd0}, _T_6560}; // @[Bitwise.scala 48:55:@6637.4]
  assign _T_6601 = _GEN_773 + _T_6600; // @[Bitwise.scala 48:55:@6637.4]
  assign _GEN_774 = {{1'd0}, _T_6599}; // @[Bitwise.scala 48:55:@6638.4]
  assign _T_6602 = _GEN_774 + _T_6601; // @[Bitwise.scala 48:55:@6638.4]
  assign _T_6603 = _T_6563 + _T_6564; // @[Bitwise.scala 48:55:@6639.4]
  assign _T_6604 = _T_6566 + _T_6567; // @[Bitwise.scala 48:55:@6640.4]
  assign _GEN_775 = {{1'd0}, _T_6565}; // @[Bitwise.scala 48:55:@6641.4]
  assign _T_6605 = _GEN_775 + _T_6604; // @[Bitwise.scala 48:55:@6641.4]
  assign _GEN_776 = {{1'd0}, _T_6603}; // @[Bitwise.scala 48:55:@6642.4]
  assign _T_6606 = _GEN_776 + _T_6605; // @[Bitwise.scala 48:55:@6642.4]
  assign _T_6607 = _T_6602 + _T_6606; // @[Bitwise.scala 48:55:@6643.4]
  assign _T_6608 = _T_6568 + _T_6569; // @[Bitwise.scala 48:55:@6644.4]
  assign _T_6609 = _T_6571 + _T_6572; // @[Bitwise.scala 48:55:@6645.4]
  assign _GEN_777 = {{1'd0}, _T_6570}; // @[Bitwise.scala 48:55:@6646.4]
  assign _T_6610 = _GEN_777 + _T_6609; // @[Bitwise.scala 48:55:@6646.4]
  assign _GEN_778 = {{1'd0}, _T_6608}; // @[Bitwise.scala 48:55:@6647.4]
  assign _T_6611 = _GEN_778 + _T_6610; // @[Bitwise.scala 48:55:@6647.4]
  assign _T_6612 = _T_6574 + _T_6575; // @[Bitwise.scala 48:55:@6648.4]
  assign _GEN_779 = {{1'd0}, _T_6573}; // @[Bitwise.scala 48:55:@6649.4]
  assign _T_6613 = _GEN_779 + _T_6612; // @[Bitwise.scala 48:55:@6649.4]
  assign _T_6614 = _T_6577 + _T_6578; // @[Bitwise.scala 48:55:@6650.4]
  assign _GEN_780 = {{1'd0}, _T_6576}; // @[Bitwise.scala 48:55:@6651.4]
  assign _T_6615 = _GEN_780 + _T_6614; // @[Bitwise.scala 48:55:@6651.4]
  assign _T_6616 = _T_6613 + _T_6615; // @[Bitwise.scala 48:55:@6652.4]
  assign _T_6617 = _T_6611 + _T_6616; // @[Bitwise.scala 48:55:@6653.4]
  assign _T_6618 = _T_6607 + _T_6617; // @[Bitwise.scala 48:55:@6654.4]
  assign _T_6619 = _T_6598 + _T_6618; // @[Bitwise.scala 48:55:@6655.4]
  assign _T_6683 = _T_2230[42:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6720.4]
  assign _T_6684 = _T_6683[0]; // @[Bitwise.scala 50:65:@6721.4]
  assign _T_6685 = _T_6683[1]; // @[Bitwise.scala 50:65:@6722.4]
  assign _T_6686 = _T_6683[2]; // @[Bitwise.scala 50:65:@6723.4]
  assign _T_6687 = _T_6683[3]; // @[Bitwise.scala 50:65:@6724.4]
  assign _T_6688 = _T_6683[4]; // @[Bitwise.scala 50:65:@6725.4]
  assign _T_6689 = _T_6683[5]; // @[Bitwise.scala 50:65:@6726.4]
  assign _T_6690 = _T_6683[6]; // @[Bitwise.scala 50:65:@6727.4]
  assign _T_6691 = _T_6683[7]; // @[Bitwise.scala 50:65:@6728.4]
  assign _T_6692 = _T_6683[8]; // @[Bitwise.scala 50:65:@6729.4]
  assign _T_6693 = _T_6683[9]; // @[Bitwise.scala 50:65:@6730.4]
  assign _T_6694 = _T_6683[10]; // @[Bitwise.scala 50:65:@6731.4]
  assign _T_6695 = _T_6683[11]; // @[Bitwise.scala 50:65:@6732.4]
  assign _T_6696 = _T_6683[12]; // @[Bitwise.scala 50:65:@6733.4]
  assign _T_6697 = _T_6683[13]; // @[Bitwise.scala 50:65:@6734.4]
  assign _T_6698 = _T_6683[14]; // @[Bitwise.scala 50:65:@6735.4]
  assign _T_6699 = _T_6683[15]; // @[Bitwise.scala 50:65:@6736.4]
  assign _T_6700 = _T_6683[16]; // @[Bitwise.scala 50:65:@6737.4]
  assign _T_6701 = _T_6683[17]; // @[Bitwise.scala 50:65:@6738.4]
  assign _T_6702 = _T_6683[18]; // @[Bitwise.scala 50:65:@6739.4]
  assign _T_6703 = _T_6683[19]; // @[Bitwise.scala 50:65:@6740.4]
  assign _T_6704 = _T_6683[20]; // @[Bitwise.scala 50:65:@6741.4]
  assign _T_6705 = _T_6683[21]; // @[Bitwise.scala 50:65:@6742.4]
  assign _T_6706 = _T_6683[22]; // @[Bitwise.scala 50:65:@6743.4]
  assign _T_6707 = _T_6683[23]; // @[Bitwise.scala 50:65:@6744.4]
  assign _T_6708 = _T_6683[24]; // @[Bitwise.scala 50:65:@6745.4]
  assign _T_6709 = _T_6683[25]; // @[Bitwise.scala 50:65:@6746.4]
  assign _T_6710 = _T_6683[26]; // @[Bitwise.scala 50:65:@6747.4]
  assign _T_6711 = _T_6683[27]; // @[Bitwise.scala 50:65:@6748.4]
  assign _T_6712 = _T_6683[28]; // @[Bitwise.scala 50:65:@6749.4]
  assign _T_6713 = _T_6683[29]; // @[Bitwise.scala 50:65:@6750.4]
  assign _T_6714 = _T_6683[30]; // @[Bitwise.scala 50:65:@6751.4]
  assign _T_6715 = _T_6683[31]; // @[Bitwise.scala 50:65:@6752.4]
  assign _T_6716 = _T_6683[32]; // @[Bitwise.scala 50:65:@6753.4]
  assign _T_6717 = _T_6683[33]; // @[Bitwise.scala 50:65:@6754.4]
  assign _T_6718 = _T_6683[34]; // @[Bitwise.scala 50:65:@6755.4]
  assign _T_6719 = _T_6683[35]; // @[Bitwise.scala 50:65:@6756.4]
  assign _T_6720 = _T_6683[36]; // @[Bitwise.scala 50:65:@6757.4]
  assign _T_6721 = _T_6683[37]; // @[Bitwise.scala 50:65:@6758.4]
  assign _T_6722 = _T_6683[38]; // @[Bitwise.scala 50:65:@6759.4]
  assign _T_6723 = _T_6683[39]; // @[Bitwise.scala 50:65:@6760.4]
  assign _T_6724 = _T_6683[40]; // @[Bitwise.scala 50:65:@6761.4]
  assign _T_6725 = _T_6683[41]; // @[Bitwise.scala 50:65:@6762.4]
  assign _T_6726 = _T_6683[42]; // @[Bitwise.scala 50:65:@6763.4]
  assign _T_6727 = _T_6684 + _T_6685; // @[Bitwise.scala 48:55:@6764.4]
  assign _T_6728 = _T_6687 + _T_6688; // @[Bitwise.scala 48:55:@6765.4]
  assign _GEN_781 = {{1'd0}, _T_6686}; // @[Bitwise.scala 48:55:@6766.4]
  assign _T_6729 = _GEN_781 + _T_6728; // @[Bitwise.scala 48:55:@6766.4]
  assign _GEN_782 = {{1'd0}, _T_6727}; // @[Bitwise.scala 48:55:@6767.4]
  assign _T_6730 = _GEN_782 + _T_6729; // @[Bitwise.scala 48:55:@6767.4]
  assign _T_6731 = _T_6689 + _T_6690; // @[Bitwise.scala 48:55:@6768.4]
  assign _T_6732 = _T_6692 + _T_6693; // @[Bitwise.scala 48:55:@6769.4]
  assign _GEN_783 = {{1'd0}, _T_6691}; // @[Bitwise.scala 48:55:@6770.4]
  assign _T_6733 = _GEN_783 + _T_6732; // @[Bitwise.scala 48:55:@6770.4]
  assign _GEN_784 = {{1'd0}, _T_6731}; // @[Bitwise.scala 48:55:@6771.4]
  assign _T_6734 = _GEN_784 + _T_6733; // @[Bitwise.scala 48:55:@6771.4]
  assign _T_6735 = _T_6730 + _T_6734; // @[Bitwise.scala 48:55:@6772.4]
  assign _T_6736 = _T_6694 + _T_6695; // @[Bitwise.scala 48:55:@6773.4]
  assign _T_6737 = _T_6697 + _T_6698; // @[Bitwise.scala 48:55:@6774.4]
  assign _GEN_785 = {{1'd0}, _T_6696}; // @[Bitwise.scala 48:55:@6775.4]
  assign _T_6738 = _GEN_785 + _T_6737; // @[Bitwise.scala 48:55:@6775.4]
  assign _GEN_786 = {{1'd0}, _T_6736}; // @[Bitwise.scala 48:55:@6776.4]
  assign _T_6739 = _GEN_786 + _T_6738; // @[Bitwise.scala 48:55:@6776.4]
  assign _T_6740 = _T_6700 + _T_6701; // @[Bitwise.scala 48:55:@6777.4]
  assign _GEN_787 = {{1'd0}, _T_6699}; // @[Bitwise.scala 48:55:@6778.4]
  assign _T_6741 = _GEN_787 + _T_6740; // @[Bitwise.scala 48:55:@6778.4]
  assign _T_6742 = _T_6703 + _T_6704; // @[Bitwise.scala 48:55:@6779.4]
  assign _GEN_788 = {{1'd0}, _T_6702}; // @[Bitwise.scala 48:55:@6780.4]
  assign _T_6743 = _GEN_788 + _T_6742; // @[Bitwise.scala 48:55:@6780.4]
  assign _T_6744 = _T_6741 + _T_6743; // @[Bitwise.scala 48:55:@6781.4]
  assign _T_6745 = _T_6739 + _T_6744; // @[Bitwise.scala 48:55:@6782.4]
  assign _T_6746 = _T_6735 + _T_6745; // @[Bitwise.scala 48:55:@6783.4]
  assign _T_6747 = _T_6705 + _T_6706; // @[Bitwise.scala 48:55:@6784.4]
  assign _T_6748 = _T_6708 + _T_6709; // @[Bitwise.scala 48:55:@6785.4]
  assign _GEN_789 = {{1'd0}, _T_6707}; // @[Bitwise.scala 48:55:@6786.4]
  assign _T_6749 = _GEN_789 + _T_6748; // @[Bitwise.scala 48:55:@6786.4]
  assign _GEN_790 = {{1'd0}, _T_6747}; // @[Bitwise.scala 48:55:@6787.4]
  assign _T_6750 = _GEN_790 + _T_6749; // @[Bitwise.scala 48:55:@6787.4]
  assign _T_6751 = _T_6711 + _T_6712; // @[Bitwise.scala 48:55:@6788.4]
  assign _GEN_791 = {{1'd0}, _T_6710}; // @[Bitwise.scala 48:55:@6789.4]
  assign _T_6752 = _GEN_791 + _T_6751; // @[Bitwise.scala 48:55:@6789.4]
  assign _T_6753 = _T_6714 + _T_6715; // @[Bitwise.scala 48:55:@6790.4]
  assign _GEN_792 = {{1'd0}, _T_6713}; // @[Bitwise.scala 48:55:@6791.4]
  assign _T_6754 = _GEN_792 + _T_6753; // @[Bitwise.scala 48:55:@6791.4]
  assign _T_6755 = _T_6752 + _T_6754; // @[Bitwise.scala 48:55:@6792.4]
  assign _T_6756 = _T_6750 + _T_6755; // @[Bitwise.scala 48:55:@6793.4]
  assign _T_6757 = _T_6716 + _T_6717; // @[Bitwise.scala 48:55:@6794.4]
  assign _T_6758 = _T_6719 + _T_6720; // @[Bitwise.scala 48:55:@6795.4]
  assign _GEN_793 = {{1'd0}, _T_6718}; // @[Bitwise.scala 48:55:@6796.4]
  assign _T_6759 = _GEN_793 + _T_6758; // @[Bitwise.scala 48:55:@6796.4]
  assign _GEN_794 = {{1'd0}, _T_6757}; // @[Bitwise.scala 48:55:@6797.4]
  assign _T_6760 = _GEN_794 + _T_6759; // @[Bitwise.scala 48:55:@6797.4]
  assign _T_6761 = _T_6722 + _T_6723; // @[Bitwise.scala 48:55:@6798.4]
  assign _GEN_795 = {{1'd0}, _T_6721}; // @[Bitwise.scala 48:55:@6799.4]
  assign _T_6762 = _GEN_795 + _T_6761; // @[Bitwise.scala 48:55:@6799.4]
  assign _T_6763 = _T_6725 + _T_6726; // @[Bitwise.scala 48:55:@6800.4]
  assign _GEN_796 = {{1'd0}, _T_6724}; // @[Bitwise.scala 48:55:@6801.4]
  assign _T_6764 = _GEN_796 + _T_6763; // @[Bitwise.scala 48:55:@6801.4]
  assign _T_6765 = _T_6762 + _T_6764; // @[Bitwise.scala 48:55:@6802.4]
  assign _T_6766 = _T_6760 + _T_6765; // @[Bitwise.scala 48:55:@6803.4]
  assign _T_6767 = _T_6756 + _T_6766; // @[Bitwise.scala 48:55:@6804.4]
  assign _T_6768 = _T_6746 + _T_6767; // @[Bitwise.scala 48:55:@6805.4]
  assign _T_6832 = _T_2230[43:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6870.4]
  assign _T_6833 = _T_6832[0]; // @[Bitwise.scala 50:65:@6871.4]
  assign _T_6834 = _T_6832[1]; // @[Bitwise.scala 50:65:@6872.4]
  assign _T_6835 = _T_6832[2]; // @[Bitwise.scala 50:65:@6873.4]
  assign _T_6836 = _T_6832[3]; // @[Bitwise.scala 50:65:@6874.4]
  assign _T_6837 = _T_6832[4]; // @[Bitwise.scala 50:65:@6875.4]
  assign _T_6838 = _T_6832[5]; // @[Bitwise.scala 50:65:@6876.4]
  assign _T_6839 = _T_6832[6]; // @[Bitwise.scala 50:65:@6877.4]
  assign _T_6840 = _T_6832[7]; // @[Bitwise.scala 50:65:@6878.4]
  assign _T_6841 = _T_6832[8]; // @[Bitwise.scala 50:65:@6879.4]
  assign _T_6842 = _T_6832[9]; // @[Bitwise.scala 50:65:@6880.4]
  assign _T_6843 = _T_6832[10]; // @[Bitwise.scala 50:65:@6881.4]
  assign _T_6844 = _T_6832[11]; // @[Bitwise.scala 50:65:@6882.4]
  assign _T_6845 = _T_6832[12]; // @[Bitwise.scala 50:65:@6883.4]
  assign _T_6846 = _T_6832[13]; // @[Bitwise.scala 50:65:@6884.4]
  assign _T_6847 = _T_6832[14]; // @[Bitwise.scala 50:65:@6885.4]
  assign _T_6848 = _T_6832[15]; // @[Bitwise.scala 50:65:@6886.4]
  assign _T_6849 = _T_6832[16]; // @[Bitwise.scala 50:65:@6887.4]
  assign _T_6850 = _T_6832[17]; // @[Bitwise.scala 50:65:@6888.4]
  assign _T_6851 = _T_6832[18]; // @[Bitwise.scala 50:65:@6889.4]
  assign _T_6852 = _T_6832[19]; // @[Bitwise.scala 50:65:@6890.4]
  assign _T_6853 = _T_6832[20]; // @[Bitwise.scala 50:65:@6891.4]
  assign _T_6854 = _T_6832[21]; // @[Bitwise.scala 50:65:@6892.4]
  assign _T_6855 = _T_6832[22]; // @[Bitwise.scala 50:65:@6893.4]
  assign _T_6856 = _T_6832[23]; // @[Bitwise.scala 50:65:@6894.4]
  assign _T_6857 = _T_6832[24]; // @[Bitwise.scala 50:65:@6895.4]
  assign _T_6858 = _T_6832[25]; // @[Bitwise.scala 50:65:@6896.4]
  assign _T_6859 = _T_6832[26]; // @[Bitwise.scala 50:65:@6897.4]
  assign _T_6860 = _T_6832[27]; // @[Bitwise.scala 50:65:@6898.4]
  assign _T_6861 = _T_6832[28]; // @[Bitwise.scala 50:65:@6899.4]
  assign _T_6862 = _T_6832[29]; // @[Bitwise.scala 50:65:@6900.4]
  assign _T_6863 = _T_6832[30]; // @[Bitwise.scala 50:65:@6901.4]
  assign _T_6864 = _T_6832[31]; // @[Bitwise.scala 50:65:@6902.4]
  assign _T_6865 = _T_6832[32]; // @[Bitwise.scala 50:65:@6903.4]
  assign _T_6866 = _T_6832[33]; // @[Bitwise.scala 50:65:@6904.4]
  assign _T_6867 = _T_6832[34]; // @[Bitwise.scala 50:65:@6905.4]
  assign _T_6868 = _T_6832[35]; // @[Bitwise.scala 50:65:@6906.4]
  assign _T_6869 = _T_6832[36]; // @[Bitwise.scala 50:65:@6907.4]
  assign _T_6870 = _T_6832[37]; // @[Bitwise.scala 50:65:@6908.4]
  assign _T_6871 = _T_6832[38]; // @[Bitwise.scala 50:65:@6909.4]
  assign _T_6872 = _T_6832[39]; // @[Bitwise.scala 50:65:@6910.4]
  assign _T_6873 = _T_6832[40]; // @[Bitwise.scala 50:65:@6911.4]
  assign _T_6874 = _T_6832[41]; // @[Bitwise.scala 50:65:@6912.4]
  assign _T_6875 = _T_6832[42]; // @[Bitwise.scala 50:65:@6913.4]
  assign _T_6876 = _T_6832[43]; // @[Bitwise.scala 50:65:@6914.4]
  assign _T_6877 = _T_6833 + _T_6834; // @[Bitwise.scala 48:55:@6915.4]
  assign _T_6878 = _T_6836 + _T_6837; // @[Bitwise.scala 48:55:@6916.4]
  assign _GEN_797 = {{1'd0}, _T_6835}; // @[Bitwise.scala 48:55:@6917.4]
  assign _T_6879 = _GEN_797 + _T_6878; // @[Bitwise.scala 48:55:@6917.4]
  assign _GEN_798 = {{1'd0}, _T_6877}; // @[Bitwise.scala 48:55:@6918.4]
  assign _T_6880 = _GEN_798 + _T_6879; // @[Bitwise.scala 48:55:@6918.4]
  assign _T_6881 = _T_6839 + _T_6840; // @[Bitwise.scala 48:55:@6919.4]
  assign _GEN_799 = {{1'd0}, _T_6838}; // @[Bitwise.scala 48:55:@6920.4]
  assign _T_6882 = _GEN_799 + _T_6881; // @[Bitwise.scala 48:55:@6920.4]
  assign _T_6883 = _T_6842 + _T_6843; // @[Bitwise.scala 48:55:@6921.4]
  assign _GEN_800 = {{1'd0}, _T_6841}; // @[Bitwise.scala 48:55:@6922.4]
  assign _T_6884 = _GEN_800 + _T_6883; // @[Bitwise.scala 48:55:@6922.4]
  assign _T_6885 = _T_6882 + _T_6884; // @[Bitwise.scala 48:55:@6923.4]
  assign _T_6886 = _T_6880 + _T_6885; // @[Bitwise.scala 48:55:@6924.4]
  assign _T_6887 = _T_6844 + _T_6845; // @[Bitwise.scala 48:55:@6925.4]
  assign _T_6888 = _T_6847 + _T_6848; // @[Bitwise.scala 48:55:@6926.4]
  assign _GEN_801 = {{1'd0}, _T_6846}; // @[Bitwise.scala 48:55:@6927.4]
  assign _T_6889 = _GEN_801 + _T_6888; // @[Bitwise.scala 48:55:@6927.4]
  assign _GEN_802 = {{1'd0}, _T_6887}; // @[Bitwise.scala 48:55:@6928.4]
  assign _T_6890 = _GEN_802 + _T_6889; // @[Bitwise.scala 48:55:@6928.4]
  assign _T_6891 = _T_6850 + _T_6851; // @[Bitwise.scala 48:55:@6929.4]
  assign _GEN_803 = {{1'd0}, _T_6849}; // @[Bitwise.scala 48:55:@6930.4]
  assign _T_6892 = _GEN_803 + _T_6891; // @[Bitwise.scala 48:55:@6930.4]
  assign _T_6893 = _T_6853 + _T_6854; // @[Bitwise.scala 48:55:@6931.4]
  assign _GEN_804 = {{1'd0}, _T_6852}; // @[Bitwise.scala 48:55:@6932.4]
  assign _T_6894 = _GEN_804 + _T_6893; // @[Bitwise.scala 48:55:@6932.4]
  assign _T_6895 = _T_6892 + _T_6894; // @[Bitwise.scala 48:55:@6933.4]
  assign _T_6896 = _T_6890 + _T_6895; // @[Bitwise.scala 48:55:@6934.4]
  assign _T_6897 = _T_6886 + _T_6896; // @[Bitwise.scala 48:55:@6935.4]
  assign _T_6898 = _T_6855 + _T_6856; // @[Bitwise.scala 48:55:@6936.4]
  assign _T_6899 = _T_6858 + _T_6859; // @[Bitwise.scala 48:55:@6937.4]
  assign _GEN_805 = {{1'd0}, _T_6857}; // @[Bitwise.scala 48:55:@6938.4]
  assign _T_6900 = _GEN_805 + _T_6899; // @[Bitwise.scala 48:55:@6938.4]
  assign _GEN_806 = {{1'd0}, _T_6898}; // @[Bitwise.scala 48:55:@6939.4]
  assign _T_6901 = _GEN_806 + _T_6900; // @[Bitwise.scala 48:55:@6939.4]
  assign _T_6902 = _T_6861 + _T_6862; // @[Bitwise.scala 48:55:@6940.4]
  assign _GEN_807 = {{1'd0}, _T_6860}; // @[Bitwise.scala 48:55:@6941.4]
  assign _T_6903 = _GEN_807 + _T_6902; // @[Bitwise.scala 48:55:@6941.4]
  assign _T_6904 = _T_6864 + _T_6865; // @[Bitwise.scala 48:55:@6942.4]
  assign _GEN_808 = {{1'd0}, _T_6863}; // @[Bitwise.scala 48:55:@6943.4]
  assign _T_6905 = _GEN_808 + _T_6904; // @[Bitwise.scala 48:55:@6943.4]
  assign _T_6906 = _T_6903 + _T_6905; // @[Bitwise.scala 48:55:@6944.4]
  assign _T_6907 = _T_6901 + _T_6906; // @[Bitwise.scala 48:55:@6945.4]
  assign _T_6908 = _T_6866 + _T_6867; // @[Bitwise.scala 48:55:@6946.4]
  assign _T_6909 = _T_6869 + _T_6870; // @[Bitwise.scala 48:55:@6947.4]
  assign _GEN_809 = {{1'd0}, _T_6868}; // @[Bitwise.scala 48:55:@6948.4]
  assign _T_6910 = _GEN_809 + _T_6909; // @[Bitwise.scala 48:55:@6948.4]
  assign _GEN_810 = {{1'd0}, _T_6908}; // @[Bitwise.scala 48:55:@6949.4]
  assign _T_6911 = _GEN_810 + _T_6910; // @[Bitwise.scala 48:55:@6949.4]
  assign _T_6912 = _T_6872 + _T_6873; // @[Bitwise.scala 48:55:@6950.4]
  assign _GEN_811 = {{1'd0}, _T_6871}; // @[Bitwise.scala 48:55:@6951.4]
  assign _T_6913 = _GEN_811 + _T_6912; // @[Bitwise.scala 48:55:@6951.4]
  assign _T_6914 = _T_6875 + _T_6876; // @[Bitwise.scala 48:55:@6952.4]
  assign _GEN_812 = {{1'd0}, _T_6874}; // @[Bitwise.scala 48:55:@6953.4]
  assign _T_6915 = _GEN_812 + _T_6914; // @[Bitwise.scala 48:55:@6953.4]
  assign _T_6916 = _T_6913 + _T_6915; // @[Bitwise.scala 48:55:@6954.4]
  assign _T_6917 = _T_6911 + _T_6916; // @[Bitwise.scala 48:55:@6955.4]
  assign _T_6918 = _T_6907 + _T_6917; // @[Bitwise.scala 48:55:@6956.4]
  assign _T_6919 = _T_6897 + _T_6918; // @[Bitwise.scala 48:55:@6957.4]
  assign _T_6983 = _T_2230[44:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7022.4]
  assign _T_6984 = _T_6983[0]; // @[Bitwise.scala 50:65:@7023.4]
  assign _T_6985 = _T_6983[1]; // @[Bitwise.scala 50:65:@7024.4]
  assign _T_6986 = _T_6983[2]; // @[Bitwise.scala 50:65:@7025.4]
  assign _T_6987 = _T_6983[3]; // @[Bitwise.scala 50:65:@7026.4]
  assign _T_6988 = _T_6983[4]; // @[Bitwise.scala 50:65:@7027.4]
  assign _T_6989 = _T_6983[5]; // @[Bitwise.scala 50:65:@7028.4]
  assign _T_6990 = _T_6983[6]; // @[Bitwise.scala 50:65:@7029.4]
  assign _T_6991 = _T_6983[7]; // @[Bitwise.scala 50:65:@7030.4]
  assign _T_6992 = _T_6983[8]; // @[Bitwise.scala 50:65:@7031.4]
  assign _T_6993 = _T_6983[9]; // @[Bitwise.scala 50:65:@7032.4]
  assign _T_6994 = _T_6983[10]; // @[Bitwise.scala 50:65:@7033.4]
  assign _T_6995 = _T_6983[11]; // @[Bitwise.scala 50:65:@7034.4]
  assign _T_6996 = _T_6983[12]; // @[Bitwise.scala 50:65:@7035.4]
  assign _T_6997 = _T_6983[13]; // @[Bitwise.scala 50:65:@7036.4]
  assign _T_6998 = _T_6983[14]; // @[Bitwise.scala 50:65:@7037.4]
  assign _T_6999 = _T_6983[15]; // @[Bitwise.scala 50:65:@7038.4]
  assign _T_7000 = _T_6983[16]; // @[Bitwise.scala 50:65:@7039.4]
  assign _T_7001 = _T_6983[17]; // @[Bitwise.scala 50:65:@7040.4]
  assign _T_7002 = _T_6983[18]; // @[Bitwise.scala 50:65:@7041.4]
  assign _T_7003 = _T_6983[19]; // @[Bitwise.scala 50:65:@7042.4]
  assign _T_7004 = _T_6983[20]; // @[Bitwise.scala 50:65:@7043.4]
  assign _T_7005 = _T_6983[21]; // @[Bitwise.scala 50:65:@7044.4]
  assign _T_7006 = _T_6983[22]; // @[Bitwise.scala 50:65:@7045.4]
  assign _T_7007 = _T_6983[23]; // @[Bitwise.scala 50:65:@7046.4]
  assign _T_7008 = _T_6983[24]; // @[Bitwise.scala 50:65:@7047.4]
  assign _T_7009 = _T_6983[25]; // @[Bitwise.scala 50:65:@7048.4]
  assign _T_7010 = _T_6983[26]; // @[Bitwise.scala 50:65:@7049.4]
  assign _T_7011 = _T_6983[27]; // @[Bitwise.scala 50:65:@7050.4]
  assign _T_7012 = _T_6983[28]; // @[Bitwise.scala 50:65:@7051.4]
  assign _T_7013 = _T_6983[29]; // @[Bitwise.scala 50:65:@7052.4]
  assign _T_7014 = _T_6983[30]; // @[Bitwise.scala 50:65:@7053.4]
  assign _T_7015 = _T_6983[31]; // @[Bitwise.scala 50:65:@7054.4]
  assign _T_7016 = _T_6983[32]; // @[Bitwise.scala 50:65:@7055.4]
  assign _T_7017 = _T_6983[33]; // @[Bitwise.scala 50:65:@7056.4]
  assign _T_7018 = _T_6983[34]; // @[Bitwise.scala 50:65:@7057.4]
  assign _T_7019 = _T_6983[35]; // @[Bitwise.scala 50:65:@7058.4]
  assign _T_7020 = _T_6983[36]; // @[Bitwise.scala 50:65:@7059.4]
  assign _T_7021 = _T_6983[37]; // @[Bitwise.scala 50:65:@7060.4]
  assign _T_7022 = _T_6983[38]; // @[Bitwise.scala 50:65:@7061.4]
  assign _T_7023 = _T_6983[39]; // @[Bitwise.scala 50:65:@7062.4]
  assign _T_7024 = _T_6983[40]; // @[Bitwise.scala 50:65:@7063.4]
  assign _T_7025 = _T_6983[41]; // @[Bitwise.scala 50:65:@7064.4]
  assign _T_7026 = _T_6983[42]; // @[Bitwise.scala 50:65:@7065.4]
  assign _T_7027 = _T_6983[43]; // @[Bitwise.scala 50:65:@7066.4]
  assign _T_7028 = _T_6983[44]; // @[Bitwise.scala 50:65:@7067.4]
  assign _T_7029 = _T_6984 + _T_6985; // @[Bitwise.scala 48:55:@7068.4]
  assign _T_7030 = _T_6987 + _T_6988; // @[Bitwise.scala 48:55:@7069.4]
  assign _GEN_813 = {{1'd0}, _T_6986}; // @[Bitwise.scala 48:55:@7070.4]
  assign _T_7031 = _GEN_813 + _T_7030; // @[Bitwise.scala 48:55:@7070.4]
  assign _GEN_814 = {{1'd0}, _T_7029}; // @[Bitwise.scala 48:55:@7071.4]
  assign _T_7032 = _GEN_814 + _T_7031; // @[Bitwise.scala 48:55:@7071.4]
  assign _T_7033 = _T_6990 + _T_6991; // @[Bitwise.scala 48:55:@7072.4]
  assign _GEN_815 = {{1'd0}, _T_6989}; // @[Bitwise.scala 48:55:@7073.4]
  assign _T_7034 = _GEN_815 + _T_7033; // @[Bitwise.scala 48:55:@7073.4]
  assign _T_7035 = _T_6993 + _T_6994; // @[Bitwise.scala 48:55:@7074.4]
  assign _GEN_816 = {{1'd0}, _T_6992}; // @[Bitwise.scala 48:55:@7075.4]
  assign _T_7036 = _GEN_816 + _T_7035; // @[Bitwise.scala 48:55:@7075.4]
  assign _T_7037 = _T_7034 + _T_7036; // @[Bitwise.scala 48:55:@7076.4]
  assign _T_7038 = _T_7032 + _T_7037; // @[Bitwise.scala 48:55:@7077.4]
  assign _T_7039 = _T_6995 + _T_6996; // @[Bitwise.scala 48:55:@7078.4]
  assign _T_7040 = _T_6998 + _T_6999; // @[Bitwise.scala 48:55:@7079.4]
  assign _GEN_817 = {{1'd0}, _T_6997}; // @[Bitwise.scala 48:55:@7080.4]
  assign _T_7041 = _GEN_817 + _T_7040; // @[Bitwise.scala 48:55:@7080.4]
  assign _GEN_818 = {{1'd0}, _T_7039}; // @[Bitwise.scala 48:55:@7081.4]
  assign _T_7042 = _GEN_818 + _T_7041; // @[Bitwise.scala 48:55:@7081.4]
  assign _T_7043 = _T_7001 + _T_7002; // @[Bitwise.scala 48:55:@7082.4]
  assign _GEN_819 = {{1'd0}, _T_7000}; // @[Bitwise.scala 48:55:@7083.4]
  assign _T_7044 = _GEN_819 + _T_7043; // @[Bitwise.scala 48:55:@7083.4]
  assign _T_7045 = _T_7004 + _T_7005; // @[Bitwise.scala 48:55:@7084.4]
  assign _GEN_820 = {{1'd0}, _T_7003}; // @[Bitwise.scala 48:55:@7085.4]
  assign _T_7046 = _GEN_820 + _T_7045; // @[Bitwise.scala 48:55:@7085.4]
  assign _T_7047 = _T_7044 + _T_7046; // @[Bitwise.scala 48:55:@7086.4]
  assign _T_7048 = _T_7042 + _T_7047; // @[Bitwise.scala 48:55:@7087.4]
  assign _T_7049 = _T_7038 + _T_7048; // @[Bitwise.scala 48:55:@7088.4]
  assign _T_7050 = _T_7006 + _T_7007; // @[Bitwise.scala 48:55:@7089.4]
  assign _T_7051 = _T_7009 + _T_7010; // @[Bitwise.scala 48:55:@7090.4]
  assign _GEN_821 = {{1'd0}, _T_7008}; // @[Bitwise.scala 48:55:@7091.4]
  assign _T_7052 = _GEN_821 + _T_7051; // @[Bitwise.scala 48:55:@7091.4]
  assign _GEN_822 = {{1'd0}, _T_7050}; // @[Bitwise.scala 48:55:@7092.4]
  assign _T_7053 = _GEN_822 + _T_7052; // @[Bitwise.scala 48:55:@7092.4]
  assign _T_7054 = _T_7012 + _T_7013; // @[Bitwise.scala 48:55:@7093.4]
  assign _GEN_823 = {{1'd0}, _T_7011}; // @[Bitwise.scala 48:55:@7094.4]
  assign _T_7055 = _GEN_823 + _T_7054; // @[Bitwise.scala 48:55:@7094.4]
  assign _T_7056 = _T_7015 + _T_7016; // @[Bitwise.scala 48:55:@7095.4]
  assign _GEN_824 = {{1'd0}, _T_7014}; // @[Bitwise.scala 48:55:@7096.4]
  assign _T_7057 = _GEN_824 + _T_7056; // @[Bitwise.scala 48:55:@7096.4]
  assign _T_7058 = _T_7055 + _T_7057; // @[Bitwise.scala 48:55:@7097.4]
  assign _T_7059 = _T_7053 + _T_7058; // @[Bitwise.scala 48:55:@7098.4]
  assign _T_7060 = _T_7018 + _T_7019; // @[Bitwise.scala 48:55:@7099.4]
  assign _GEN_825 = {{1'd0}, _T_7017}; // @[Bitwise.scala 48:55:@7100.4]
  assign _T_7061 = _GEN_825 + _T_7060; // @[Bitwise.scala 48:55:@7100.4]
  assign _T_7062 = _T_7021 + _T_7022; // @[Bitwise.scala 48:55:@7101.4]
  assign _GEN_826 = {{1'd0}, _T_7020}; // @[Bitwise.scala 48:55:@7102.4]
  assign _T_7063 = _GEN_826 + _T_7062; // @[Bitwise.scala 48:55:@7102.4]
  assign _T_7064 = _T_7061 + _T_7063; // @[Bitwise.scala 48:55:@7103.4]
  assign _T_7065 = _T_7024 + _T_7025; // @[Bitwise.scala 48:55:@7104.4]
  assign _GEN_827 = {{1'd0}, _T_7023}; // @[Bitwise.scala 48:55:@7105.4]
  assign _T_7066 = _GEN_827 + _T_7065; // @[Bitwise.scala 48:55:@7105.4]
  assign _T_7067 = _T_7027 + _T_7028; // @[Bitwise.scala 48:55:@7106.4]
  assign _GEN_828 = {{1'd0}, _T_7026}; // @[Bitwise.scala 48:55:@7107.4]
  assign _T_7068 = _GEN_828 + _T_7067; // @[Bitwise.scala 48:55:@7107.4]
  assign _T_7069 = _T_7066 + _T_7068; // @[Bitwise.scala 48:55:@7108.4]
  assign _T_7070 = _T_7064 + _T_7069; // @[Bitwise.scala 48:55:@7109.4]
  assign _T_7071 = _T_7059 + _T_7070; // @[Bitwise.scala 48:55:@7110.4]
  assign _T_7072 = _T_7049 + _T_7071; // @[Bitwise.scala 48:55:@7111.4]
  assign _T_7136 = _T_2230[45:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7176.4]
  assign _T_7137 = _T_7136[0]; // @[Bitwise.scala 50:65:@7177.4]
  assign _T_7138 = _T_7136[1]; // @[Bitwise.scala 50:65:@7178.4]
  assign _T_7139 = _T_7136[2]; // @[Bitwise.scala 50:65:@7179.4]
  assign _T_7140 = _T_7136[3]; // @[Bitwise.scala 50:65:@7180.4]
  assign _T_7141 = _T_7136[4]; // @[Bitwise.scala 50:65:@7181.4]
  assign _T_7142 = _T_7136[5]; // @[Bitwise.scala 50:65:@7182.4]
  assign _T_7143 = _T_7136[6]; // @[Bitwise.scala 50:65:@7183.4]
  assign _T_7144 = _T_7136[7]; // @[Bitwise.scala 50:65:@7184.4]
  assign _T_7145 = _T_7136[8]; // @[Bitwise.scala 50:65:@7185.4]
  assign _T_7146 = _T_7136[9]; // @[Bitwise.scala 50:65:@7186.4]
  assign _T_7147 = _T_7136[10]; // @[Bitwise.scala 50:65:@7187.4]
  assign _T_7148 = _T_7136[11]; // @[Bitwise.scala 50:65:@7188.4]
  assign _T_7149 = _T_7136[12]; // @[Bitwise.scala 50:65:@7189.4]
  assign _T_7150 = _T_7136[13]; // @[Bitwise.scala 50:65:@7190.4]
  assign _T_7151 = _T_7136[14]; // @[Bitwise.scala 50:65:@7191.4]
  assign _T_7152 = _T_7136[15]; // @[Bitwise.scala 50:65:@7192.4]
  assign _T_7153 = _T_7136[16]; // @[Bitwise.scala 50:65:@7193.4]
  assign _T_7154 = _T_7136[17]; // @[Bitwise.scala 50:65:@7194.4]
  assign _T_7155 = _T_7136[18]; // @[Bitwise.scala 50:65:@7195.4]
  assign _T_7156 = _T_7136[19]; // @[Bitwise.scala 50:65:@7196.4]
  assign _T_7157 = _T_7136[20]; // @[Bitwise.scala 50:65:@7197.4]
  assign _T_7158 = _T_7136[21]; // @[Bitwise.scala 50:65:@7198.4]
  assign _T_7159 = _T_7136[22]; // @[Bitwise.scala 50:65:@7199.4]
  assign _T_7160 = _T_7136[23]; // @[Bitwise.scala 50:65:@7200.4]
  assign _T_7161 = _T_7136[24]; // @[Bitwise.scala 50:65:@7201.4]
  assign _T_7162 = _T_7136[25]; // @[Bitwise.scala 50:65:@7202.4]
  assign _T_7163 = _T_7136[26]; // @[Bitwise.scala 50:65:@7203.4]
  assign _T_7164 = _T_7136[27]; // @[Bitwise.scala 50:65:@7204.4]
  assign _T_7165 = _T_7136[28]; // @[Bitwise.scala 50:65:@7205.4]
  assign _T_7166 = _T_7136[29]; // @[Bitwise.scala 50:65:@7206.4]
  assign _T_7167 = _T_7136[30]; // @[Bitwise.scala 50:65:@7207.4]
  assign _T_7168 = _T_7136[31]; // @[Bitwise.scala 50:65:@7208.4]
  assign _T_7169 = _T_7136[32]; // @[Bitwise.scala 50:65:@7209.4]
  assign _T_7170 = _T_7136[33]; // @[Bitwise.scala 50:65:@7210.4]
  assign _T_7171 = _T_7136[34]; // @[Bitwise.scala 50:65:@7211.4]
  assign _T_7172 = _T_7136[35]; // @[Bitwise.scala 50:65:@7212.4]
  assign _T_7173 = _T_7136[36]; // @[Bitwise.scala 50:65:@7213.4]
  assign _T_7174 = _T_7136[37]; // @[Bitwise.scala 50:65:@7214.4]
  assign _T_7175 = _T_7136[38]; // @[Bitwise.scala 50:65:@7215.4]
  assign _T_7176 = _T_7136[39]; // @[Bitwise.scala 50:65:@7216.4]
  assign _T_7177 = _T_7136[40]; // @[Bitwise.scala 50:65:@7217.4]
  assign _T_7178 = _T_7136[41]; // @[Bitwise.scala 50:65:@7218.4]
  assign _T_7179 = _T_7136[42]; // @[Bitwise.scala 50:65:@7219.4]
  assign _T_7180 = _T_7136[43]; // @[Bitwise.scala 50:65:@7220.4]
  assign _T_7181 = _T_7136[44]; // @[Bitwise.scala 50:65:@7221.4]
  assign _T_7182 = _T_7136[45]; // @[Bitwise.scala 50:65:@7222.4]
  assign _T_7183 = _T_7137 + _T_7138; // @[Bitwise.scala 48:55:@7223.4]
  assign _T_7184 = _T_7140 + _T_7141; // @[Bitwise.scala 48:55:@7224.4]
  assign _GEN_829 = {{1'd0}, _T_7139}; // @[Bitwise.scala 48:55:@7225.4]
  assign _T_7185 = _GEN_829 + _T_7184; // @[Bitwise.scala 48:55:@7225.4]
  assign _GEN_830 = {{1'd0}, _T_7183}; // @[Bitwise.scala 48:55:@7226.4]
  assign _T_7186 = _GEN_830 + _T_7185; // @[Bitwise.scala 48:55:@7226.4]
  assign _T_7187 = _T_7143 + _T_7144; // @[Bitwise.scala 48:55:@7227.4]
  assign _GEN_831 = {{1'd0}, _T_7142}; // @[Bitwise.scala 48:55:@7228.4]
  assign _T_7188 = _GEN_831 + _T_7187; // @[Bitwise.scala 48:55:@7228.4]
  assign _T_7189 = _T_7146 + _T_7147; // @[Bitwise.scala 48:55:@7229.4]
  assign _GEN_832 = {{1'd0}, _T_7145}; // @[Bitwise.scala 48:55:@7230.4]
  assign _T_7190 = _GEN_832 + _T_7189; // @[Bitwise.scala 48:55:@7230.4]
  assign _T_7191 = _T_7188 + _T_7190; // @[Bitwise.scala 48:55:@7231.4]
  assign _T_7192 = _T_7186 + _T_7191; // @[Bitwise.scala 48:55:@7232.4]
  assign _T_7193 = _T_7149 + _T_7150; // @[Bitwise.scala 48:55:@7233.4]
  assign _GEN_833 = {{1'd0}, _T_7148}; // @[Bitwise.scala 48:55:@7234.4]
  assign _T_7194 = _GEN_833 + _T_7193; // @[Bitwise.scala 48:55:@7234.4]
  assign _T_7195 = _T_7152 + _T_7153; // @[Bitwise.scala 48:55:@7235.4]
  assign _GEN_834 = {{1'd0}, _T_7151}; // @[Bitwise.scala 48:55:@7236.4]
  assign _T_7196 = _GEN_834 + _T_7195; // @[Bitwise.scala 48:55:@7236.4]
  assign _T_7197 = _T_7194 + _T_7196; // @[Bitwise.scala 48:55:@7237.4]
  assign _T_7198 = _T_7155 + _T_7156; // @[Bitwise.scala 48:55:@7238.4]
  assign _GEN_835 = {{1'd0}, _T_7154}; // @[Bitwise.scala 48:55:@7239.4]
  assign _T_7199 = _GEN_835 + _T_7198; // @[Bitwise.scala 48:55:@7239.4]
  assign _T_7200 = _T_7158 + _T_7159; // @[Bitwise.scala 48:55:@7240.4]
  assign _GEN_836 = {{1'd0}, _T_7157}; // @[Bitwise.scala 48:55:@7241.4]
  assign _T_7201 = _GEN_836 + _T_7200; // @[Bitwise.scala 48:55:@7241.4]
  assign _T_7202 = _T_7199 + _T_7201; // @[Bitwise.scala 48:55:@7242.4]
  assign _T_7203 = _T_7197 + _T_7202; // @[Bitwise.scala 48:55:@7243.4]
  assign _T_7204 = _T_7192 + _T_7203; // @[Bitwise.scala 48:55:@7244.4]
  assign _T_7205 = _T_7160 + _T_7161; // @[Bitwise.scala 48:55:@7245.4]
  assign _T_7206 = _T_7163 + _T_7164; // @[Bitwise.scala 48:55:@7246.4]
  assign _GEN_837 = {{1'd0}, _T_7162}; // @[Bitwise.scala 48:55:@7247.4]
  assign _T_7207 = _GEN_837 + _T_7206; // @[Bitwise.scala 48:55:@7247.4]
  assign _GEN_838 = {{1'd0}, _T_7205}; // @[Bitwise.scala 48:55:@7248.4]
  assign _T_7208 = _GEN_838 + _T_7207; // @[Bitwise.scala 48:55:@7248.4]
  assign _T_7209 = _T_7166 + _T_7167; // @[Bitwise.scala 48:55:@7249.4]
  assign _GEN_839 = {{1'd0}, _T_7165}; // @[Bitwise.scala 48:55:@7250.4]
  assign _T_7210 = _GEN_839 + _T_7209; // @[Bitwise.scala 48:55:@7250.4]
  assign _T_7211 = _T_7169 + _T_7170; // @[Bitwise.scala 48:55:@7251.4]
  assign _GEN_840 = {{1'd0}, _T_7168}; // @[Bitwise.scala 48:55:@7252.4]
  assign _T_7212 = _GEN_840 + _T_7211; // @[Bitwise.scala 48:55:@7252.4]
  assign _T_7213 = _T_7210 + _T_7212; // @[Bitwise.scala 48:55:@7253.4]
  assign _T_7214 = _T_7208 + _T_7213; // @[Bitwise.scala 48:55:@7254.4]
  assign _T_7215 = _T_7172 + _T_7173; // @[Bitwise.scala 48:55:@7255.4]
  assign _GEN_841 = {{1'd0}, _T_7171}; // @[Bitwise.scala 48:55:@7256.4]
  assign _T_7216 = _GEN_841 + _T_7215; // @[Bitwise.scala 48:55:@7256.4]
  assign _T_7217 = _T_7175 + _T_7176; // @[Bitwise.scala 48:55:@7257.4]
  assign _GEN_842 = {{1'd0}, _T_7174}; // @[Bitwise.scala 48:55:@7258.4]
  assign _T_7218 = _GEN_842 + _T_7217; // @[Bitwise.scala 48:55:@7258.4]
  assign _T_7219 = _T_7216 + _T_7218; // @[Bitwise.scala 48:55:@7259.4]
  assign _T_7220 = _T_7178 + _T_7179; // @[Bitwise.scala 48:55:@7260.4]
  assign _GEN_843 = {{1'd0}, _T_7177}; // @[Bitwise.scala 48:55:@7261.4]
  assign _T_7221 = _GEN_843 + _T_7220; // @[Bitwise.scala 48:55:@7261.4]
  assign _T_7222 = _T_7181 + _T_7182; // @[Bitwise.scala 48:55:@7262.4]
  assign _GEN_844 = {{1'd0}, _T_7180}; // @[Bitwise.scala 48:55:@7263.4]
  assign _T_7223 = _GEN_844 + _T_7222; // @[Bitwise.scala 48:55:@7263.4]
  assign _T_7224 = _T_7221 + _T_7223; // @[Bitwise.scala 48:55:@7264.4]
  assign _T_7225 = _T_7219 + _T_7224; // @[Bitwise.scala 48:55:@7265.4]
  assign _T_7226 = _T_7214 + _T_7225; // @[Bitwise.scala 48:55:@7266.4]
  assign _T_7227 = _T_7204 + _T_7226; // @[Bitwise.scala 48:55:@7267.4]
  assign _T_7291 = _T_2230[46:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7332.4]
  assign _T_7292 = _T_7291[0]; // @[Bitwise.scala 50:65:@7333.4]
  assign _T_7293 = _T_7291[1]; // @[Bitwise.scala 50:65:@7334.4]
  assign _T_7294 = _T_7291[2]; // @[Bitwise.scala 50:65:@7335.4]
  assign _T_7295 = _T_7291[3]; // @[Bitwise.scala 50:65:@7336.4]
  assign _T_7296 = _T_7291[4]; // @[Bitwise.scala 50:65:@7337.4]
  assign _T_7297 = _T_7291[5]; // @[Bitwise.scala 50:65:@7338.4]
  assign _T_7298 = _T_7291[6]; // @[Bitwise.scala 50:65:@7339.4]
  assign _T_7299 = _T_7291[7]; // @[Bitwise.scala 50:65:@7340.4]
  assign _T_7300 = _T_7291[8]; // @[Bitwise.scala 50:65:@7341.4]
  assign _T_7301 = _T_7291[9]; // @[Bitwise.scala 50:65:@7342.4]
  assign _T_7302 = _T_7291[10]; // @[Bitwise.scala 50:65:@7343.4]
  assign _T_7303 = _T_7291[11]; // @[Bitwise.scala 50:65:@7344.4]
  assign _T_7304 = _T_7291[12]; // @[Bitwise.scala 50:65:@7345.4]
  assign _T_7305 = _T_7291[13]; // @[Bitwise.scala 50:65:@7346.4]
  assign _T_7306 = _T_7291[14]; // @[Bitwise.scala 50:65:@7347.4]
  assign _T_7307 = _T_7291[15]; // @[Bitwise.scala 50:65:@7348.4]
  assign _T_7308 = _T_7291[16]; // @[Bitwise.scala 50:65:@7349.4]
  assign _T_7309 = _T_7291[17]; // @[Bitwise.scala 50:65:@7350.4]
  assign _T_7310 = _T_7291[18]; // @[Bitwise.scala 50:65:@7351.4]
  assign _T_7311 = _T_7291[19]; // @[Bitwise.scala 50:65:@7352.4]
  assign _T_7312 = _T_7291[20]; // @[Bitwise.scala 50:65:@7353.4]
  assign _T_7313 = _T_7291[21]; // @[Bitwise.scala 50:65:@7354.4]
  assign _T_7314 = _T_7291[22]; // @[Bitwise.scala 50:65:@7355.4]
  assign _T_7315 = _T_7291[23]; // @[Bitwise.scala 50:65:@7356.4]
  assign _T_7316 = _T_7291[24]; // @[Bitwise.scala 50:65:@7357.4]
  assign _T_7317 = _T_7291[25]; // @[Bitwise.scala 50:65:@7358.4]
  assign _T_7318 = _T_7291[26]; // @[Bitwise.scala 50:65:@7359.4]
  assign _T_7319 = _T_7291[27]; // @[Bitwise.scala 50:65:@7360.4]
  assign _T_7320 = _T_7291[28]; // @[Bitwise.scala 50:65:@7361.4]
  assign _T_7321 = _T_7291[29]; // @[Bitwise.scala 50:65:@7362.4]
  assign _T_7322 = _T_7291[30]; // @[Bitwise.scala 50:65:@7363.4]
  assign _T_7323 = _T_7291[31]; // @[Bitwise.scala 50:65:@7364.4]
  assign _T_7324 = _T_7291[32]; // @[Bitwise.scala 50:65:@7365.4]
  assign _T_7325 = _T_7291[33]; // @[Bitwise.scala 50:65:@7366.4]
  assign _T_7326 = _T_7291[34]; // @[Bitwise.scala 50:65:@7367.4]
  assign _T_7327 = _T_7291[35]; // @[Bitwise.scala 50:65:@7368.4]
  assign _T_7328 = _T_7291[36]; // @[Bitwise.scala 50:65:@7369.4]
  assign _T_7329 = _T_7291[37]; // @[Bitwise.scala 50:65:@7370.4]
  assign _T_7330 = _T_7291[38]; // @[Bitwise.scala 50:65:@7371.4]
  assign _T_7331 = _T_7291[39]; // @[Bitwise.scala 50:65:@7372.4]
  assign _T_7332 = _T_7291[40]; // @[Bitwise.scala 50:65:@7373.4]
  assign _T_7333 = _T_7291[41]; // @[Bitwise.scala 50:65:@7374.4]
  assign _T_7334 = _T_7291[42]; // @[Bitwise.scala 50:65:@7375.4]
  assign _T_7335 = _T_7291[43]; // @[Bitwise.scala 50:65:@7376.4]
  assign _T_7336 = _T_7291[44]; // @[Bitwise.scala 50:65:@7377.4]
  assign _T_7337 = _T_7291[45]; // @[Bitwise.scala 50:65:@7378.4]
  assign _T_7338 = _T_7291[46]; // @[Bitwise.scala 50:65:@7379.4]
  assign _T_7339 = _T_7292 + _T_7293; // @[Bitwise.scala 48:55:@7380.4]
  assign _T_7340 = _T_7295 + _T_7296; // @[Bitwise.scala 48:55:@7381.4]
  assign _GEN_845 = {{1'd0}, _T_7294}; // @[Bitwise.scala 48:55:@7382.4]
  assign _T_7341 = _GEN_845 + _T_7340; // @[Bitwise.scala 48:55:@7382.4]
  assign _GEN_846 = {{1'd0}, _T_7339}; // @[Bitwise.scala 48:55:@7383.4]
  assign _T_7342 = _GEN_846 + _T_7341; // @[Bitwise.scala 48:55:@7383.4]
  assign _T_7343 = _T_7298 + _T_7299; // @[Bitwise.scala 48:55:@7384.4]
  assign _GEN_847 = {{1'd0}, _T_7297}; // @[Bitwise.scala 48:55:@7385.4]
  assign _T_7344 = _GEN_847 + _T_7343; // @[Bitwise.scala 48:55:@7385.4]
  assign _T_7345 = _T_7301 + _T_7302; // @[Bitwise.scala 48:55:@7386.4]
  assign _GEN_848 = {{1'd0}, _T_7300}; // @[Bitwise.scala 48:55:@7387.4]
  assign _T_7346 = _GEN_848 + _T_7345; // @[Bitwise.scala 48:55:@7387.4]
  assign _T_7347 = _T_7344 + _T_7346; // @[Bitwise.scala 48:55:@7388.4]
  assign _T_7348 = _T_7342 + _T_7347; // @[Bitwise.scala 48:55:@7389.4]
  assign _T_7349 = _T_7304 + _T_7305; // @[Bitwise.scala 48:55:@7390.4]
  assign _GEN_849 = {{1'd0}, _T_7303}; // @[Bitwise.scala 48:55:@7391.4]
  assign _T_7350 = _GEN_849 + _T_7349; // @[Bitwise.scala 48:55:@7391.4]
  assign _T_7351 = _T_7307 + _T_7308; // @[Bitwise.scala 48:55:@7392.4]
  assign _GEN_850 = {{1'd0}, _T_7306}; // @[Bitwise.scala 48:55:@7393.4]
  assign _T_7352 = _GEN_850 + _T_7351; // @[Bitwise.scala 48:55:@7393.4]
  assign _T_7353 = _T_7350 + _T_7352; // @[Bitwise.scala 48:55:@7394.4]
  assign _T_7354 = _T_7310 + _T_7311; // @[Bitwise.scala 48:55:@7395.4]
  assign _GEN_851 = {{1'd0}, _T_7309}; // @[Bitwise.scala 48:55:@7396.4]
  assign _T_7355 = _GEN_851 + _T_7354; // @[Bitwise.scala 48:55:@7396.4]
  assign _T_7356 = _T_7313 + _T_7314; // @[Bitwise.scala 48:55:@7397.4]
  assign _GEN_852 = {{1'd0}, _T_7312}; // @[Bitwise.scala 48:55:@7398.4]
  assign _T_7357 = _GEN_852 + _T_7356; // @[Bitwise.scala 48:55:@7398.4]
  assign _T_7358 = _T_7355 + _T_7357; // @[Bitwise.scala 48:55:@7399.4]
  assign _T_7359 = _T_7353 + _T_7358; // @[Bitwise.scala 48:55:@7400.4]
  assign _T_7360 = _T_7348 + _T_7359; // @[Bitwise.scala 48:55:@7401.4]
  assign _T_7361 = _T_7316 + _T_7317; // @[Bitwise.scala 48:55:@7402.4]
  assign _GEN_853 = {{1'd0}, _T_7315}; // @[Bitwise.scala 48:55:@7403.4]
  assign _T_7362 = _GEN_853 + _T_7361; // @[Bitwise.scala 48:55:@7403.4]
  assign _T_7363 = _T_7319 + _T_7320; // @[Bitwise.scala 48:55:@7404.4]
  assign _GEN_854 = {{1'd0}, _T_7318}; // @[Bitwise.scala 48:55:@7405.4]
  assign _T_7364 = _GEN_854 + _T_7363; // @[Bitwise.scala 48:55:@7405.4]
  assign _T_7365 = _T_7362 + _T_7364; // @[Bitwise.scala 48:55:@7406.4]
  assign _T_7366 = _T_7322 + _T_7323; // @[Bitwise.scala 48:55:@7407.4]
  assign _GEN_855 = {{1'd0}, _T_7321}; // @[Bitwise.scala 48:55:@7408.4]
  assign _T_7367 = _GEN_855 + _T_7366; // @[Bitwise.scala 48:55:@7408.4]
  assign _T_7368 = _T_7325 + _T_7326; // @[Bitwise.scala 48:55:@7409.4]
  assign _GEN_856 = {{1'd0}, _T_7324}; // @[Bitwise.scala 48:55:@7410.4]
  assign _T_7369 = _GEN_856 + _T_7368; // @[Bitwise.scala 48:55:@7410.4]
  assign _T_7370 = _T_7367 + _T_7369; // @[Bitwise.scala 48:55:@7411.4]
  assign _T_7371 = _T_7365 + _T_7370; // @[Bitwise.scala 48:55:@7412.4]
  assign _T_7372 = _T_7328 + _T_7329; // @[Bitwise.scala 48:55:@7413.4]
  assign _GEN_857 = {{1'd0}, _T_7327}; // @[Bitwise.scala 48:55:@7414.4]
  assign _T_7373 = _GEN_857 + _T_7372; // @[Bitwise.scala 48:55:@7414.4]
  assign _T_7374 = _T_7331 + _T_7332; // @[Bitwise.scala 48:55:@7415.4]
  assign _GEN_858 = {{1'd0}, _T_7330}; // @[Bitwise.scala 48:55:@7416.4]
  assign _T_7375 = _GEN_858 + _T_7374; // @[Bitwise.scala 48:55:@7416.4]
  assign _T_7376 = _T_7373 + _T_7375; // @[Bitwise.scala 48:55:@7417.4]
  assign _T_7377 = _T_7334 + _T_7335; // @[Bitwise.scala 48:55:@7418.4]
  assign _GEN_859 = {{1'd0}, _T_7333}; // @[Bitwise.scala 48:55:@7419.4]
  assign _T_7378 = _GEN_859 + _T_7377; // @[Bitwise.scala 48:55:@7419.4]
  assign _T_7379 = _T_7337 + _T_7338; // @[Bitwise.scala 48:55:@7420.4]
  assign _GEN_860 = {{1'd0}, _T_7336}; // @[Bitwise.scala 48:55:@7421.4]
  assign _T_7380 = _GEN_860 + _T_7379; // @[Bitwise.scala 48:55:@7421.4]
  assign _T_7381 = _T_7378 + _T_7380; // @[Bitwise.scala 48:55:@7422.4]
  assign _T_7382 = _T_7376 + _T_7381; // @[Bitwise.scala 48:55:@7423.4]
  assign _T_7383 = _T_7371 + _T_7382; // @[Bitwise.scala 48:55:@7424.4]
  assign _T_7384 = _T_7360 + _T_7383; // @[Bitwise.scala 48:55:@7425.4]
  assign _T_7448 = _T_2230[47:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7490.4]
  assign _T_7449 = _T_7448[0]; // @[Bitwise.scala 50:65:@7491.4]
  assign _T_7450 = _T_7448[1]; // @[Bitwise.scala 50:65:@7492.4]
  assign _T_7451 = _T_7448[2]; // @[Bitwise.scala 50:65:@7493.4]
  assign _T_7452 = _T_7448[3]; // @[Bitwise.scala 50:65:@7494.4]
  assign _T_7453 = _T_7448[4]; // @[Bitwise.scala 50:65:@7495.4]
  assign _T_7454 = _T_7448[5]; // @[Bitwise.scala 50:65:@7496.4]
  assign _T_7455 = _T_7448[6]; // @[Bitwise.scala 50:65:@7497.4]
  assign _T_7456 = _T_7448[7]; // @[Bitwise.scala 50:65:@7498.4]
  assign _T_7457 = _T_7448[8]; // @[Bitwise.scala 50:65:@7499.4]
  assign _T_7458 = _T_7448[9]; // @[Bitwise.scala 50:65:@7500.4]
  assign _T_7459 = _T_7448[10]; // @[Bitwise.scala 50:65:@7501.4]
  assign _T_7460 = _T_7448[11]; // @[Bitwise.scala 50:65:@7502.4]
  assign _T_7461 = _T_7448[12]; // @[Bitwise.scala 50:65:@7503.4]
  assign _T_7462 = _T_7448[13]; // @[Bitwise.scala 50:65:@7504.4]
  assign _T_7463 = _T_7448[14]; // @[Bitwise.scala 50:65:@7505.4]
  assign _T_7464 = _T_7448[15]; // @[Bitwise.scala 50:65:@7506.4]
  assign _T_7465 = _T_7448[16]; // @[Bitwise.scala 50:65:@7507.4]
  assign _T_7466 = _T_7448[17]; // @[Bitwise.scala 50:65:@7508.4]
  assign _T_7467 = _T_7448[18]; // @[Bitwise.scala 50:65:@7509.4]
  assign _T_7468 = _T_7448[19]; // @[Bitwise.scala 50:65:@7510.4]
  assign _T_7469 = _T_7448[20]; // @[Bitwise.scala 50:65:@7511.4]
  assign _T_7470 = _T_7448[21]; // @[Bitwise.scala 50:65:@7512.4]
  assign _T_7471 = _T_7448[22]; // @[Bitwise.scala 50:65:@7513.4]
  assign _T_7472 = _T_7448[23]; // @[Bitwise.scala 50:65:@7514.4]
  assign _T_7473 = _T_7448[24]; // @[Bitwise.scala 50:65:@7515.4]
  assign _T_7474 = _T_7448[25]; // @[Bitwise.scala 50:65:@7516.4]
  assign _T_7475 = _T_7448[26]; // @[Bitwise.scala 50:65:@7517.4]
  assign _T_7476 = _T_7448[27]; // @[Bitwise.scala 50:65:@7518.4]
  assign _T_7477 = _T_7448[28]; // @[Bitwise.scala 50:65:@7519.4]
  assign _T_7478 = _T_7448[29]; // @[Bitwise.scala 50:65:@7520.4]
  assign _T_7479 = _T_7448[30]; // @[Bitwise.scala 50:65:@7521.4]
  assign _T_7480 = _T_7448[31]; // @[Bitwise.scala 50:65:@7522.4]
  assign _T_7481 = _T_7448[32]; // @[Bitwise.scala 50:65:@7523.4]
  assign _T_7482 = _T_7448[33]; // @[Bitwise.scala 50:65:@7524.4]
  assign _T_7483 = _T_7448[34]; // @[Bitwise.scala 50:65:@7525.4]
  assign _T_7484 = _T_7448[35]; // @[Bitwise.scala 50:65:@7526.4]
  assign _T_7485 = _T_7448[36]; // @[Bitwise.scala 50:65:@7527.4]
  assign _T_7486 = _T_7448[37]; // @[Bitwise.scala 50:65:@7528.4]
  assign _T_7487 = _T_7448[38]; // @[Bitwise.scala 50:65:@7529.4]
  assign _T_7488 = _T_7448[39]; // @[Bitwise.scala 50:65:@7530.4]
  assign _T_7489 = _T_7448[40]; // @[Bitwise.scala 50:65:@7531.4]
  assign _T_7490 = _T_7448[41]; // @[Bitwise.scala 50:65:@7532.4]
  assign _T_7491 = _T_7448[42]; // @[Bitwise.scala 50:65:@7533.4]
  assign _T_7492 = _T_7448[43]; // @[Bitwise.scala 50:65:@7534.4]
  assign _T_7493 = _T_7448[44]; // @[Bitwise.scala 50:65:@7535.4]
  assign _T_7494 = _T_7448[45]; // @[Bitwise.scala 50:65:@7536.4]
  assign _T_7495 = _T_7448[46]; // @[Bitwise.scala 50:65:@7537.4]
  assign _T_7496 = _T_7448[47]; // @[Bitwise.scala 50:65:@7538.4]
  assign _T_7497 = _T_7450 + _T_7451; // @[Bitwise.scala 48:55:@7539.4]
  assign _GEN_861 = {{1'd0}, _T_7449}; // @[Bitwise.scala 48:55:@7540.4]
  assign _T_7498 = _GEN_861 + _T_7497; // @[Bitwise.scala 48:55:@7540.4]
  assign _T_7499 = _T_7453 + _T_7454; // @[Bitwise.scala 48:55:@7541.4]
  assign _GEN_862 = {{1'd0}, _T_7452}; // @[Bitwise.scala 48:55:@7542.4]
  assign _T_7500 = _GEN_862 + _T_7499; // @[Bitwise.scala 48:55:@7542.4]
  assign _T_7501 = _T_7498 + _T_7500; // @[Bitwise.scala 48:55:@7543.4]
  assign _T_7502 = _T_7456 + _T_7457; // @[Bitwise.scala 48:55:@7544.4]
  assign _GEN_863 = {{1'd0}, _T_7455}; // @[Bitwise.scala 48:55:@7545.4]
  assign _T_7503 = _GEN_863 + _T_7502; // @[Bitwise.scala 48:55:@7545.4]
  assign _T_7504 = _T_7459 + _T_7460; // @[Bitwise.scala 48:55:@7546.4]
  assign _GEN_864 = {{1'd0}, _T_7458}; // @[Bitwise.scala 48:55:@7547.4]
  assign _T_7505 = _GEN_864 + _T_7504; // @[Bitwise.scala 48:55:@7547.4]
  assign _T_7506 = _T_7503 + _T_7505; // @[Bitwise.scala 48:55:@7548.4]
  assign _T_7507 = _T_7501 + _T_7506; // @[Bitwise.scala 48:55:@7549.4]
  assign _T_7508 = _T_7462 + _T_7463; // @[Bitwise.scala 48:55:@7550.4]
  assign _GEN_865 = {{1'd0}, _T_7461}; // @[Bitwise.scala 48:55:@7551.4]
  assign _T_7509 = _GEN_865 + _T_7508; // @[Bitwise.scala 48:55:@7551.4]
  assign _T_7510 = _T_7465 + _T_7466; // @[Bitwise.scala 48:55:@7552.4]
  assign _GEN_866 = {{1'd0}, _T_7464}; // @[Bitwise.scala 48:55:@7553.4]
  assign _T_7511 = _GEN_866 + _T_7510; // @[Bitwise.scala 48:55:@7553.4]
  assign _T_7512 = _T_7509 + _T_7511; // @[Bitwise.scala 48:55:@7554.4]
  assign _T_7513 = _T_7468 + _T_7469; // @[Bitwise.scala 48:55:@7555.4]
  assign _GEN_867 = {{1'd0}, _T_7467}; // @[Bitwise.scala 48:55:@7556.4]
  assign _T_7514 = _GEN_867 + _T_7513; // @[Bitwise.scala 48:55:@7556.4]
  assign _T_7515 = _T_7471 + _T_7472; // @[Bitwise.scala 48:55:@7557.4]
  assign _GEN_868 = {{1'd0}, _T_7470}; // @[Bitwise.scala 48:55:@7558.4]
  assign _T_7516 = _GEN_868 + _T_7515; // @[Bitwise.scala 48:55:@7558.4]
  assign _T_7517 = _T_7514 + _T_7516; // @[Bitwise.scala 48:55:@7559.4]
  assign _T_7518 = _T_7512 + _T_7517; // @[Bitwise.scala 48:55:@7560.4]
  assign _T_7519 = _T_7507 + _T_7518; // @[Bitwise.scala 48:55:@7561.4]
  assign _T_7520 = _T_7474 + _T_7475; // @[Bitwise.scala 48:55:@7562.4]
  assign _GEN_869 = {{1'd0}, _T_7473}; // @[Bitwise.scala 48:55:@7563.4]
  assign _T_7521 = _GEN_869 + _T_7520; // @[Bitwise.scala 48:55:@7563.4]
  assign _T_7522 = _T_7477 + _T_7478; // @[Bitwise.scala 48:55:@7564.4]
  assign _GEN_870 = {{1'd0}, _T_7476}; // @[Bitwise.scala 48:55:@7565.4]
  assign _T_7523 = _GEN_870 + _T_7522; // @[Bitwise.scala 48:55:@7565.4]
  assign _T_7524 = _T_7521 + _T_7523; // @[Bitwise.scala 48:55:@7566.4]
  assign _T_7525 = _T_7480 + _T_7481; // @[Bitwise.scala 48:55:@7567.4]
  assign _GEN_871 = {{1'd0}, _T_7479}; // @[Bitwise.scala 48:55:@7568.4]
  assign _T_7526 = _GEN_871 + _T_7525; // @[Bitwise.scala 48:55:@7568.4]
  assign _T_7527 = _T_7483 + _T_7484; // @[Bitwise.scala 48:55:@7569.4]
  assign _GEN_872 = {{1'd0}, _T_7482}; // @[Bitwise.scala 48:55:@7570.4]
  assign _T_7528 = _GEN_872 + _T_7527; // @[Bitwise.scala 48:55:@7570.4]
  assign _T_7529 = _T_7526 + _T_7528; // @[Bitwise.scala 48:55:@7571.4]
  assign _T_7530 = _T_7524 + _T_7529; // @[Bitwise.scala 48:55:@7572.4]
  assign _T_7531 = _T_7486 + _T_7487; // @[Bitwise.scala 48:55:@7573.4]
  assign _GEN_873 = {{1'd0}, _T_7485}; // @[Bitwise.scala 48:55:@7574.4]
  assign _T_7532 = _GEN_873 + _T_7531; // @[Bitwise.scala 48:55:@7574.4]
  assign _T_7533 = _T_7489 + _T_7490; // @[Bitwise.scala 48:55:@7575.4]
  assign _GEN_874 = {{1'd0}, _T_7488}; // @[Bitwise.scala 48:55:@7576.4]
  assign _T_7534 = _GEN_874 + _T_7533; // @[Bitwise.scala 48:55:@7576.4]
  assign _T_7535 = _T_7532 + _T_7534; // @[Bitwise.scala 48:55:@7577.4]
  assign _T_7536 = _T_7492 + _T_7493; // @[Bitwise.scala 48:55:@7578.4]
  assign _GEN_875 = {{1'd0}, _T_7491}; // @[Bitwise.scala 48:55:@7579.4]
  assign _T_7537 = _GEN_875 + _T_7536; // @[Bitwise.scala 48:55:@7579.4]
  assign _T_7538 = _T_7495 + _T_7496; // @[Bitwise.scala 48:55:@7580.4]
  assign _GEN_876 = {{1'd0}, _T_7494}; // @[Bitwise.scala 48:55:@7581.4]
  assign _T_7539 = _GEN_876 + _T_7538; // @[Bitwise.scala 48:55:@7581.4]
  assign _T_7540 = _T_7537 + _T_7539; // @[Bitwise.scala 48:55:@7582.4]
  assign _T_7541 = _T_7535 + _T_7540; // @[Bitwise.scala 48:55:@7583.4]
  assign _T_7542 = _T_7530 + _T_7541; // @[Bitwise.scala 48:55:@7584.4]
  assign _T_7543 = _T_7519 + _T_7542; // @[Bitwise.scala 48:55:@7585.4]
  assign _T_7607 = _T_2230[48:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7650.4]
  assign _T_7608 = _T_7607[0]; // @[Bitwise.scala 50:65:@7651.4]
  assign _T_7609 = _T_7607[1]; // @[Bitwise.scala 50:65:@7652.4]
  assign _T_7610 = _T_7607[2]; // @[Bitwise.scala 50:65:@7653.4]
  assign _T_7611 = _T_7607[3]; // @[Bitwise.scala 50:65:@7654.4]
  assign _T_7612 = _T_7607[4]; // @[Bitwise.scala 50:65:@7655.4]
  assign _T_7613 = _T_7607[5]; // @[Bitwise.scala 50:65:@7656.4]
  assign _T_7614 = _T_7607[6]; // @[Bitwise.scala 50:65:@7657.4]
  assign _T_7615 = _T_7607[7]; // @[Bitwise.scala 50:65:@7658.4]
  assign _T_7616 = _T_7607[8]; // @[Bitwise.scala 50:65:@7659.4]
  assign _T_7617 = _T_7607[9]; // @[Bitwise.scala 50:65:@7660.4]
  assign _T_7618 = _T_7607[10]; // @[Bitwise.scala 50:65:@7661.4]
  assign _T_7619 = _T_7607[11]; // @[Bitwise.scala 50:65:@7662.4]
  assign _T_7620 = _T_7607[12]; // @[Bitwise.scala 50:65:@7663.4]
  assign _T_7621 = _T_7607[13]; // @[Bitwise.scala 50:65:@7664.4]
  assign _T_7622 = _T_7607[14]; // @[Bitwise.scala 50:65:@7665.4]
  assign _T_7623 = _T_7607[15]; // @[Bitwise.scala 50:65:@7666.4]
  assign _T_7624 = _T_7607[16]; // @[Bitwise.scala 50:65:@7667.4]
  assign _T_7625 = _T_7607[17]; // @[Bitwise.scala 50:65:@7668.4]
  assign _T_7626 = _T_7607[18]; // @[Bitwise.scala 50:65:@7669.4]
  assign _T_7627 = _T_7607[19]; // @[Bitwise.scala 50:65:@7670.4]
  assign _T_7628 = _T_7607[20]; // @[Bitwise.scala 50:65:@7671.4]
  assign _T_7629 = _T_7607[21]; // @[Bitwise.scala 50:65:@7672.4]
  assign _T_7630 = _T_7607[22]; // @[Bitwise.scala 50:65:@7673.4]
  assign _T_7631 = _T_7607[23]; // @[Bitwise.scala 50:65:@7674.4]
  assign _T_7632 = _T_7607[24]; // @[Bitwise.scala 50:65:@7675.4]
  assign _T_7633 = _T_7607[25]; // @[Bitwise.scala 50:65:@7676.4]
  assign _T_7634 = _T_7607[26]; // @[Bitwise.scala 50:65:@7677.4]
  assign _T_7635 = _T_7607[27]; // @[Bitwise.scala 50:65:@7678.4]
  assign _T_7636 = _T_7607[28]; // @[Bitwise.scala 50:65:@7679.4]
  assign _T_7637 = _T_7607[29]; // @[Bitwise.scala 50:65:@7680.4]
  assign _T_7638 = _T_7607[30]; // @[Bitwise.scala 50:65:@7681.4]
  assign _T_7639 = _T_7607[31]; // @[Bitwise.scala 50:65:@7682.4]
  assign _T_7640 = _T_7607[32]; // @[Bitwise.scala 50:65:@7683.4]
  assign _T_7641 = _T_7607[33]; // @[Bitwise.scala 50:65:@7684.4]
  assign _T_7642 = _T_7607[34]; // @[Bitwise.scala 50:65:@7685.4]
  assign _T_7643 = _T_7607[35]; // @[Bitwise.scala 50:65:@7686.4]
  assign _T_7644 = _T_7607[36]; // @[Bitwise.scala 50:65:@7687.4]
  assign _T_7645 = _T_7607[37]; // @[Bitwise.scala 50:65:@7688.4]
  assign _T_7646 = _T_7607[38]; // @[Bitwise.scala 50:65:@7689.4]
  assign _T_7647 = _T_7607[39]; // @[Bitwise.scala 50:65:@7690.4]
  assign _T_7648 = _T_7607[40]; // @[Bitwise.scala 50:65:@7691.4]
  assign _T_7649 = _T_7607[41]; // @[Bitwise.scala 50:65:@7692.4]
  assign _T_7650 = _T_7607[42]; // @[Bitwise.scala 50:65:@7693.4]
  assign _T_7651 = _T_7607[43]; // @[Bitwise.scala 50:65:@7694.4]
  assign _T_7652 = _T_7607[44]; // @[Bitwise.scala 50:65:@7695.4]
  assign _T_7653 = _T_7607[45]; // @[Bitwise.scala 50:65:@7696.4]
  assign _T_7654 = _T_7607[46]; // @[Bitwise.scala 50:65:@7697.4]
  assign _T_7655 = _T_7607[47]; // @[Bitwise.scala 50:65:@7698.4]
  assign _T_7656 = _T_7607[48]; // @[Bitwise.scala 50:65:@7699.4]
  assign _T_7657 = _T_7609 + _T_7610; // @[Bitwise.scala 48:55:@7700.4]
  assign _GEN_877 = {{1'd0}, _T_7608}; // @[Bitwise.scala 48:55:@7701.4]
  assign _T_7658 = _GEN_877 + _T_7657; // @[Bitwise.scala 48:55:@7701.4]
  assign _T_7659 = _T_7612 + _T_7613; // @[Bitwise.scala 48:55:@7702.4]
  assign _GEN_878 = {{1'd0}, _T_7611}; // @[Bitwise.scala 48:55:@7703.4]
  assign _T_7660 = _GEN_878 + _T_7659; // @[Bitwise.scala 48:55:@7703.4]
  assign _T_7661 = _T_7658 + _T_7660; // @[Bitwise.scala 48:55:@7704.4]
  assign _T_7662 = _T_7615 + _T_7616; // @[Bitwise.scala 48:55:@7705.4]
  assign _GEN_879 = {{1'd0}, _T_7614}; // @[Bitwise.scala 48:55:@7706.4]
  assign _T_7663 = _GEN_879 + _T_7662; // @[Bitwise.scala 48:55:@7706.4]
  assign _T_7664 = _T_7618 + _T_7619; // @[Bitwise.scala 48:55:@7707.4]
  assign _GEN_880 = {{1'd0}, _T_7617}; // @[Bitwise.scala 48:55:@7708.4]
  assign _T_7665 = _GEN_880 + _T_7664; // @[Bitwise.scala 48:55:@7708.4]
  assign _T_7666 = _T_7663 + _T_7665; // @[Bitwise.scala 48:55:@7709.4]
  assign _T_7667 = _T_7661 + _T_7666; // @[Bitwise.scala 48:55:@7710.4]
  assign _T_7668 = _T_7621 + _T_7622; // @[Bitwise.scala 48:55:@7711.4]
  assign _GEN_881 = {{1'd0}, _T_7620}; // @[Bitwise.scala 48:55:@7712.4]
  assign _T_7669 = _GEN_881 + _T_7668; // @[Bitwise.scala 48:55:@7712.4]
  assign _T_7670 = _T_7624 + _T_7625; // @[Bitwise.scala 48:55:@7713.4]
  assign _GEN_882 = {{1'd0}, _T_7623}; // @[Bitwise.scala 48:55:@7714.4]
  assign _T_7671 = _GEN_882 + _T_7670; // @[Bitwise.scala 48:55:@7714.4]
  assign _T_7672 = _T_7669 + _T_7671; // @[Bitwise.scala 48:55:@7715.4]
  assign _T_7673 = _T_7627 + _T_7628; // @[Bitwise.scala 48:55:@7716.4]
  assign _GEN_883 = {{1'd0}, _T_7626}; // @[Bitwise.scala 48:55:@7717.4]
  assign _T_7674 = _GEN_883 + _T_7673; // @[Bitwise.scala 48:55:@7717.4]
  assign _T_7675 = _T_7630 + _T_7631; // @[Bitwise.scala 48:55:@7718.4]
  assign _GEN_884 = {{1'd0}, _T_7629}; // @[Bitwise.scala 48:55:@7719.4]
  assign _T_7676 = _GEN_884 + _T_7675; // @[Bitwise.scala 48:55:@7719.4]
  assign _T_7677 = _T_7674 + _T_7676; // @[Bitwise.scala 48:55:@7720.4]
  assign _T_7678 = _T_7672 + _T_7677; // @[Bitwise.scala 48:55:@7721.4]
  assign _T_7679 = _T_7667 + _T_7678; // @[Bitwise.scala 48:55:@7722.4]
  assign _T_7680 = _T_7633 + _T_7634; // @[Bitwise.scala 48:55:@7723.4]
  assign _GEN_885 = {{1'd0}, _T_7632}; // @[Bitwise.scala 48:55:@7724.4]
  assign _T_7681 = _GEN_885 + _T_7680; // @[Bitwise.scala 48:55:@7724.4]
  assign _T_7682 = _T_7636 + _T_7637; // @[Bitwise.scala 48:55:@7725.4]
  assign _GEN_886 = {{1'd0}, _T_7635}; // @[Bitwise.scala 48:55:@7726.4]
  assign _T_7683 = _GEN_886 + _T_7682; // @[Bitwise.scala 48:55:@7726.4]
  assign _T_7684 = _T_7681 + _T_7683; // @[Bitwise.scala 48:55:@7727.4]
  assign _T_7685 = _T_7639 + _T_7640; // @[Bitwise.scala 48:55:@7728.4]
  assign _GEN_887 = {{1'd0}, _T_7638}; // @[Bitwise.scala 48:55:@7729.4]
  assign _T_7686 = _GEN_887 + _T_7685; // @[Bitwise.scala 48:55:@7729.4]
  assign _T_7687 = _T_7642 + _T_7643; // @[Bitwise.scala 48:55:@7730.4]
  assign _GEN_888 = {{1'd0}, _T_7641}; // @[Bitwise.scala 48:55:@7731.4]
  assign _T_7688 = _GEN_888 + _T_7687; // @[Bitwise.scala 48:55:@7731.4]
  assign _T_7689 = _T_7686 + _T_7688; // @[Bitwise.scala 48:55:@7732.4]
  assign _T_7690 = _T_7684 + _T_7689; // @[Bitwise.scala 48:55:@7733.4]
  assign _T_7691 = _T_7645 + _T_7646; // @[Bitwise.scala 48:55:@7734.4]
  assign _GEN_889 = {{1'd0}, _T_7644}; // @[Bitwise.scala 48:55:@7735.4]
  assign _T_7692 = _GEN_889 + _T_7691; // @[Bitwise.scala 48:55:@7735.4]
  assign _T_7693 = _T_7648 + _T_7649; // @[Bitwise.scala 48:55:@7736.4]
  assign _GEN_890 = {{1'd0}, _T_7647}; // @[Bitwise.scala 48:55:@7737.4]
  assign _T_7694 = _GEN_890 + _T_7693; // @[Bitwise.scala 48:55:@7737.4]
  assign _T_7695 = _T_7692 + _T_7694; // @[Bitwise.scala 48:55:@7738.4]
  assign _T_7696 = _T_7651 + _T_7652; // @[Bitwise.scala 48:55:@7739.4]
  assign _GEN_891 = {{1'd0}, _T_7650}; // @[Bitwise.scala 48:55:@7740.4]
  assign _T_7697 = _GEN_891 + _T_7696; // @[Bitwise.scala 48:55:@7740.4]
  assign _T_7698 = _T_7653 + _T_7654; // @[Bitwise.scala 48:55:@7741.4]
  assign _T_7699 = _T_7655 + _T_7656; // @[Bitwise.scala 48:55:@7742.4]
  assign _T_7700 = _T_7698 + _T_7699; // @[Bitwise.scala 48:55:@7743.4]
  assign _T_7701 = _T_7697 + _T_7700; // @[Bitwise.scala 48:55:@7744.4]
  assign _T_7702 = _T_7695 + _T_7701; // @[Bitwise.scala 48:55:@7745.4]
  assign _T_7703 = _T_7690 + _T_7702; // @[Bitwise.scala 48:55:@7746.4]
  assign _T_7704 = _T_7679 + _T_7703; // @[Bitwise.scala 48:55:@7747.4]
  assign _T_7768 = _T_2230[49:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7812.4]
  assign _T_7769 = _T_7768[0]; // @[Bitwise.scala 50:65:@7813.4]
  assign _T_7770 = _T_7768[1]; // @[Bitwise.scala 50:65:@7814.4]
  assign _T_7771 = _T_7768[2]; // @[Bitwise.scala 50:65:@7815.4]
  assign _T_7772 = _T_7768[3]; // @[Bitwise.scala 50:65:@7816.4]
  assign _T_7773 = _T_7768[4]; // @[Bitwise.scala 50:65:@7817.4]
  assign _T_7774 = _T_7768[5]; // @[Bitwise.scala 50:65:@7818.4]
  assign _T_7775 = _T_7768[6]; // @[Bitwise.scala 50:65:@7819.4]
  assign _T_7776 = _T_7768[7]; // @[Bitwise.scala 50:65:@7820.4]
  assign _T_7777 = _T_7768[8]; // @[Bitwise.scala 50:65:@7821.4]
  assign _T_7778 = _T_7768[9]; // @[Bitwise.scala 50:65:@7822.4]
  assign _T_7779 = _T_7768[10]; // @[Bitwise.scala 50:65:@7823.4]
  assign _T_7780 = _T_7768[11]; // @[Bitwise.scala 50:65:@7824.4]
  assign _T_7781 = _T_7768[12]; // @[Bitwise.scala 50:65:@7825.4]
  assign _T_7782 = _T_7768[13]; // @[Bitwise.scala 50:65:@7826.4]
  assign _T_7783 = _T_7768[14]; // @[Bitwise.scala 50:65:@7827.4]
  assign _T_7784 = _T_7768[15]; // @[Bitwise.scala 50:65:@7828.4]
  assign _T_7785 = _T_7768[16]; // @[Bitwise.scala 50:65:@7829.4]
  assign _T_7786 = _T_7768[17]; // @[Bitwise.scala 50:65:@7830.4]
  assign _T_7787 = _T_7768[18]; // @[Bitwise.scala 50:65:@7831.4]
  assign _T_7788 = _T_7768[19]; // @[Bitwise.scala 50:65:@7832.4]
  assign _T_7789 = _T_7768[20]; // @[Bitwise.scala 50:65:@7833.4]
  assign _T_7790 = _T_7768[21]; // @[Bitwise.scala 50:65:@7834.4]
  assign _T_7791 = _T_7768[22]; // @[Bitwise.scala 50:65:@7835.4]
  assign _T_7792 = _T_7768[23]; // @[Bitwise.scala 50:65:@7836.4]
  assign _T_7793 = _T_7768[24]; // @[Bitwise.scala 50:65:@7837.4]
  assign _T_7794 = _T_7768[25]; // @[Bitwise.scala 50:65:@7838.4]
  assign _T_7795 = _T_7768[26]; // @[Bitwise.scala 50:65:@7839.4]
  assign _T_7796 = _T_7768[27]; // @[Bitwise.scala 50:65:@7840.4]
  assign _T_7797 = _T_7768[28]; // @[Bitwise.scala 50:65:@7841.4]
  assign _T_7798 = _T_7768[29]; // @[Bitwise.scala 50:65:@7842.4]
  assign _T_7799 = _T_7768[30]; // @[Bitwise.scala 50:65:@7843.4]
  assign _T_7800 = _T_7768[31]; // @[Bitwise.scala 50:65:@7844.4]
  assign _T_7801 = _T_7768[32]; // @[Bitwise.scala 50:65:@7845.4]
  assign _T_7802 = _T_7768[33]; // @[Bitwise.scala 50:65:@7846.4]
  assign _T_7803 = _T_7768[34]; // @[Bitwise.scala 50:65:@7847.4]
  assign _T_7804 = _T_7768[35]; // @[Bitwise.scala 50:65:@7848.4]
  assign _T_7805 = _T_7768[36]; // @[Bitwise.scala 50:65:@7849.4]
  assign _T_7806 = _T_7768[37]; // @[Bitwise.scala 50:65:@7850.4]
  assign _T_7807 = _T_7768[38]; // @[Bitwise.scala 50:65:@7851.4]
  assign _T_7808 = _T_7768[39]; // @[Bitwise.scala 50:65:@7852.4]
  assign _T_7809 = _T_7768[40]; // @[Bitwise.scala 50:65:@7853.4]
  assign _T_7810 = _T_7768[41]; // @[Bitwise.scala 50:65:@7854.4]
  assign _T_7811 = _T_7768[42]; // @[Bitwise.scala 50:65:@7855.4]
  assign _T_7812 = _T_7768[43]; // @[Bitwise.scala 50:65:@7856.4]
  assign _T_7813 = _T_7768[44]; // @[Bitwise.scala 50:65:@7857.4]
  assign _T_7814 = _T_7768[45]; // @[Bitwise.scala 50:65:@7858.4]
  assign _T_7815 = _T_7768[46]; // @[Bitwise.scala 50:65:@7859.4]
  assign _T_7816 = _T_7768[47]; // @[Bitwise.scala 50:65:@7860.4]
  assign _T_7817 = _T_7768[48]; // @[Bitwise.scala 50:65:@7861.4]
  assign _T_7818 = _T_7768[49]; // @[Bitwise.scala 50:65:@7862.4]
  assign _T_7819 = _T_7770 + _T_7771; // @[Bitwise.scala 48:55:@7863.4]
  assign _GEN_892 = {{1'd0}, _T_7769}; // @[Bitwise.scala 48:55:@7864.4]
  assign _T_7820 = _GEN_892 + _T_7819; // @[Bitwise.scala 48:55:@7864.4]
  assign _T_7821 = _T_7773 + _T_7774; // @[Bitwise.scala 48:55:@7865.4]
  assign _GEN_893 = {{1'd0}, _T_7772}; // @[Bitwise.scala 48:55:@7866.4]
  assign _T_7822 = _GEN_893 + _T_7821; // @[Bitwise.scala 48:55:@7866.4]
  assign _T_7823 = _T_7820 + _T_7822; // @[Bitwise.scala 48:55:@7867.4]
  assign _T_7824 = _T_7776 + _T_7777; // @[Bitwise.scala 48:55:@7868.4]
  assign _GEN_894 = {{1'd0}, _T_7775}; // @[Bitwise.scala 48:55:@7869.4]
  assign _T_7825 = _GEN_894 + _T_7824; // @[Bitwise.scala 48:55:@7869.4]
  assign _T_7826 = _T_7779 + _T_7780; // @[Bitwise.scala 48:55:@7870.4]
  assign _GEN_895 = {{1'd0}, _T_7778}; // @[Bitwise.scala 48:55:@7871.4]
  assign _T_7827 = _GEN_895 + _T_7826; // @[Bitwise.scala 48:55:@7871.4]
  assign _T_7828 = _T_7825 + _T_7827; // @[Bitwise.scala 48:55:@7872.4]
  assign _T_7829 = _T_7823 + _T_7828; // @[Bitwise.scala 48:55:@7873.4]
  assign _T_7830 = _T_7782 + _T_7783; // @[Bitwise.scala 48:55:@7874.4]
  assign _GEN_896 = {{1'd0}, _T_7781}; // @[Bitwise.scala 48:55:@7875.4]
  assign _T_7831 = _GEN_896 + _T_7830; // @[Bitwise.scala 48:55:@7875.4]
  assign _T_7832 = _T_7785 + _T_7786; // @[Bitwise.scala 48:55:@7876.4]
  assign _GEN_897 = {{1'd0}, _T_7784}; // @[Bitwise.scala 48:55:@7877.4]
  assign _T_7833 = _GEN_897 + _T_7832; // @[Bitwise.scala 48:55:@7877.4]
  assign _T_7834 = _T_7831 + _T_7833; // @[Bitwise.scala 48:55:@7878.4]
  assign _T_7835 = _T_7788 + _T_7789; // @[Bitwise.scala 48:55:@7879.4]
  assign _GEN_898 = {{1'd0}, _T_7787}; // @[Bitwise.scala 48:55:@7880.4]
  assign _T_7836 = _GEN_898 + _T_7835; // @[Bitwise.scala 48:55:@7880.4]
  assign _T_7837 = _T_7790 + _T_7791; // @[Bitwise.scala 48:55:@7881.4]
  assign _T_7838 = _T_7792 + _T_7793; // @[Bitwise.scala 48:55:@7882.4]
  assign _T_7839 = _T_7837 + _T_7838; // @[Bitwise.scala 48:55:@7883.4]
  assign _T_7840 = _T_7836 + _T_7839; // @[Bitwise.scala 48:55:@7884.4]
  assign _T_7841 = _T_7834 + _T_7840; // @[Bitwise.scala 48:55:@7885.4]
  assign _T_7842 = _T_7829 + _T_7841; // @[Bitwise.scala 48:55:@7886.4]
  assign _T_7843 = _T_7795 + _T_7796; // @[Bitwise.scala 48:55:@7887.4]
  assign _GEN_899 = {{1'd0}, _T_7794}; // @[Bitwise.scala 48:55:@7888.4]
  assign _T_7844 = _GEN_899 + _T_7843; // @[Bitwise.scala 48:55:@7888.4]
  assign _T_7845 = _T_7798 + _T_7799; // @[Bitwise.scala 48:55:@7889.4]
  assign _GEN_900 = {{1'd0}, _T_7797}; // @[Bitwise.scala 48:55:@7890.4]
  assign _T_7846 = _GEN_900 + _T_7845; // @[Bitwise.scala 48:55:@7890.4]
  assign _T_7847 = _T_7844 + _T_7846; // @[Bitwise.scala 48:55:@7891.4]
  assign _T_7848 = _T_7801 + _T_7802; // @[Bitwise.scala 48:55:@7892.4]
  assign _GEN_901 = {{1'd0}, _T_7800}; // @[Bitwise.scala 48:55:@7893.4]
  assign _T_7849 = _GEN_901 + _T_7848; // @[Bitwise.scala 48:55:@7893.4]
  assign _T_7850 = _T_7804 + _T_7805; // @[Bitwise.scala 48:55:@7894.4]
  assign _GEN_902 = {{1'd0}, _T_7803}; // @[Bitwise.scala 48:55:@7895.4]
  assign _T_7851 = _GEN_902 + _T_7850; // @[Bitwise.scala 48:55:@7895.4]
  assign _T_7852 = _T_7849 + _T_7851; // @[Bitwise.scala 48:55:@7896.4]
  assign _T_7853 = _T_7847 + _T_7852; // @[Bitwise.scala 48:55:@7897.4]
  assign _T_7854 = _T_7807 + _T_7808; // @[Bitwise.scala 48:55:@7898.4]
  assign _GEN_903 = {{1'd0}, _T_7806}; // @[Bitwise.scala 48:55:@7899.4]
  assign _T_7855 = _GEN_903 + _T_7854; // @[Bitwise.scala 48:55:@7899.4]
  assign _T_7856 = _T_7810 + _T_7811; // @[Bitwise.scala 48:55:@7900.4]
  assign _GEN_904 = {{1'd0}, _T_7809}; // @[Bitwise.scala 48:55:@7901.4]
  assign _T_7857 = _GEN_904 + _T_7856; // @[Bitwise.scala 48:55:@7901.4]
  assign _T_7858 = _T_7855 + _T_7857; // @[Bitwise.scala 48:55:@7902.4]
  assign _T_7859 = _T_7813 + _T_7814; // @[Bitwise.scala 48:55:@7903.4]
  assign _GEN_905 = {{1'd0}, _T_7812}; // @[Bitwise.scala 48:55:@7904.4]
  assign _T_7860 = _GEN_905 + _T_7859; // @[Bitwise.scala 48:55:@7904.4]
  assign _T_7861 = _T_7815 + _T_7816; // @[Bitwise.scala 48:55:@7905.4]
  assign _T_7862 = _T_7817 + _T_7818; // @[Bitwise.scala 48:55:@7906.4]
  assign _T_7863 = _T_7861 + _T_7862; // @[Bitwise.scala 48:55:@7907.4]
  assign _T_7864 = _T_7860 + _T_7863; // @[Bitwise.scala 48:55:@7908.4]
  assign _T_7865 = _T_7858 + _T_7864; // @[Bitwise.scala 48:55:@7909.4]
  assign _T_7866 = _T_7853 + _T_7865; // @[Bitwise.scala 48:55:@7910.4]
  assign _T_7867 = _T_7842 + _T_7866; // @[Bitwise.scala 48:55:@7911.4]
  assign _T_7931 = _T_2230[50:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7976.4]
  assign _T_7932 = _T_7931[0]; // @[Bitwise.scala 50:65:@7977.4]
  assign _T_7933 = _T_7931[1]; // @[Bitwise.scala 50:65:@7978.4]
  assign _T_7934 = _T_7931[2]; // @[Bitwise.scala 50:65:@7979.4]
  assign _T_7935 = _T_7931[3]; // @[Bitwise.scala 50:65:@7980.4]
  assign _T_7936 = _T_7931[4]; // @[Bitwise.scala 50:65:@7981.4]
  assign _T_7937 = _T_7931[5]; // @[Bitwise.scala 50:65:@7982.4]
  assign _T_7938 = _T_7931[6]; // @[Bitwise.scala 50:65:@7983.4]
  assign _T_7939 = _T_7931[7]; // @[Bitwise.scala 50:65:@7984.4]
  assign _T_7940 = _T_7931[8]; // @[Bitwise.scala 50:65:@7985.4]
  assign _T_7941 = _T_7931[9]; // @[Bitwise.scala 50:65:@7986.4]
  assign _T_7942 = _T_7931[10]; // @[Bitwise.scala 50:65:@7987.4]
  assign _T_7943 = _T_7931[11]; // @[Bitwise.scala 50:65:@7988.4]
  assign _T_7944 = _T_7931[12]; // @[Bitwise.scala 50:65:@7989.4]
  assign _T_7945 = _T_7931[13]; // @[Bitwise.scala 50:65:@7990.4]
  assign _T_7946 = _T_7931[14]; // @[Bitwise.scala 50:65:@7991.4]
  assign _T_7947 = _T_7931[15]; // @[Bitwise.scala 50:65:@7992.4]
  assign _T_7948 = _T_7931[16]; // @[Bitwise.scala 50:65:@7993.4]
  assign _T_7949 = _T_7931[17]; // @[Bitwise.scala 50:65:@7994.4]
  assign _T_7950 = _T_7931[18]; // @[Bitwise.scala 50:65:@7995.4]
  assign _T_7951 = _T_7931[19]; // @[Bitwise.scala 50:65:@7996.4]
  assign _T_7952 = _T_7931[20]; // @[Bitwise.scala 50:65:@7997.4]
  assign _T_7953 = _T_7931[21]; // @[Bitwise.scala 50:65:@7998.4]
  assign _T_7954 = _T_7931[22]; // @[Bitwise.scala 50:65:@7999.4]
  assign _T_7955 = _T_7931[23]; // @[Bitwise.scala 50:65:@8000.4]
  assign _T_7956 = _T_7931[24]; // @[Bitwise.scala 50:65:@8001.4]
  assign _T_7957 = _T_7931[25]; // @[Bitwise.scala 50:65:@8002.4]
  assign _T_7958 = _T_7931[26]; // @[Bitwise.scala 50:65:@8003.4]
  assign _T_7959 = _T_7931[27]; // @[Bitwise.scala 50:65:@8004.4]
  assign _T_7960 = _T_7931[28]; // @[Bitwise.scala 50:65:@8005.4]
  assign _T_7961 = _T_7931[29]; // @[Bitwise.scala 50:65:@8006.4]
  assign _T_7962 = _T_7931[30]; // @[Bitwise.scala 50:65:@8007.4]
  assign _T_7963 = _T_7931[31]; // @[Bitwise.scala 50:65:@8008.4]
  assign _T_7964 = _T_7931[32]; // @[Bitwise.scala 50:65:@8009.4]
  assign _T_7965 = _T_7931[33]; // @[Bitwise.scala 50:65:@8010.4]
  assign _T_7966 = _T_7931[34]; // @[Bitwise.scala 50:65:@8011.4]
  assign _T_7967 = _T_7931[35]; // @[Bitwise.scala 50:65:@8012.4]
  assign _T_7968 = _T_7931[36]; // @[Bitwise.scala 50:65:@8013.4]
  assign _T_7969 = _T_7931[37]; // @[Bitwise.scala 50:65:@8014.4]
  assign _T_7970 = _T_7931[38]; // @[Bitwise.scala 50:65:@8015.4]
  assign _T_7971 = _T_7931[39]; // @[Bitwise.scala 50:65:@8016.4]
  assign _T_7972 = _T_7931[40]; // @[Bitwise.scala 50:65:@8017.4]
  assign _T_7973 = _T_7931[41]; // @[Bitwise.scala 50:65:@8018.4]
  assign _T_7974 = _T_7931[42]; // @[Bitwise.scala 50:65:@8019.4]
  assign _T_7975 = _T_7931[43]; // @[Bitwise.scala 50:65:@8020.4]
  assign _T_7976 = _T_7931[44]; // @[Bitwise.scala 50:65:@8021.4]
  assign _T_7977 = _T_7931[45]; // @[Bitwise.scala 50:65:@8022.4]
  assign _T_7978 = _T_7931[46]; // @[Bitwise.scala 50:65:@8023.4]
  assign _T_7979 = _T_7931[47]; // @[Bitwise.scala 50:65:@8024.4]
  assign _T_7980 = _T_7931[48]; // @[Bitwise.scala 50:65:@8025.4]
  assign _T_7981 = _T_7931[49]; // @[Bitwise.scala 50:65:@8026.4]
  assign _T_7982 = _T_7931[50]; // @[Bitwise.scala 50:65:@8027.4]
  assign _T_7983 = _T_7933 + _T_7934; // @[Bitwise.scala 48:55:@8028.4]
  assign _GEN_906 = {{1'd0}, _T_7932}; // @[Bitwise.scala 48:55:@8029.4]
  assign _T_7984 = _GEN_906 + _T_7983; // @[Bitwise.scala 48:55:@8029.4]
  assign _T_7985 = _T_7936 + _T_7937; // @[Bitwise.scala 48:55:@8030.4]
  assign _GEN_907 = {{1'd0}, _T_7935}; // @[Bitwise.scala 48:55:@8031.4]
  assign _T_7986 = _GEN_907 + _T_7985; // @[Bitwise.scala 48:55:@8031.4]
  assign _T_7987 = _T_7984 + _T_7986; // @[Bitwise.scala 48:55:@8032.4]
  assign _T_7988 = _T_7939 + _T_7940; // @[Bitwise.scala 48:55:@8033.4]
  assign _GEN_908 = {{1'd0}, _T_7938}; // @[Bitwise.scala 48:55:@8034.4]
  assign _T_7989 = _GEN_908 + _T_7988; // @[Bitwise.scala 48:55:@8034.4]
  assign _T_7990 = _T_7942 + _T_7943; // @[Bitwise.scala 48:55:@8035.4]
  assign _GEN_909 = {{1'd0}, _T_7941}; // @[Bitwise.scala 48:55:@8036.4]
  assign _T_7991 = _GEN_909 + _T_7990; // @[Bitwise.scala 48:55:@8036.4]
  assign _T_7992 = _T_7989 + _T_7991; // @[Bitwise.scala 48:55:@8037.4]
  assign _T_7993 = _T_7987 + _T_7992; // @[Bitwise.scala 48:55:@8038.4]
  assign _T_7994 = _T_7945 + _T_7946; // @[Bitwise.scala 48:55:@8039.4]
  assign _GEN_910 = {{1'd0}, _T_7944}; // @[Bitwise.scala 48:55:@8040.4]
  assign _T_7995 = _GEN_910 + _T_7994; // @[Bitwise.scala 48:55:@8040.4]
  assign _T_7996 = _T_7948 + _T_7949; // @[Bitwise.scala 48:55:@8041.4]
  assign _GEN_911 = {{1'd0}, _T_7947}; // @[Bitwise.scala 48:55:@8042.4]
  assign _T_7997 = _GEN_911 + _T_7996; // @[Bitwise.scala 48:55:@8042.4]
  assign _T_7998 = _T_7995 + _T_7997; // @[Bitwise.scala 48:55:@8043.4]
  assign _T_7999 = _T_7951 + _T_7952; // @[Bitwise.scala 48:55:@8044.4]
  assign _GEN_912 = {{1'd0}, _T_7950}; // @[Bitwise.scala 48:55:@8045.4]
  assign _T_8000 = _GEN_912 + _T_7999; // @[Bitwise.scala 48:55:@8045.4]
  assign _T_8001 = _T_7953 + _T_7954; // @[Bitwise.scala 48:55:@8046.4]
  assign _T_8002 = _T_7955 + _T_7956; // @[Bitwise.scala 48:55:@8047.4]
  assign _T_8003 = _T_8001 + _T_8002; // @[Bitwise.scala 48:55:@8048.4]
  assign _T_8004 = _T_8000 + _T_8003; // @[Bitwise.scala 48:55:@8049.4]
  assign _T_8005 = _T_7998 + _T_8004; // @[Bitwise.scala 48:55:@8050.4]
  assign _T_8006 = _T_7993 + _T_8005; // @[Bitwise.scala 48:55:@8051.4]
  assign _T_8007 = _T_7958 + _T_7959; // @[Bitwise.scala 48:55:@8052.4]
  assign _GEN_913 = {{1'd0}, _T_7957}; // @[Bitwise.scala 48:55:@8053.4]
  assign _T_8008 = _GEN_913 + _T_8007; // @[Bitwise.scala 48:55:@8053.4]
  assign _T_8009 = _T_7961 + _T_7962; // @[Bitwise.scala 48:55:@8054.4]
  assign _GEN_914 = {{1'd0}, _T_7960}; // @[Bitwise.scala 48:55:@8055.4]
  assign _T_8010 = _GEN_914 + _T_8009; // @[Bitwise.scala 48:55:@8055.4]
  assign _T_8011 = _T_8008 + _T_8010; // @[Bitwise.scala 48:55:@8056.4]
  assign _T_8012 = _T_7964 + _T_7965; // @[Bitwise.scala 48:55:@8057.4]
  assign _GEN_915 = {{1'd0}, _T_7963}; // @[Bitwise.scala 48:55:@8058.4]
  assign _T_8013 = _GEN_915 + _T_8012; // @[Bitwise.scala 48:55:@8058.4]
  assign _T_8014 = _T_7966 + _T_7967; // @[Bitwise.scala 48:55:@8059.4]
  assign _T_8015 = _T_7968 + _T_7969; // @[Bitwise.scala 48:55:@8060.4]
  assign _T_8016 = _T_8014 + _T_8015; // @[Bitwise.scala 48:55:@8061.4]
  assign _T_8017 = _T_8013 + _T_8016; // @[Bitwise.scala 48:55:@8062.4]
  assign _T_8018 = _T_8011 + _T_8017; // @[Bitwise.scala 48:55:@8063.4]
  assign _T_8019 = _T_7971 + _T_7972; // @[Bitwise.scala 48:55:@8064.4]
  assign _GEN_916 = {{1'd0}, _T_7970}; // @[Bitwise.scala 48:55:@8065.4]
  assign _T_8020 = _GEN_916 + _T_8019; // @[Bitwise.scala 48:55:@8065.4]
  assign _T_8021 = _T_7974 + _T_7975; // @[Bitwise.scala 48:55:@8066.4]
  assign _GEN_917 = {{1'd0}, _T_7973}; // @[Bitwise.scala 48:55:@8067.4]
  assign _T_8022 = _GEN_917 + _T_8021; // @[Bitwise.scala 48:55:@8067.4]
  assign _T_8023 = _T_8020 + _T_8022; // @[Bitwise.scala 48:55:@8068.4]
  assign _T_8024 = _T_7977 + _T_7978; // @[Bitwise.scala 48:55:@8069.4]
  assign _GEN_918 = {{1'd0}, _T_7976}; // @[Bitwise.scala 48:55:@8070.4]
  assign _T_8025 = _GEN_918 + _T_8024; // @[Bitwise.scala 48:55:@8070.4]
  assign _T_8026 = _T_7979 + _T_7980; // @[Bitwise.scala 48:55:@8071.4]
  assign _T_8027 = _T_7981 + _T_7982; // @[Bitwise.scala 48:55:@8072.4]
  assign _T_8028 = _T_8026 + _T_8027; // @[Bitwise.scala 48:55:@8073.4]
  assign _T_8029 = _T_8025 + _T_8028; // @[Bitwise.scala 48:55:@8074.4]
  assign _T_8030 = _T_8023 + _T_8029; // @[Bitwise.scala 48:55:@8075.4]
  assign _T_8031 = _T_8018 + _T_8030; // @[Bitwise.scala 48:55:@8076.4]
  assign _T_8032 = _T_8006 + _T_8031; // @[Bitwise.scala 48:55:@8077.4]
  assign _T_8096 = _T_2230[51:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@8142.4]
  assign _T_8097 = _T_8096[0]; // @[Bitwise.scala 50:65:@8143.4]
  assign _T_8098 = _T_8096[1]; // @[Bitwise.scala 50:65:@8144.4]
  assign _T_8099 = _T_8096[2]; // @[Bitwise.scala 50:65:@8145.4]
  assign _T_8100 = _T_8096[3]; // @[Bitwise.scala 50:65:@8146.4]
  assign _T_8101 = _T_8096[4]; // @[Bitwise.scala 50:65:@8147.4]
  assign _T_8102 = _T_8096[5]; // @[Bitwise.scala 50:65:@8148.4]
  assign _T_8103 = _T_8096[6]; // @[Bitwise.scala 50:65:@8149.4]
  assign _T_8104 = _T_8096[7]; // @[Bitwise.scala 50:65:@8150.4]
  assign _T_8105 = _T_8096[8]; // @[Bitwise.scala 50:65:@8151.4]
  assign _T_8106 = _T_8096[9]; // @[Bitwise.scala 50:65:@8152.4]
  assign _T_8107 = _T_8096[10]; // @[Bitwise.scala 50:65:@8153.4]
  assign _T_8108 = _T_8096[11]; // @[Bitwise.scala 50:65:@8154.4]
  assign _T_8109 = _T_8096[12]; // @[Bitwise.scala 50:65:@8155.4]
  assign _T_8110 = _T_8096[13]; // @[Bitwise.scala 50:65:@8156.4]
  assign _T_8111 = _T_8096[14]; // @[Bitwise.scala 50:65:@8157.4]
  assign _T_8112 = _T_8096[15]; // @[Bitwise.scala 50:65:@8158.4]
  assign _T_8113 = _T_8096[16]; // @[Bitwise.scala 50:65:@8159.4]
  assign _T_8114 = _T_8096[17]; // @[Bitwise.scala 50:65:@8160.4]
  assign _T_8115 = _T_8096[18]; // @[Bitwise.scala 50:65:@8161.4]
  assign _T_8116 = _T_8096[19]; // @[Bitwise.scala 50:65:@8162.4]
  assign _T_8117 = _T_8096[20]; // @[Bitwise.scala 50:65:@8163.4]
  assign _T_8118 = _T_8096[21]; // @[Bitwise.scala 50:65:@8164.4]
  assign _T_8119 = _T_8096[22]; // @[Bitwise.scala 50:65:@8165.4]
  assign _T_8120 = _T_8096[23]; // @[Bitwise.scala 50:65:@8166.4]
  assign _T_8121 = _T_8096[24]; // @[Bitwise.scala 50:65:@8167.4]
  assign _T_8122 = _T_8096[25]; // @[Bitwise.scala 50:65:@8168.4]
  assign _T_8123 = _T_8096[26]; // @[Bitwise.scala 50:65:@8169.4]
  assign _T_8124 = _T_8096[27]; // @[Bitwise.scala 50:65:@8170.4]
  assign _T_8125 = _T_8096[28]; // @[Bitwise.scala 50:65:@8171.4]
  assign _T_8126 = _T_8096[29]; // @[Bitwise.scala 50:65:@8172.4]
  assign _T_8127 = _T_8096[30]; // @[Bitwise.scala 50:65:@8173.4]
  assign _T_8128 = _T_8096[31]; // @[Bitwise.scala 50:65:@8174.4]
  assign _T_8129 = _T_8096[32]; // @[Bitwise.scala 50:65:@8175.4]
  assign _T_8130 = _T_8096[33]; // @[Bitwise.scala 50:65:@8176.4]
  assign _T_8131 = _T_8096[34]; // @[Bitwise.scala 50:65:@8177.4]
  assign _T_8132 = _T_8096[35]; // @[Bitwise.scala 50:65:@8178.4]
  assign _T_8133 = _T_8096[36]; // @[Bitwise.scala 50:65:@8179.4]
  assign _T_8134 = _T_8096[37]; // @[Bitwise.scala 50:65:@8180.4]
  assign _T_8135 = _T_8096[38]; // @[Bitwise.scala 50:65:@8181.4]
  assign _T_8136 = _T_8096[39]; // @[Bitwise.scala 50:65:@8182.4]
  assign _T_8137 = _T_8096[40]; // @[Bitwise.scala 50:65:@8183.4]
  assign _T_8138 = _T_8096[41]; // @[Bitwise.scala 50:65:@8184.4]
  assign _T_8139 = _T_8096[42]; // @[Bitwise.scala 50:65:@8185.4]
  assign _T_8140 = _T_8096[43]; // @[Bitwise.scala 50:65:@8186.4]
  assign _T_8141 = _T_8096[44]; // @[Bitwise.scala 50:65:@8187.4]
  assign _T_8142 = _T_8096[45]; // @[Bitwise.scala 50:65:@8188.4]
  assign _T_8143 = _T_8096[46]; // @[Bitwise.scala 50:65:@8189.4]
  assign _T_8144 = _T_8096[47]; // @[Bitwise.scala 50:65:@8190.4]
  assign _T_8145 = _T_8096[48]; // @[Bitwise.scala 50:65:@8191.4]
  assign _T_8146 = _T_8096[49]; // @[Bitwise.scala 50:65:@8192.4]
  assign _T_8147 = _T_8096[50]; // @[Bitwise.scala 50:65:@8193.4]
  assign _T_8148 = _T_8096[51]; // @[Bitwise.scala 50:65:@8194.4]
  assign _T_8149 = _T_8098 + _T_8099; // @[Bitwise.scala 48:55:@8195.4]
  assign _GEN_919 = {{1'd0}, _T_8097}; // @[Bitwise.scala 48:55:@8196.4]
  assign _T_8150 = _GEN_919 + _T_8149; // @[Bitwise.scala 48:55:@8196.4]
  assign _T_8151 = _T_8101 + _T_8102; // @[Bitwise.scala 48:55:@8197.4]
  assign _GEN_920 = {{1'd0}, _T_8100}; // @[Bitwise.scala 48:55:@8198.4]
  assign _T_8152 = _GEN_920 + _T_8151; // @[Bitwise.scala 48:55:@8198.4]
  assign _T_8153 = _T_8150 + _T_8152; // @[Bitwise.scala 48:55:@8199.4]
  assign _T_8154 = _T_8104 + _T_8105; // @[Bitwise.scala 48:55:@8200.4]
  assign _GEN_921 = {{1'd0}, _T_8103}; // @[Bitwise.scala 48:55:@8201.4]
  assign _T_8155 = _GEN_921 + _T_8154; // @[Bitwise.scala 48:55:@8201.4]
  assign _T_8156 = _T_8106 + _T_8107; // @[Bitwise.scala 48:55:@8202.4]
  assign _T_8157 = _T_8108 + _T_8109; // @[Bitwise.scala 48:55:@8203.4]
  assign _T_8158 = _T_8156 + _T_8157; // @[Bitwise.scala 48:55:@8204.4]
  assign _T_8159 = _T_8155 + _T_8158; // @[Bitwise.scala 48:55:@8205.4]
  assign _T_8160 = _T_8153 + _T_8159; // @[Bitwise.scala 48:55:@8206.4]
  assign _T_8161 = _T_8111 + _T_8112; // @[Bitwise.scala 48:55:@8207.4]
  assign _GEN_922 = {{1'd0}, _T_8110}; // @[Bitwise.scala 48:55:@8208.4]
  assign _T_8162 = _GEN_922 + _T_8161; // @[Bitwise.scala 48:55:@8208.4]
  assign _T_8163 = _T_8114 + _T_8115; // @[Bitwise.scala 48:55:@8209.4]
  assign _GEN_923 = {{1'd0}, _T_8113}; // @[Bitwise.scala 48:55:@8210.4]
  assign _T_8164 = _GEN_923 + _T_8163; // @[Bitwise.scala 48:55:@8210.4]
  assign _T_8165 = _T_8162 + _T_8164; // @[Bitwise.scala 48:55:@8211.4]
  assign _T_8166 = _T_8117 + _T_8118; // @[Bitwise.scala 48:55:@8212.4]
  assign _GEN_924 = {{1'd0}, _T_8116}; // @[Bitwise.scala 48:55:@8213.4]
  assign _T_8167 = _GEN_924 + _T_8166; // @[Bitwise.scala 48:55:@8213.4]
  assign _T_8168 = _T_8119 + _T_8120; // @[Bitwise.scala 48:55:@8214.4]
  assign _T_8169 = _T_8121 + _T_8122; // @[Bitwise.scala 48:55:@8215.4]
  assign _T_8170 = _T_8168 + _T_8169; // @[Bitwise.scala 48:55:@8216.4]
  assign _T_8171 = _T_8167 + _T_8170; // @[Bitwise.scala 48:55:@8217.4]
  assign _T_8172 = _T_8165 + _T_8171; // @[Bitwise.scala 48:55:@8218.4]
  assign _T_8173 = _T_8160 + _T_8172; // @[Bitwise.scala 48:55:@8219.4]
  assign _T_8174 = _T_8124 + _T_8125; // @[Bitwise.scala 48:55:@8220.4]
  assign _GEN_925 = {{1'd0}, _T_8123}; // @[Bitwise.scala 48:55:@8221.4]
  assign _T_8175 = _GEN_925 + _T_8174; // @[Bitwise.scala 48:55:@8221.4]
  assign _T_8176 = _T_8127 + _T_8128; // @[Bitwise.scala 48:55:@8222.4]
  assign _GEN_926 = {{1'd0}, _T_8126}; // @[Bitwise.scala 48:55:@8223.4]
  assign _T_8177 = _GEN_926 + _T_8176; // @[Bitwise.scala 48:55:@8223.4]
  assign _T_8178 = _T_8175 + _T_8177; // @[Bitwise.scala 48:55:@8224.4]
  assign _T_8179 = _T_8130 + _T_8131; // @[Bitwise.scala 48:55:@8225.4]
  assign _GEN_927 = {{1'd0}, _T_8129}; // @[Bitwise.scala 48:55:@8226.4]
  assign _T_8180 = _GEN_927 + _T_8179; // @[Bitwise.scala 48:55:@8226.4]
  assign _T_8181 = _T_8132 + _T_8133; // @[Bitwise.scala 48:55:@8227.4]
  assign _T_8182 = _T_8134 + _T_8135; // @[Bitwise.scala 48:55:@8228.4]
  assign _T_8183 = _T_8181 + _T_8182; // @[Bitwise.scala 48:55:@8229.4]
  assign _T_8184 = _T_8180 + _T_8183; // @[Bitwise.scala 48:55:@8230.4]
  assign _T_8185 = _T_8178 + _T_8184; // @[Bitwise.scala 48:55:@8231.4]
  assign _T_8186 = _T_8137 + _T_8138; // @[Bitwise.scala 48:55:@8232.4]
  assign _GEN_928 = {{1'd0}, _T_8136}; // @[Bitwise.scala 48:55:@8233.4]
  assign _T_8187 = _GEN_928 + _T_8186; // @[Bitwise.scala 48:55:@8233.4]
  assign _T_8188 = _T_8140 + _T_8141; // @[Bitwise.scala 48:55:@8234.4]
  assign _GEN_929 = {{1'd0}, _T_8139}; // @[Bitwise.scala 48:55:@8235.4]
  assign _T_8189 = _GEN_929 + _T_8188; // @[Bitwise.scala 48:55:@8235.4]
  assign _T_8190 = _T_8187 + _T_8189; // @[Bitwise.scala 48:55:@8236.4]
  assign _T_8191 = _T_8143 + _T_8144; // @[Bitwise.scala 48:55:@8237.4]
  assign _GEN_930 = {{1'd0}, _T_8142}; // @[Bitwise.scala 48:55:@8238.4]
  assign _T_8192 = _GEN_930 + _T_8191; // @[Bitwise.scala 48:55:@8238.4]
  assign _T_8193 = _T_8145 + _T_8146; // @[Bitwise.scala 48:55:@8239.4]
  assign _T_8194 = _T_8147 + _T_8148; // @[Bitwise.scala 48:55:@8240.4]
  assign _T_8195 = _T_8193 + _T_8194; // @[Bitwise.scala 48:55:@8241.4]
  assign _T_8196 = _T_8192 + _T_8195; // @[Bitwise.scala 48:55:@8242.4]
  assign _T_8197 = _T_8190 + _T_8196; // @[Bitwise.scala 48:55:@8243.4]
  assign _T_8198 = _T_8185 + _T_8197; // @[Bitwise.scala 48:55:@8244.4]
  assign _T_8199 = _T_8173 + _T_8198; // @[Bitwise.scala 48:55:@8245.4]
  assign _T_8263 = _T_2230[52:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@8310.4]
  assign _T_8264 = _T_8263[0]; // @[Bitwise.scala 50:65:@8311.4]
  assign _T_8265 = _T_8263[1]; // @[Bitwise.scala 50:65:@8312.4]
  assign _T_8266 = _T_8263[2]; // @[Bitwise.scala 50:65:@8313.4]
  assign _T_8267 = _T_8263[3]; // @[Bitwise.scala 50:65:@8314.4]
  assign _T_8268 = _T_8263[4]; // @[Bitwise.scala 50:65:@8315.4]
  assign _T_8269 = _T_8263[5]; // @[Bitwise.scala 50:65:@8316.4]
  assign _T_8270 = _T_8263[6]; // @[Bitwise.scala 50:65:@8317.4]
  assign _T_8271 = _T_8263[7]; // @[Bitwise.scala 50:65:@8318.4]
  assign _T_8272 = _T_8263[8]; // @[Bitwise.scala 50:65:@8319.4]
  assign _T_8273 = _T_8263[9]; // @[Bitwise.scala 50:65:@8320.4]
  assign _T_8274 = _T_8263[10]; // @[Bitwise.scala 50:65:@8321.4]
  assign _T_8275 = _T_8263[11]; // @[Bitwise.scala 50:65:@8322.4]
  assign _T_8276 = _T_8263[12]; // @[Bitwise.scala 50:65:@8323.4]
  assign _T_8277 = _T_8263[13]; // @[Bitwise.scala 50:65:@8324.4]
  assign _T_8278 = _T_8263[14]; // @[Bitwise.scala 50:65:@8325.4]
  assign _T_8279 = _T_8263[15]; // @[Bitwise.scala 50:65:@8326.4]
  assign _T_8280 = _T_8263[16]; // @[Bitwise.scala 50:65:@8327.4]
  assign _T_8281 = _T_8263[17]; // @[Bitwise.scala 50:65:@8328.4]
  assign _T_8282 = _T_8263[18]; // @[Bitwise.scala 50:65:@8329.4]
  assign _T_8283 = _T_8263[19]; // @[Bitwise.scala 50:65:@8330.4]
  assign _T_8284 = _T_8263[20]; // @[Bitwise.scala 50:65:@8331.4]
  assign _T_8285 = _T_8263[21]; // @[Bitwise.scala 50:65:@8332.4]
  assign _T_8286 = _T_8263[22]; // @[Bitwise.scala 50:65:@8333.4]
  assign _T_8287 = _T_8263[23]; // @[Bitwise.scala 50:65:@8334.4]
  assign _T_8288 = _T_8263[24]; // @[Bitwise.scala 50:65:@8335.4]
  assign _T_8289 = _T_8263[25]; // @[Bitwise.scala 50:65:@8336.4]
  assign _T_8290 = _T_8263[26]; // @[Bitwise.scala 50:65:@8337.4]
  assign _T_8291 = _T_8263[27]; // @[Bitwise.scala 50:65:@8338.4]
  assign _T_8292 = _T_8263[28]; // @[Bitwise.scala 50:65:@8339.4]
  assign _T_8293 = _T_8263[29]; // @[Bitwise.scala 50:65:@8340.4]
  assign _T_8294 = _T_8263[30]; // @[Bitwise.scala 50:65:@8341.4]
  assign _T_8295 = _T_8263[31]; // @[Bitwise.scala 50:65:@8342.4]
  assign _T_8296 = _T_8263[32]; // @[Bitwise.scala 50:65:@8343.4]
  assign _T_8297 = _T_8263[33]; // @[Bitwise.scala 50:65:@8344.4]
  assign _T_8298 = _T_8263[34]; // @[Bitwise.scala 50:65:@8345.4]
  assign _T_8299 = _T_8263[35]; // @[Bitwise.scala 50:65:@8346.4]
  assign _T_8300 = _T_8263[36]; // @[Bitwise.scala 50:65:@8347.4]
  assign _T_8301 = _T_8263[37]; // @[Bitwise.scala 50:65:@8348.4]
  assign _T_8302 = _T_8263[38]; // @[Bitwise.scala 50:65:@8349.4]
  assign _T_8303 = _T_8263[39]; // @[Bitwise.scala 50:65:@8350.4]
  assign _T_8304 = _T_8263[40]; // @[Bitwise.scala 50:65:@8351.4]
  assign _T_8305 = _T_8263[41]; // @[Bitwise.scala 50:65:@8352.4]
  assign _T_8306 = _T_8263[42]; // @[Bitwise.scala 50:65:@8353.4]
  assign _T_8307 = _T_8263[43]; // @[Bitwise.scala 50:65:@8354.4]
  assign _T_8308 = _T_8263[44]; // @[Bitwise.scala 50:65:@8355.4]
  assign _T_8309 = _T_8263[45]; // @[Bitwise.scala 50:65:@8356.4]
  assign _T_8310 = _T_8263[46]; // @[Bitwise.scala 50:65:@8357.4]
  assign _T_8311 = _T_8263[47]; // @[Bitwise.scala 50:65:@8358.4]
  assign _T_8312 = _T_8263[48]; // @[Bitwise.scala 50:65:@8359.4]
  assign _T_8313 = _T_8263[49]; // @[Bitwise.scala 50:65:@8360.4]
  assign _T_8314 = _T_8263[50]; // @[Bitwise.scala 50:65:@8361.4]
  assign _T_8315 = _T_8263[51]; // @[Bitwise.scala 50:65:@8362.4]
  assign _T_8316 = _T_8263[52]; // @[Bitwise.scala 50:65:@8363.4]
  assign _T_8317 = _T_8265 + _T_8266; // @[Bitwise.scala 48:55:@8364.4]
  assign _GEN_931 = {{1'd0}, _T_8264}; // @[Bitwise.scala 48:55:@8365.4]
  assign _T_8318 = _GEN_931 + _T_8317; // @[Bitwise.scala 48:55:@8365.4]
  assign _T_8319 = _T_8268 + _T_8269; // @[Bitwise.scala 48:55:@8366.4]
  assign _GEN_932 = {{1'd0}, _T_8267}; // @[Bitwise.scala 48:55:@8367.4]
  assign _T_8320 = _GEN_932 + _T_8319; // @[Bitwise.scala 48:55:@8367.4]
  assign _T_8321 = _T_8318 + _T_8320; // @[Bitwise.scala 48:55:@8368.4]
  assign _T_8322 = _T_8271 + _T_8272; // @[Bitwise.scala 48:55:@8369.4]
  assign _GEN_933 = {{1'd0}, _T_8270}; // @[Bitwise.scala 48:55:@8370.4]
  assign _T_8323 = _GEN_933 + _T_8322; // @[Bitwise.scala 48:55:@8370.4]
  assign _T_8324 = _T_8273 + _T_8274; // @[Bitwise.scala 48:55:@8371.4]
  assign _T_8325 = _T_8275 + _T_8276; // @[Bitwise.scala 48:55:@8372.4]
  assign _T_8326 = _T_8324 + _T_8325; // @[Bitwise.scala 48:55:@8373.4]
  assign _T_8327 = _T_8323 + _T_8326; // @[Bitwise.scala 48:55:@8374.4]
  assign _T_8328 = _T_8321 + _T_8327; // @[Bitwise.scala 48:55:@8375.4]
  assign _T_8329 = _T_8278 + _T_8279; // @[Bitwise.scala 48:55:@8376.4]
  assign _GEN_934 = {{1'd0}, _T_8277}; // @[Bitwise.scala 48:55:@8377.4]
  assign _T_8330 = _GEN_934 + _T_8329; // @[Bitwise.scala 48:55:@8377.4]
  assign _T_8331 = _T_8281 + _T_8282; // @[Bitwise.scala 48:55:@8378.4]
  assign _GEN_935 = {{1'd0}, _T_8280}; // @[Bitwise.scala 48:55:@8379.4]
  assign _T_8332 = _GEN_935 + _T_8331; // @[Bitwise.scala 48:55:@8379.4]
  assign _T_8333 = _T_8330 + _T_8332; // @[Bitwise.scala 48:55:@8380.4]
  assign _T_8334 = _T_8284 + _T_8285; // @[Bitwise.scala 48:55:@8381.4]
  assign _GEN_936 = {{1'd0}, _T_8283}; // @[Bitwise.scala 48:55:@8382.4]
  assign _T_8335 = _GEN_936 + _T_8334; // @[Bitwise.scala 48:55:@8382.4]
  assign _T_8336 = _T_8286 + _T_8287; // @[Bitwise.scala 48:55:@8383.4]
  assign _T_8337 = _T_8288 + _T_8289; // @[Bitwise.scala 48:55:@8384.4]
  assign _T_8338 = _T_8336 + _T_8337; // @[Bitwise.scala 48:55:@8385.4]
  assign _T_8339 = _T_8335 + _T_8338; // @[Bitwise.scala 48:55:@8386.4]
  assign _T_8340 = _T_8333 + _T_8339; // @[Bitwise.scala 48:55:@8387.4]
  assign _T_8341 = _T_8328 + _T_8340; // @[Bitwise.scala 48:55:@8388.4]
  assign _T_8342 = _T_8291 + _T_8292; // @[Bitwise.scala 48:55:@8389.4]
  assign _GEN_937 = {{1'd0}, _T_8290}; // @[Bitwise.scala 48:55:@8390.4]
  assign _T_8343 = _GEN_937 + _T_8342; // @[Bitwise.scala 48:55:@8390.4]
  assign _T_8344 = _T_8294 + _T_8295; // @[Bitwise.scala 48:55:@8391.4]
  assign _GEN_938 = {{1'd0}, _T_8293}; // @[Bitwise.scala 48:55:@8392.4]
  assign _T_8345 = _GEN_938 + _T_8344; // @[Bitwise.scala 48:55:@8392.4]
  assign _T_8346 = _T_8343 + _T_8345; // @[Bitwise.scala 48:55:@8393.4]
  assign _T_8347 = _T_8297 + _T_8298; // @[Bitwise.scala 48:55:@8394.4]
  assign _GEN_939 = {{1'd0}, _T_8296}; // @[Bitwise.scala 48:55:@8395.4]
  assign _T_8348 = _GEN_939 + _T_8347; // @[Bitwise.scala 48:55:@8395.4]
  assign _T_8349 = _T_8299 + _T_8300; // @[Bitwise.scala 48:55:@8396.4]
  assign _T_8350 = _T_8301 + _T_8302; // @[Bitwise.scala 48:55:@8397.4]
  assign _T_8351 = _T_8349 + _T_8350; // @[Bitwise.scala 48:55:@8398.4]
  assign _T_8352 = _T_8348 + _T_8351; // @[Bitwise.scala 48:55:@8399.4]
  assign _T_8353 = _T_8346 + _T_8352; // @[Bitwise.scala 48:55:@8400.4]
  assign _T_8354 = _T_8304 + _T_8305; // @[Bitwise.scala 48:55:@8401.4]
  assign _GEN_940 = {{1'd0}, _T_8303}; // @[Bitwise.scala 48:55:@8402.4]
  assign _T_8355 = _GEN_940 + _T_8354; // @[Bitwise.scala 48:55:@8402.4]
  assign _T_8356 = _T_8306 + _T_8307; // @[Bitwise.scala 48:55:@8403.4]
  assign _T_8357 = _T_8308 + _T_8309; // @[Bitwise.scala 48:55:@8404.4]
  assign _T_8358 = _T_8356 + _T_8357; // @[Bitwise.scala 48:55:@8405.4]
  assign _T_8359 = _T_8355 + _T_8358; // @[Bitwise.scala 48:55:@8406.4]
  assign _T_8360 = _T_8311 + _T_8312; // @[Bitwise.scala 48:55:@8407.4]
  assign _GEN_941 = {{1'd0}, _T_8310}; // @[Bitwise.scala 48:55:@8408.4]
  assign _T_8361 = _GEN_941 + _T_8360; // @[Bitwise.scala 48:55:@8408.4]
  assign _T_8362 = _T_8313 + _T_8314; // @[Bitwise.scala 48:55:@8409.4]
  assign _T_8363 = _T_8315 + _T_8316; // @[Bitwise.scala 48:55:@8410.4]
  assign _T_8364 = _T_8362 + _T_8363; // @[Bitwise.scala 48:55:@8411.4]
  assign _T_8365 = _T_8361 + _T_8364; // @[Bitwise.scala 48:55:@8412.4]
  assign _T_8366 = _T_8359 + _T_8365; // @[Bitwise.scala 48:55:@8413.4]
  assign _T_8367 = _T_8353 + _T_8366; // @[Bitwise.scala 48:55:@8414.4]
  assign _T_8368 = _T_8341 + _T_8367; // @[Bitwise.scala 48:55:@8415.4]
  assign _T_8432 = _T_2230[53:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@8480.4]
  assign _T_8433 = _T_8432[0]; // @[Bitwise.scala 50:65:@8481.4]
  assign _T_8434 = _T_8432[1]; // @[Bitwise.scala 50:65:@8482.4]
  assign _T_8435 = _T_8432[2]; // @[Bitwise.scala 50:65:@8483.4]
  assign _T_8436 = _T_8432[3]; // @[Bitwise.scala 50:65:@8484.4]
  assign _T_8437 = _T_8432[4]; // @[Bitwise.scala 50:65:@8485.4]
  assign _T_8438 = _T_8432[5]; // @[Bitwise.scala 50:65:@8486.4]
  assign _T_8439 = _T_8432[6]; // @[Bitwise.scala 50:65:@8487.4]
  assign _T_8440 = _T_8432[7]; // @[Bitwise.scala 50:65:@8488.4]
  assign _T_8441 = _T_8432[8]; // @[Bitwise.scala 50:65:@8489.4]
  assign _T_8442 = _T_8432[9]; // @[Bitwise.scala 50:65:@8490.4]
  assign _T_8443 = _T_8432[10]; // @[Bitwise.scala 50:65:@8491.4]
  assign _T_8444 = _T_8432[11]; // @[Bitwise.scala 50:65:@8492.4]
  assign _T_8445 = _T_8432[12]; // @[Bitwise.scala 50:65:@8493.4]
  assign _T_8446 = _T_8432[13]; // @[Bitwise.scala 50:65:@8494.4]
  assign _T_8447 = _T_8432[14]; // @[Bitwise.scala 50:65:@8495.4]
  assign _T_8448 = _T_8432[15]; // @[Bitwise.scala 50:65:@8496.4]
  assign _T_8449 = _T_8432[16]; // @[Bitwise.scala 50:65:@8497.4]
  assign _T_8450 = _T_8432[17]; // @[Bitwise.scala 50:65:@8498.4]
  assign _T_8451 = _T_8432[18]; // @[Bitwise.scala 50:65:@8499.4]
  assign _T_8452 = _T_8432[19]; // @[Bitwise.scala 50:65:@8500.4]
  assign _T_8453 = _T_8432[20]; // @[Bitwise.scala 50:65:@8501.4]
  assign _T_8454 = _T_8432[21]; // @[Bitwise.scala 50:65:@8502.4]
  assign _T_8455 = _T_8432[22]; // @[Bitwise.scala 50:65:@8503.4]
  assign _T_8456 = _T_8432[23]; // @[Bitwise.scala 50:65:@8504.4]
  assign _T_8457 = _T_8432[24]; // @[Bitwise.scala 50:65:@8505.4]
  assign _T_8458 = _T_8432[25]; // @[Bitwise.scala 50:65:@8506.4]
  assign _T_8459 = _T_8432[26]; // @[Bitwise.scala 50:65:@8507.4]
  assign _T_8460 = _T_8432[27]; // @[Bitwise.scala 50:65:@8508.4]
  assign _T_8461 = _T_8432[28]; // @[Bitwise.scala 50:65:@8509.4]
  assign _T_8462 = _T_8432[29]; // @[Bitwise.scala 50:65:@8510.4]
  assign _T_8463 = _T_8432[30]; // @[Bitwise.scala 50:65:@8511.4]
  assign _T_8464 = _T_8432[31]; // @[Bitwise.scala 50:65:@8512.4]
  assign _T_8465 = _T_8432[32]; // @[Bitwise.scala 50:65:@8513.4]
  assign _T_8466 = _T_8432[33]; // @[Bitwise.scala 50:65:@8514.4]
  assign _T_8467 = _T_8432[34]; // @[Bitwise.scala 50:65:@8515.4]
  assign _T_8468 = _T_8432[35]; // @[Bitwise.scala 50:65:@8516.4]
  assign _T_8469 = _T_8432[36]; // @[Bitwise.scala 50:65:@8517.4]
  assign _T_8470 = _T_8432[37]; // @[Bitwise.scala 50:65:@8518.4]
  assign _T_8471 = _T_8432[38]; // @[Bitwise.scala 50:65:@8519.4]
  assign _T_8472 = _T_8432[39]; // @[Bitwise.scala 50:65:@8520.4]
  assign _T_8473 = _T_8432[40]; // @[Bitwise.scala 50:65:@8521.4]
  assign _T_8474 = _T_8432[41]; // @[Bitwise.scala 50:65:@8522.4]
  assign _T_8475 = _T_8432[42]; // @[Bitwise.scala 50:65:@8523.4]
  assign _T_8476 = _T_8432[43]; // @[Bitwise.scala 50:65:@8524.4]
  assign _T_8477 = _T_8432[44]; // @[Bitwise.scala 50:65:@8525.4]
  assign _T_8478 = _T_8432[45]; // @[Bitwise.scala 50:65:@8526.4]
  assign _T_8479 = _T_8432[46]; // @[Bitwise.scala 50:65:@8527.4]
  assign _T_8480 = _T_8432[47]; // @[Bitwise.scala 50:65:@8528.4]
  assign _T_8481 = _T_8432[48]; // @[Bitwise.scala 50:65:@8529.4]
  assign _T_8482 = _T_8432[49]; // @[Bitwise.scala 50:65:@8530.4]
  assign _T_8483 = _T_8432[50]; // @[Bitwise.scala 50:65:@8531.4]
  assign _T_8484 = _T_8432[51]; // @[Bitwise.scala 50:65:@8532.4]
  assign _T_8485 = _T_8432[52]; // @[Bitwise.scala 50:65:@8533.4]
  assign _T_8486 = _T_8432[53]; // @[Bitwise.scala 50:65:@8534.4]
  assign _T_8487 = _T_8434 + _T_8435; // @[Bitwise.scala 48:55:@8535.4]
  assign _GEN_942 = {{1'd0}, _T_8433}; // @[Bitwise.scala 48:55:@8536.4]
  assign _T_8488 = _GEN_942 + _T_8487; // @[Bitwise.scala 48:55:@8536.4]
  assign _T_8489 = _T_8437 + _T_8438; // @[Bitwise.scala 48:55:@8537.4]
  assign _GEN_943 = {{1'd0}, _T_8436}; // @[Bitwise.scala 48:55:@8538.4]
  assign _T_8490 = _GEN_943 + _T_8489; // @[Bitwise.scala 48:55:@8538.4]
  assign _T_8491 = _T_8488 + _T_8490; // @[Bitwise.scala 48:55:@8539.4]
  assign _T_8492 = _T_8440 + _T_8441; // @[Bitwise.scala 48:55:@8540.4]
  assign _GEN_944 = {{1'd0}, _T_8439}; // @[Bitwise.scala 48:55:@8541.4]
  assign _T_8493 = _GEN_944 + _T_8492; // @[Bitwise.scala 48:55:@8541.4]
  assign _T_8494 = _T_8442 + _T_8443; // @[Bitwise.scala 48:55:@8542.4]
  assign _T_8495 = _T_8444 + _T_8445; // @[Bitwise.scala 48:55:@8543.4]
  assign _T_8496 = _T_8494 + _T_8495; // @[Bitwise.scala 48:55:@8544.4]
  assign _T_8497 = _T_8493 + _T_8496; // @[Bitwise.scala 48:55:@8545.4]
  assign _T_8498 = _T_8491 + _T_8497; // @[Bitwise.scala 48:55:@8546.4]
  assign _T_8499 = _T_8447 + _T_8448; // @[Bitwise.scala 48:55:@8547.4]
  assign _GEN_945 = {{1'd0}, _T_8446}; // @[Bitwise.scala 48:55:@8548.4]
  assign _T_8500 = _GEN_945 + _T_8499; // @[Bitwise.scala 48:55:@8548.4]
  assign _T_8501 = _T_8449 + _T_8450; // @[Bitwise.scala 48:55:@8549.4]
  assign _T_8502 = _T_8451 + _T_8452; // @[Bitwise.scala 48:55:@8550.4]
  assign _T_8503 = _T_8501 + _T_8502; // @[Bitwise.scala 48:55:@8551.4]
  assign _T_8504 = _T_8500 + _T_8503; // @[Bitwise.scala 48:55:@8552.4]
  assign _T_8505 = _T_8454 + _T_8455; // @[Bitwise.scala 48:55:@8553.4]
  assign _GEN_946 = {{1'd0}, _T_8453}; // @[Bitwise.scala 48:55:@8554.4]
  assign _T_8506 = _GEN_946 + _T_8505; // @[Bitwise.scala 48:55:@8554.4]
  assign _T_8507 = _T_8456 + _T_8457; // @[Bitwise.scala 48:55:@8555.4]
  assign _T_8508 = _T_8458 + _T_8459; // @[Bitwise.scala 48:55:@8556.4]
  assign _T_8509 = _T_8507 + _T_8508; // @[Bitwise.scala 48:55:@8557.4]
  assign _T_8510 = _T_8506 + _T_8509; // @[Bitwise.scala 48:55:@8558.4]
  assign _T_8511 = _T_8504 + _T_8510; // @[Bitwise.scala 48:55:@8559.4]
  assign _T_8512 = _T_8498 + _T_8511; // @[Bitwise.scala 48:55:@8560.4]
  assign _T_8513 = _T_8461 + _T_8462; // @[Bitwise.scala 48:55:@8561.4]
  assign _GEN_947 = {{1'd0}, _T_8460}; // @[Bitwise.scala 48:55:@8562.4]
  assign _T_8514 = _GEN_947 + _T_8513; // @[Bitwise.scala 48:55:@8562.4]
  assign _T_8515 = _T_8464 + _T_8465; // @[Bitwise.scala 48:55:@8563.4]
  assign _GEN_948 = {{1'd0}, _T_8463}; // @[Bitwise.scala 48:55:@8564.4]
  assign _T_8516 = _GEN_948 + _T_8515; // @[Bitwise.scala 48:55:@8564.4]
  assign _T_8517 = _T_8514 + _T_8516; // @[Bitwise.scala 48:55:@8565.4]
  assign _T_8518 = _T_8467 + _T_8468; // @[Bitwise.scala 48:55:@8566.4]
  assign _GEN_949 = {{1'd0}, _T_8466}; // @[Bitwise.scala 48:55:@8567.4]
  assign _T_8519 = _GEN_949 + _T_8518; // @[Bitwise.scala 48:55:@8567.4]
  assign _T_8520 = _T_8469 + _T_8470; // @[Bitwise.scala 48:55:@8568.4]
  assign _T_8521 = _T_8471 + _T_8472; // @[Bitwise.scala 48:55:@8569.4]
  assign _T_8522 = _T_8520 + _T_8521; // @[Bitwise.scala 48:55:@8570.4]
  assign _T_8523 = _T_8519 + _T_8522; // @[Bitwise.scala 48:55:@8571.4]
  assign _T_8524 = _T_8517 + _T_8523; // @[Bitwise.scala 48:55:@8572.4]
  assign _T_8525 = _T_8474 + _T_8475; // @[Bitwise.scala 48:55:@8573.4]
  assign _GEN_950 = {{1'd0}, _T_8473}; // @[Bitwise.scala 48:55:@8574.4]
  assign _T_8526 = _GEN_950 + _T_8525; // @[Bitwise.scala 48:55:@8574.4]
  assign _T_8527 = _T_8476 + _T_8477; // @[Bitwise.scala 48:55:@8575.4]
  assign _T_8528 = _T_8478 + _T_8479; // @[Bitwise.scala 48:55:@8576.4]
  assign _T_8529 = _T_8527 + _T_8528; // @[Bitwise.scala 48:55:@8577.4]
  assign _T_8530 = _T_8526 + _T_8529; // @[Bitwise.scala 48:55:@8578.4]
  assign _T_8531 = _T_8481 + _T_8482; // @[Bitwise.scala 48:55:@8579.4]
  assign _GEN_951 = {{1'd0}, _T_8480}; // @[Bitwise.scala 48:55:@8580.4]
  assign _T_8532 = _GEN_951 + _T_8531; // @[Bitwise.scala 48:55:@8580.4]
  assign _T_8533 = _T_8483 + _T_8484; // @[Bitwise.scala 48:55:@8581.4]
  assign _T_8534 = _T_8485 + _T_8486; // @[Bitwise.scala 48:55:@8582.4]
  assign _T_8535 = _T_8533 + _T_8534; // @[Bitwise.scala 48:55:@8583.4]
  assign _T_8536 = _T_8532 + _T_8535; // @[Bitwise.scala 48:55:@8584.4]
  assign _T_8537 = _T_8530 + _T_8536; // @[Bitwise.scala 48:55:@8585.4]
  assign _T_8538 = _T_8524 + _T_8537; // @[Bitwise.scala 48:55:@8586.4]
  assign _T_8539 = _T_8512 + _T_8538; // @[Bitwise.scala 48:55:@8587.4]
  assign _T_8603 = _T_2230[54:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@8652.4]
  assign _T_8604 = _T_8603[0]; // @[Bitwise.scala 50:65:@8653.4]
  assign _T_8605 = _T_8603[1]; // @[Bitwise.scala 50:65:@8654.4]
  assign _T_8606 = _T_8603[2]; // @[Bitwise.scala 50:65:@8655.4]
  assign _T_8607 = _T_8603[3]; // @[Bitwise.scala 50:65:@8656.4]
  assign _T_8608 = _T_8603[4]; // @[Bitwise.scala 50:65:@8657.4]
  assign _T_8609 = _T_8603[5]; // @[Bitwise.scala 50:65:@8658.4]
  assign _T_8610 = _T_8603[6]; // @[Bitwise.scala 50:65:@8659.4]
  assign _T_8611 = _T_8603[7]; // @[Bitwise.scala 50:65:@8660.4]
  assign _T_8612 = _T_8603[8]; // @[Bitwise.scala 50:65:@8661.4]
  assign _T_8613 = _T_8603[9]; // @[Bitwise.scala 50:65:@8662.4]
  assign _T_8614 = _T_8603[10]; // @[Bitwise.scala 50:65:@8663.4]
  assign _T_8615 = _T_8603[11]; // @[Bitwise.scala 50:65:@8664.4]
  assign _T_8616 = _T_8603[12]; // @[Bitwise.scala 50:65:@8665.4]
  assign _T_8617 = _T_8603[13]; // @[Bitwise.scala 50:65:@8666.4]
  assign _T_8618 = _T_8603[14]; // @[Bitwise.scala 50:65:@8667.4]
  assign _T_8619 = _T_8603[15]; // @[Bitwise.scala 50:65:@8668.4]
  assign _T_8620 = _T_8603[16]; // @[Bitwise.scala 50:65:@8669.4]
  assign _T_8621 = _T_8603[17]; // @[Bitwise.scala 50:65:@8670.4]
  assign _T_8622 = _T_8603[18]; // @[Bitwise.scala 50:65:@8671.4]
  assign _T_8623 = _T_8603[19]; // @[Bitwise.scala 50:65:@8672.4]
  assign _T_8624 = _T_8603[20]; // @[Bitwise.scala 50:65:@8673.4]
  assign _T_8625 = _T_8603[21]; // @[Bitwise.scala 50:65:@8674.4]
  assign _T_8626 = _T_8603[22]; // @[Bitwise.scala 50:65:@8675.4]
  assign _T_8627 = _T_8603[23]; // @[Bitwise.scala 50:65:@8676.4]
  assign _T_8628 = _T_8603[24]; // @[Bitwise.scala 50:65:@8677.4]
  assign _T_8629 = _T_8603[25]; // @[Bitwise.scala 50:65:@8678.4]
  assign _T_8630 = _T_8603[26]; // @[Bitwise.scala 50:65:@8679.4]
  assign _T_8631 = _T_8603[27]; // @[Bitwise.scala 50:65:@8680.4]
  assign _T_8632 = _T_8603[28]; // @[Bitwise.scala 50:65:@8681.4]
  assign _T_8633 = _T_8603[29]; // @[Bitwise.scala 50:65:@8682.4]
  assign _T_8634 = _T_8603[30]; // @[Bitwise.scala 50:65:@8683.4]
  assign _T_8635 = _T_8603[31]; // @[Bitwise.scala 50:65:@8684.4]
  assign _T_8636 = _T_8603[32]; // @[Bitwise.scala 50:65:@8685.4]
  assign _T_8637 = _T_8603[33]; // @[Bitwise.scala 50:65:@8686.4]
  assign _T_8638 = _T_8603[34]; // @[Bitwise.scala 50:65:@8687.4]
  assign _T_8639 = _T_8603[35]; // @[Bitwise.scala 50:65:@8688.4]
  assign _T_8640 = _T_8603[36]; // @[Bitwise.scala 50:65:@8689.4]
  assign _T_8641 = _T_8603[37]; // @[Bitwise.scala 50:65:@8690.4]
  assign _T_8642 = _T_8603[38]; // @[Bitwise.scala 50:65:@8691.4]
  assign _T_8643 = _T_8603[39]; // @[Bitwise.scala 50:65:@8692.4]
  assign _T_8644 = _T_8603[40]; // @[Bitwise.scala 50:65:@8693.4]
  assign _T_8645 = _T_8603[41]; // @[Bitwise.scala 50:65:@8694.4]
  assign _T_8646 = _T_8603[42]; // @[Bitwise.scala 50:65:@8695.4]
  assign _T_8647 = _T_8603[43]; // @[Bitwise.scala 50:65:@8696.4]
  assign _T_8648 = _T_8603[44]; // @[Bitwise.scala 50:65:@8697.4]
  assign _T_8649 = _T_8603[45]; // @[Bitwise.scala 50:65:@8698.4]
  assign _T_8650 = _T_8603[46]; // @[Bitwise.scala 50:65:@8699.4]
  assign _T_8651 = _T_8603[47]; // @[Bitwise.scala 50:65:@8700.4]
  assign _T_8652 = _T_8603[48]; // @[Bitwise.scala 50:65:@8701.4]
  assign _T_8653 = _T_8603[49]; // @[Bitwise.scala 50:65:@8702.4]
  assign _T_8654 = _T_8603[50]; // @[Bitwise.scala 50:65:@8703.4]
  assign _T_8655 = _T_8603[51]; // @[Bitwise.scala 50:65:@8704.4]
  assign _T_8656 = _T_8603[52]; // @[Bitwise.scala 50:65:@8705.4]
  assign _T_8657 = _T_8603[53]; // @[Bitwise.scala 50:65:@8706.4]
  assign _T_8658 = _T_8603[54]; // @[Bitwise.scala 50:65:@8707.4]
  assign _T_8659 = _T_8605 + _T_8606; // @[Bitwise.scala 48:55:@8708.4]
  assign _GEN_952 = {{1'd0}, _T_8604}; // @[Bitwise.scala 48:55:@8709.4]
  assign _T_8660 = _GEN_952 + _T_8659; // @[Bitwise.scala 48:55:@8709.4]
  assign _T_8661 = _T_8608 + _T_8609; // @[Bitwise.scala 48:55:@8710.4]
  assign _GEN_953 = {{1'd0}, _T_8607}; // @[Bitwise.scala 48:55:@8711.4]
  assign _T_8662 = _GEN_953 + _T_8661; // @[Bitwise.scala 48:55:@8711.4]
  assign _T_8663 = _T_8660 + _T_8662; // @[Bitwise.scala 48:55:@8712.4]
  assign _T_8664 = _T_8611 + _T_8612; // @[Bitwise.scala 48:55:@8713.4]
  assign _GEN_954 = {{1'd0}, _T_8610}; // @[Bitwise.scala 48:55:@8714.4]
  assign _T_8665 = _GEN_954 + _T_8664; // @[Bitwise.scala 48:55:@8714.4]
  assign _T_8666 = _T_8613 + _T_8614; // @[Bitwise.scala 48:55:@8715.4]
  assign _T_8667 = _T_8615 + _T_8616; // @[Bitwise.scala 48:55:@8716.4]
  assign _T_8668 = _T_8666 + _T_8667; // @[Bitwise.scala 48:55:@8717.4]
  assign _T_8669 = _T_8665 + _T_8668; // @[Bitwise.scala 48:55:@8718.4]
  assign _T_8670 = _T_8663 + _T_8669; // @[Bitwise.scala 48:55:@8719.4]
  assign _T_8671 = _T_8618 + _T_8619; // @[Bitwise.scala 48:55:@8720.4]
  assign _GEN_955 = {{1'd0}, _T_8617}; // @[Bitwise.scala 48:55:@8721.4]
  assign _T_8672 = _GEN_955 + _T_8671; // @[Bitwise.scala 48:55:@8721.4]
  assign _T_8673 = _T_8620 + _T_8621; // @[Bitwise.scala 48:55:@8722.4]
  assign _T_8674 = _T_8622 + _T_8623; // @[Bitwise.scala 48:55:@8723.4]
  assign _T_8675 = _T_8673 + _T_8674; // @[Bitwise.scala 48:55:@8724.4]
  assign _T_8676 = _T_8672 + _T_8675; // @[Bitwise.scala 48:55:@8725.4]
  assign _T_8677 = _T_8625 + _T_8626; // @[Bitwise.scala 48:55:@8726.4]
  assign _GEN_956 = {{1'd0}, _T_8624}; // @[Bitwise.scala 48:55:@8727.4]
  assign _T_8678 = _GEN_956 + _T_8677; // @[Bitwise.scala 48:55:@8727.4]
  assign _T_8679 = _T_8627 + _T_8628; // @[Bitwise.scala 48:55:@8728.4]
  assign _T_8680 = _T_8629 + _T_8630; // @[Bitwise.scala 48:55:@8729.4]
  assign _T_8681 = _T_8679 + _T_8680; // @[Bitwise.scala 48:55:@8730.4]
  assign _T_8682 = _T_8678 + _T_8681; // @[Bitwise.scala 48:55:@8731.4]
  assign _T_8683 = _T_8676 + _T_8682; // @[Bitwise.scala 48:55:@8732.4]
  assign _T_8684 = _T_8670 + _T_8683; // @[Bitwise.scala 48:55:@8733.4]
  assign _T_8685 = _T_8632 + _T_8633; // @[Bitwise.scala 48:55:@8734.4]
  assign _GEN_957 = {{1'd0}, _T_8631}; // @[Bitwise.scala 48:55:@8735.4]
  assign _T_8686 = _GEN_957 + _T_8685; // @[Bitwise.scala 48:55:@8735.4]
  assign _T_8687 = _T_8634 + _T_8635; // @[Bitwise.scala 48:55:@8736.4]
  assign _T_8688 = _T_8636 + _T_8637; // @[Bitwise.scala 48:55:@8737.4]
  assign _T_8689 = _T_8687 + _T_8688; // @[Bitwise.scala 48:55:@8738.4]
  assign _T_8690 = _T_8686 + _T_8689; // @[Bitwise.scala 48:55:@8739.4]
  assign _T_8691 = _T_8639 + _T_8640; // @[Bitwise.scala 48:55:@8740.4]
  assign _GEN_958 = {{1'd0}, _T_8638}; // @[Bitwise.scala 48:55:@8741.4]
  assign _T_8692 = _GEN_958 + _T_8691; // @[Bitwise.scala 48:55:@8741.4]
  assign _T_8693 = _T_8641 + _T_8642; // @[Bitwise.scala 48:55:@8742.4]
  assign _T_8694 = _T_8643 + _T_8644; // @[Bitwise.scala 48:55:@8743.4]
  assign _T_8695 = _T_8693 + _T_8694; // @[Bitwise.scala 48:55:@8744.4]
  assign _T_8696 = _T_8692 + _T_8695; // @[Bitwise.scala 48:55:@8745.4]
  assign _T_8697 = _T_8690 + _T_8696; // @[Bitwise.scala 48:55:@8746.4]
  assign _T_8698 = _T_8646 + _T_8647; // @[Bitwise.scala 48:55:@8747.4]
  assign _GEN_959 = {{1'd0}, _T_8645}; // @[Bitwise.scala 48:55:@8748.4]
  assign _T_8699 = _GEN_959 + _T_8698; // @[Bitwise.scala 48:55:@8748.4]
  assign _T_8700 = _T_8648 + _T_8649; // @[Bitwise.scala 48:55:@8749.4]
  assign _T_8701 = _T_8650 + _T_8651; // @[Bitwise.scala 48:55:@8750.4]
  assign _T_8702 = _T_8700 + _T_8701; // @[Bitwise.scala 48:55:@8751.4]
  assign _T_8703 = _T_8699 + _T_8702; // @[Bitwise.scala 48:55:@8752.4]
  assign _T_8704 = _T_8653 + _T_8654; // @[Bitwise.scala 48:55:@8753.4]
  assign _GEN_960 = {{1'd0}, _T_8652}; // @[Bitwise.scala 48:55:@8754.4]
  assign _T_8705 = _GEN_960 + _T_8704; // @[Bitwise.scala 48:55:@8754.4]
  assign _T_8706 = _T_8655 + _T_8656; // @[Bitwise.scala 48:55:@8755.4]
  assign _T_8707 = _T_8657 + _T_8658; // @[Bitwise.scala 48:55:@8756.4]
  assign _T_8708 = _T_8706 + _T_8707; // @[Bitwise.scala 48:55:@8757.4]
  assign _T_8709 = _T_8705 + _T_8708; // @[Bitwise.scala 48:55:@8758.4]
  assign _T_8710 = _T_8703 + _T_8709; // @[Bitwise.scala 48:55:@8759.4]
  assign _T_8711 = _T_8697 + _T_8710; // @[Bitwise.scala 48:55:@8760.4]
  assign _T_8712 = _T_8684 + _T_8711; // @[Bitwise.scala 48:55:@8761.4]
  assign _T_8776 = _T_2230[55:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@8826.4]
  assign _T_8777 = _T_8776[0]; // @[Bitwise.scala 50:65:@8827.4]
  assign _T_8778 = _T_8776[1]; // @[Bitwise.scala 50:65:@8828.4]
  assign _T_8779 = _T_8776[2]; // @[Bitwise.scala 50:65:@8829.4]
  assign _T_8780 = _T_8776[3]; // @[Bitwise.scala 50:65:@8830.4]
  assign _T_8781 = _T_8776[4]; // @[Bitwise.scala 50:65:@8831.4]
  assign _T_8782 = _T_8776[5]; // @[Bitwise.scala 50:65:@8832.4]
  assign _T_8783 = _T_8776[6]; // @[Bitwise.scala 50:65:@8833.4]
  assign _T_8784 = _T_8776[7]; // @[Bitwise.scala 50:65:@8834.4]
  assign _T_8785 = _T_8776[8]; // @[Bitwise.scala 50:65:@8835.4]
  assign _T_8786 = _T_8776[9]; // @[Bitwise.scala 50:65:@8836.4]
  assign _T_8787 = _T_8776[10]; // @[Bitwise.scala 50:65:@8837.4]
  assign _T_8788 = _T_8776[11]; // @[Bitwise.scala 50:65:@8838.4]
  assign _T_8789 = _T_8776[12]; // @[Bitwise.scala 50:65:@8839.4]
  assign _T_8790 = _T_8776[13]; // @[Bitwise.scala 50:65:@8840.4]
  assign _T_8791 = _T_8776[14]; // @[Bitwise.scala 50:65:@8841.4]
  assign _T_8792 = _T_8776[15]; // @[Bitwise.scala 50:65:@8842.4]
  assign _T_8793 = _T_8776[16]; // @[Bitwise.scala 50:65:@8843.4]
  assign _T_8794 = _T_8776[17]; // @[Bitwise.scala 50:65:@8844.4]
  assign _T_8795 = _T_8776[18]; // @[Bitwise.scala 50:65:@8845.4]
  assign _T_8796 = _T_8776[19]; // @[Bitwise.scala 50:65:@8846.4]
  assign _T_8797 = _T_8776[20]; // @[Bitwise.scala 50:65:@8847.4]
  assign _T_8798 = _T_8776[21]; // @[Bitwise.scala 50:65:@8848.4]
  assign _T_8799 = _T_8776[22]; // @[Bitwise.scala 50:65:@8849.4]
  assign _T_8800 = _T_8776[23]; // @[Bitwise.scala 50:65:@8850.4]
  assign _T_8801 = _T_8776[24]; // @[Bitwise.scala 50:65:@8851.4]
  assign _T_8802 = _T_8776[25]; // @[Bitwise.scala 50:65:@8852.4]
  assign _T_8803 = _T_8776[26]; // @[Bitwise.scala 50:65:@8853.4]
  assign _T_8804 = _T_8776[27]; // @[Bitwise.scala 50:65:@8854.4]
  assign _T_8805 = _T_8776[28]; // @[Bitwise.scala 50:65:@8855.4]
  assign _T_8806 = _T_8776[29]; // @[Bitwise.scala 50:65:@8856.4]
  assign _T_8807 = _T_8776[30]; // @[Bitwise.scala 50:65:@8857.4]
  assign _T_8808 = _T_8776[31]; // @[Bitwise.scala 50:65:@8858.4]
  assign _T_8809 = _T_8776[32]; // @[Bitwise.scala 50:65:@8859.4]
  assign _T_8810 = _T_8776[33]; // @[Bitwise.scala 50:65:@8860.4]
  assign _T_8811 = _T_8776[34]; // @[Bitwise.scala 50:65:@8861.4]
  assign _T_8812 = _T_8776[35]; // @[Bitwise.scala 50:65:@8862.4]
  assign _T_8813 = _T_8776[36]; // @[Bitwise.scala 50:65:@8863.4]
  assign _T_8814 = _T_8776[37]; // @[Bitwise.scala 50:65:@8864.4]
  assign _T_8815 = _T_8776[38]; // @[Bitwise.scala 50:65:@8865.4]
  assign _T_8816 = _T_8776[39]; // @[Bitwise.scala 50:65:@8866.4]
  assign _T_8817 = _T_8776[40]; // @[Bitwise.scala 50:65:@8867.4]
  assign _T_8818 = _T_8776[41]; // @[Bitwise.scala 50:65:@8868.4]
  assign _T_8819 = _T_8776[42]; // @[Bitwise.scala 50:65:@8869.4]
  assign _T_8820 = _T_8776[43]; // @[Bitwise.scala 50:65:@8870.4]
  assign _T_8821 = _T_8776[44]; // @[Bitwise.scala 50:65:@8871.4]
  assign _T_8822 = _T_8776[45]; // @[Bitwise.scala 50:65:@8872.4]
  assign _T_8823 = _T_8776[46]; // @[Bitwise.scala 50:65:@8873.4]
  assign _T_8824 = _T_8776[47]; // @[Bitwise.scala 50:65:@8874.4]
  assign _T_8825 = _T_8776[48]; // @[Bitwise.scala 50:65:@8875.4]
  assign _T_8826 = _T_8776[49]; // @[Bitwise.scala 50:65:@8876.4]
  assign _T_8827 = _T_8776[50]; // @[Bitwise.scala 50:65:@8877.4]
  assign _T_8828 = _T_8776[51]; // @[Bitwise.scala 50:65:@8878.4]
  assign _T_8829 = _T_8776[52]; // @[Bitwise.scala 50:65:@8879.4]
  assign _T_8830 = _T_8776[53]; // @[Bitwise.scala 50:65:@8880.4]
  assign _T_8831 = _T_8776[54]; // @[Bitwise.scala 50:65:@8881.4]
  assign _T_8832 = _T_8776[55]; // @[Bitwise.scala 50:65:@8882.4]
  assign _T_8833 = _T_8778 + _T_8779; // @[Bitwise.scala 48:55:@8883.4]
  assign _GEN_961 = {{1'd0}, _T_8777}; // @[Bitwise.scala 48:55:@8884.4]
  assign _T_8834 = _GEN_961 + _T_8833; // @[Bitwise.scala 48:55:@8884.4]
  assign _T_8835 = _T_8780 + _T_8781; // @[Bitwise.scala 48:55:@8885.4]
  assign _T_8836 = _T_8782 + _T_8783; // @[Bitwise.scala 48:55:@8886.4]
  assign _T_8837 = _T_8835 + _T_8836; // @[Bitwise.scala 48:55:@8887.4]
  assign _T_8838 = _T_8834 + _T_8837; // @[Bitwise.scala 48:55:@8888.4]
  assign _T_8839 = _T_8785 + _T_8786; // @[Bitwise.scala 48:55:@8889.4]
  assign _GEN_962 = {{1'd0}, _T_8784}; // @[Bitwise.scala 48:55:@8890.4]
  assign _T_8840 = _GEN_962 + _T_8839; // @[Bitwise.scala 48:55:@8890.4]
  assign _T_8841 = _T_8787 + _T_8788; // @[Bitwise.scala 48:55:@8891.4]
  assign _T_8842 = _T_8789 + _T_8790; // @[Bitwise.scala 48:55:@8892.4]
  assign _T_8843 = _T_8841 + _T_8842; // @[Bitwise.scala 48:55:@8893.4]
  assign _T_8844 = _T_8840 + _T_8843; // @[Bitwise.scala 48:55:@8894.4]
  assign _T_8845 = _T_8838 + _T_8844; // @[Bitwise.scala 48:55:@8895.4]
  assign _T_8846 = _T_8792 + _T_8793; // @[Bitwise.scala 48:55:@8896.4]
  assign _GEN_963 = {{1'd0}, _T_8791}; // @[Bitwise.scala 48:55:@8897.4]
  assign _T_8847 = _GEN_963 + _T_8846; // @[Bitwise.scala 48:55:@8897.4]
  assign _T_8848 = _T_8794 + _T_8795; // @[Bitwise.scala 48:55:@8898.4]
  assign _T_8849 = _T_8796 + _T_8797; // @[Bitwise.scala 48:55:@8899.4]
  assign _T_8850 = _T_8848 + _T_8849; // @[Bitwise.scala 48:55:@8900.4]
  assign _T_8851 = _T_8847 + _T_8850; // @[Bitwise.scala 48:55:@8901.4]
  assign _T_8852 = _T_8799 + _T_8800; // @[Bitwise.scala 48:55:@8902.4]
  assign _GEN_964 = {{1'd0}, _T_8798}; // @[Bitwise.scala 48:55:@8903.4]
  assign _T_8853 = _GEN_964 + _T_8852; // @[Bitwise.scala 48:55:@8903.4]
  assign _T_8854 = _T_8801 + _T_8802; // @[Bitwise.scala 48:55:@8904.4]
  assign _T_8855 = _T_8803 + _T_8804; // @[Bitwise.scala 48:55:@8905.4]
  assign _T_8856 = _T_8854 + _T_8855; // @[Bitwise.scala 48:55:@8906.4]
  assign _T_8857 = _T_8853 + _T_8856; // @[Bitwise.scala 48:55:@8907.4]
  assign _T_8858 = _T_8851 + _T_8857; // @[Bitwise.scala 48:55:@8908.4]
  assign _T_8859 = _T_8845 + _T_8858; // @[Bitwise.scala 48:55:@8909.4]
  assign _T_8860 = _T_8806 + _T_8807; // @[Bitwise.scala 48:55:@8910.4]
  assign _GEN_965 = {{1'd0}, _T_8805}; // @[Bitwise.scala 48:55:@8911.4]
  assign _T_8861 = _GEN_965 + _T_8860; // @[Bitwise.scala 48:55:@8911.4]
  assign _T_8862 = _T_8808 + _T_8809; // @[Bitwise.scala 48:55:@8912.4]
  assign _T_8863 = _T_8810 + _T_8811; // @[Bitwise.scala 48:55:@8913.4]
  assign _T_8864 = _T_8862 + _T_8863; // @[Bitwise.scala 48:55:@8914.4]
  assign _T_8865 = _T_8861 + _T_8864; // @[Bitwise.scala 48:55:@8915.4]
  assign _T_8866 = _T_8813 + _T_8814; // @[Bitwise.scala 48:55:@8916.4]
  assign _GEN_966 = {{1'd0}, _T_8812}; // @[Bitwise.scala 48:55:@8917.4]
  assign _T_8867 = _GEN_966 + _T_8866; // @[Bitwise.scala 48:55:@8917.4]
  assign _T_8868 = _T_8815 + _T_8816; // @[Bitwise.scala 48:55:@8918.4]
  assign _T_8869 = _T_8817 + _T_8818; // @[Bitwise.scala 48:55:@8919.4]
  assign _T_8870 = _T_8868 + _T_8869; // @[Bitwise.scala 48:55:@8920.4]
  assign _T_8871 = _T_8867 + _T_8870; // @[Bitwise.scala 48:55:@8921.4]
  assign _T_8872 = _T_8865 + _T_8871; // @[Bitwise.scala 48:55:@8922.4]
  assign _T_8873 = _T_8820 + _T_8821; // @[Bitwise.scala 48:55:@8923.4]
  assign _GEN_967 = {{1'd0}, _T_8819}; // @[Bitwise.scala 48:55:@8924.4]
  assign _T_8874 = _GEN_967 + _T_8873; // @[Bitwise.scala 48:55:@8924.4]
  assign _T_8875 = _T_8822 + _T_8823; // @[Bitwise.scala 48:55:@8925.4]
  assign _T_8876 = _T_8824 + _T_8825; // @[Bitwise.scala 48:55:@8926.4]
  assign _T_8877 = _T_8875 + _T_8876; // @[Bitwise.scala 48:55:@8927.4]
  assign _T_8878 = _T_8874 + _T_8877; // @[Bitwise.scala 48:55:@8928.4]
  assign _T_8879 = _T_8827 + _T_8828; // @[Bitwise.scala 48:55:@8929.4]
  assign _GEN_968 = {{1'd0}, _T_8826}; // @[Bitwise.scala 48:55:@8930.4]
  assign _T_8880 = _GEN_968 + _T_8879; // @[Bitwise.scala 48:55:@8930.4]
  assign _T_8881 = _T_8829 + _T_8830; // @[Bitwise.scala 48:55:@8931.4]
  assign _T_8882 = _T_8831 + _T_8832; // @[Bitwise.scala 48:55:@8932.4]
  assign _T_8883 = _T_8881 + _T_8882; // @[Bitwise.scala 48:55:@8933.4]
  assign _T_8884 = _T_8880 + _T_8883; // @[Bitwise.scala 48:55:@8934.4]
  assign _T_8885 = _T_8878 + _T_8884; // @[Bitwise.scala 48:55:@8935.4]
  assign _T_8886 = _T_8872 + _T_8885; // @[Bitwise.scala 48:55:@8936.4]
  assign _T_8887 = _T_8859 + _T_8886; // @[Bitwise.scala 48:55:@8937.4]
  assign _T_8951 = _T_2230[56:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@9002.4]
  assign _T_8952 = _T_8951[0]; // @[Bitwise.scala 50:65:@9003.4]
  assign _T_8953 = _T_8951[1]; // @[Bitwise.scala 50:65:@9004.4]
  assign _T_8954 = _T_8951[2]; // @[Bitwise.scala 50:65:@9005.4]
  assign _T_8955 = _T_8951[3]; // @[Bitwise.scala 50:65:@9006.4]
  assign _T_8956 = _T_8951[4]; // @[Bitwise.scala 50:65:@9007.4]
  assign _T_8957 = _T_8951[5]; // @[Bitwise.scala 50:65:@9008.4]
  assign _T_8958 = _T_8951[6]; // @[Bitwise.scala 50:65:@9009.4]
  assign _T_8959 = _T_8951[7]; // @[Bitwise.scala 50:65:@9010.4]
  assign _T_8960 = _T_8951[8]; // @[Bitwise.scala 50:65:@9011.4]
  assign _T_8961 = _T_8951[9]; // @[Bitwise.scala 50:65:@9012.4]
  assign _T_8962 = _T_8951[10]; // @[Bitwise.scala 50:65:@9013.4]
  assign _T_8963 = _T_8951[11]; // @[Bitwise.scala 50:65:@9014.4]
  assign _T_8964 = _T_8951[12]; // @[Bitwise.scala 50:65:@9015.4]
  assign _T_8965 = _T_8951[13]; // @[Bitwise.scala 50:65:@9016.4]
  assign _T_8966 = _T_8951[14]; // @[Bitwise.scala 50:65:@9017.4]
  assign _T_8967 = _T_8951[15]; // @[Bitwise.scala 50:65:@9018.4]
  assign _T_8968 = _T_8951[16]; // @[Bitwise.scala 50:65:@9019.4]
  assign _T_8969 = _T_8951[17]; // @[Bitwise.scala 50:65:@9020.4]
  assign _T_8970 = _T_8951[18]; // @[Bitwise.scala 50:65:@9021.4]
  assign _T_8971 = _T_8951[19]; // @[Bitwise.scala 50:65:@9022.4]
  assign _T_8972 = _T_8951[20]; // @[Bitwise.scala 50:65:@9023.4]
  assign _T_8973 = _T_8951[21]; // @[Bitwise.scala 50:65:@9024.4]
  assign _T_8974 = _T_8951[22]; // @[Bitwise.scala 50:65:@9025.4]
  assign _T_8975 = _T_8951[23]; // @[Bitwise.scala 50:65:@9026.4]
  assign _T_8976 = _T_8951[24]; // @[Bitwise.scala 50:65:@9027.4]
  assign _T_8977 = _T_8951[25]; // @[Bitwise.scala 50:65:@9028.4]
  assign _T_8978 = _T_8951[26]; // @[Bitwise.scala 50:65:@9029.4]
  assign _T_8979 = _T_8951[27]; // @[Bitwise.scala 50:65:@9030.4]
  assign _T_8980 = _T_8951[28]; // @[Bitwise.scala 50:65:@9031.4]
  assign _T_8981 = _T_8951[29]; // @[Bitwise.scala 50:65:@9032.4]
  assign _T_8982 = _T_8951[30]; // @[Bitwise.scala 50:65:@9033.4]
  assign _T_8983 = _T_8951[31]; // @[Bitwise.scala 50:65:@9034.4]
  assign _T_8984 = _T_8951[32]; // @[Bitwise.scala 50:65:@9035.4]
  assign _T_8985 = _T_8951[33]; // @[Bitwise.scala 50:65:@9036.4]
  assign _T_8986 = _T_8951[34]; // @[Bitwise.scala 50:65:@9037.4]
  assign _T_8987 = _T_8951[35]; // @[Bitwise.scala 50:65:@9038.4]
  assign _T_8988 = _T_8951[36]; // @[Bitwise.scala 50:65:@9039.4]
  assign _T_8989 = _T_8951[37]; // @[Bitwise.scala 50:65:@9040.4]
  assign _T_8990 = _T_8951[38]; // @[Bitwise.scala 50:65:@9041.4]
  assign _T_8991 = _T_8951[39]; // @[Bitwise.scala 50:65:@9042.4]
  assign _T_8992 = _T_8951[40]; // @[Bitwise.scala 50:65:@9043.4]
  assign _T_8993 = _T_8951[41]; // @[Bitwise.scala 50:65:@9044.4]
  assign _T_8994 = _T_8951[42]; // @[Bitwise.scala 50:65:@9045.4]
  assign _T_8995 = _T_8951[43]; // @[Bitwise.scala 50:65:@9046.4]
  assign _T_8996 = _T_8951[44]; // @[Bitwise.scala 50:65:@9047.4]
  assign _T_8997 = _T_8951[45]; // @[Bitwise.scala 50:65:@9048.4]
  assign _T_8998 = _T_8951[46]; // @[Bitwise.scala 50:65:@9049.4]
  assign _T_8999 = _T_8951[47]; // @[Bitwise.scala 50:65:@9050.4]
  assign _T_9000 = _T_8951[48]; // @[Bitwise.scala 50:65:@9051.4]
  assign _T_9001 = _T_8951[49]; // @[Bitwise.scala 50:65:@9052.4]
  assign _T_9002 = _T_8951[50]; // @[Bitwise.scala 50:65:@9053.4]
  assign _T_9003 = _T_8951[51]; // @[Bitwise.scala 50:65:@9054.4]
  assign _T_9004 = _T_8951[52]; // @[Bitwise.scala 50:65:@9055.4]
  assign _T_9005 = _T_8951[53]; // @[Bitwise.scala 50:65:@9056.4]
  assign _T_9006 = _T_8951[54]; // @[Bitwise.scala 50:65:@9057.4]
  assign _T_9007 = _T_8951[55]; // @[Bitwise.scala 50:65:@9058.4]
  assign _T_9008 = _T_8951[56]; // @[Bitwise.scala 50:65:@9059.4]
  assign _T_9009 = _T_8953 + _T_8954; // @[Bitwise.scala 48:55:@9060.4]
  assign _GEN_969 = {{1'd0}, _T_8952}; // @[Bitwise.scala 48:55:@9061.4]
  assign _T_9010 = _GEN_969 + _T_9009; // @[Bitwise.scala 48:55:@9061.4]
  assign _T_9011 = _T_8955 + _T_8956; // @[Bitwise.scala 48:55:@9062.4]
  assign _T_9012 = _T_8957 + _T_8958; // @[Bitwise.scala 48:55:@9063.4]
  assign _T_9013 = _T_9011 + _T_9012; // @[Bitwise.scala 48:55:@9064.4]
  assign _T_9014 = _T_9010 + _T_9013; // @[Bitwise.scala 48:55:@9065.4]
  assign _T_9015 = _T_8960 + _T_8961; // @[Bitwise.scala 48:55:@9066.4]
  assign _GEN_970 = {{1'd0}, _T_8959}; // @[Bitwise.scala 48:55:@9067.4]
  assign _T_9016 = _GEN_970 + _T_9015; // @[Bitwise.scala 48:55:@9067.4]
  assign _T_9017 = _T_8962 + _T_8963; // @[Bitwise.scala 48:55:@9068.4]
  assign _T_9018 = _T_8964 + _T_8965; // @[Bitwise.scala 48:55:@9069.4]
  assign _T_9019 = _T_9017 + _T_9018; // @[Bitwise.scala 48:55:@9070.4]
  assign _T_9020 = _T_9016 + _T_9019; // @[Bitwise.scala 48:55:@9071.4]
  assign _T_9021 = _T_9014 + _T_9020; // @[Bitwise.scala 48:55:@9072.4]
  assign _T_9022 = _T_8967 + _T_8968; // @[Bitwise.scala 48:55:@9073.4]
  assign _GEN_971 = {{1'd0}, _T_8966}; // @[Bitwise.scala 48:55:@9074.4]
  assign _T_9023 = _GEN_971 + _T_9022; // @[Bitwise.scala 48:55:@9074.4]
  assign _T_9024 = _T_8969 + _T_8970; // @[Bitwise.scala 48:55:@9075.4]
  assign _T_9025 = _T_8971 + _T_8972; // @[Bitwise.scala 48:55:@9076.4]
  assign _T_9026 = _T_9024 + _T_9025; // @[Bitwise.scala 48:55:@9077.4]
  assign _T_9027 = _T_9023 + _T_9026; // @[Bitwise.scala 48:55:@9078.4]
  assign _T_9028 = _T_8974 + _T_8975; // @[Bitwise.scala 48:55:@9079.4]
  assign _GEN_972 = {{1'd0}, _T_8973}; // @[Bitwise.scala 48:55:@9080.4]
  assign _T_9029 = _GEN_972 + _T_9028; // @[Bitwise.scala 48:55:@9080.4]
  assign _T_9030 = _T_8976 + _T_8977; // @[Bitwise.scala 48:55:@9081.4]
  assign _T_9031 = _T_8978 + _T_8979; // @[Bitwise.scala 48:55:@9082.4]
  assign _T_9032 = _T_9030 + _T_9031; // @[Bitwise.scala 48:55:@9083.4]
  assign _T_9033 = _T_9029 + _T_9032; // @[Bitwise.scala 48:55:@9084.4]
  assign _T_9034 = _T_9027 + _T_9033; // @[Bitwise.scala 48:55:@9085.4]
  assign _T_9035 = _T_9021 + _T_9034; // @[Bitwise.scala 48:55:@9086.4]
  assign _T_9036 = _T_8981 + _T_8982; // @[Bitwise.scala 48:55:@9087.4]
  assign _GEN_973 = {{1'd0}, _T_8980}; // @[Bitwise.scala 48:55:@9088.4]
  assign _T_9037 = _GEN_973 + _T_9036; // @[Bitwise.scala 48:55:@9088.4]
  assign _T_9038 = _T_8983 + _T_8984; // @[Bitwise.scala 48:55:@9089.4]
  assign _T_9039 = _T_8985 + _T_8986; // @[Bitwise.scala 48:55:@9090.4]
  assign _T_9040 = _T_9038 + _T_9039; // @[Bitwise.scala 48:55:@9091.4]
  assign _T_9041 = _T_9037 + _T_9040; // @[Bitwise.scala 48:55:@9092.4]
  assign _T_9042 = _T_8988 + _T_8989; // @[Bitwise.scala 48:55:@9093.4]
  assign _GEN_974 = {{1'd0}, _T_8987}; // @[Bitwise.scala 48:55:@9094.4]
  assign _T_9043 = _GEN_974 + _T_9042; // @[Bitwise.scala 48:55:@9094.4]
  assign _T_9044 = _T_8990 + _T_8991; // @[Bitwise.scala 48:55:@9095.4]
  assign _T_9045 = _T_8992 + _T_8993; // @[Bitwise.scala 48:55:@9096.4]
  assign _T_9046 = _T_9044 + _T_9045; // @[Bitwise.scala 48:55:@9097.4]
  assign _T_9047 = _T_9043 + _T_9046; // @[Bitwise.scala 48:55:@9098.4]
  assign _T_9048 = _T_9041 + _T_9047; // @[Bitwise.scala 48:55:@9099.4]
  assign _T_9049 = _T_8995 + _T_8996; // @[Bitwise.scala 48:55:@9100.4]
  assign _GEN_975 = {{1'd0}, _T_8994}; // @[Bitwise.scala 48:55:@9101.4]
  assign _T_9050 = _GEN_975 + _T_9049; // @[Bitwise.scala 48:55:@9101.4]
  assign _T_9051 = _T_8997 + _T_8998; // @[Bitwise.scala 48:55:@9102.4]
  assign _T_9052 = _T_8999 + _T_9000; // @[Bitwise.scala 48:55:@9103.4]
  assign _T_9053 = _T_9051 + _T_9052; // @[Bitwise.scala 48:55:@9104.4]
  assign _T_9054 = _T_9050 + _T_9053; // @[Bitwise.scala 48:55:@9105.4]
  assign _T_9055 = _T_9001 + _T_9002; // @[Bitwise.scala 48:55:@9106.4]
  assign _T_9056 = _T_9003 + _T_9004; // @[Bitwise.scala 48:55:@9107.4]
  assign _T_9057 = _T_9055 + _T_9056; // @[Bitwise.scala 48:55:@9108.4]
  assign _T_9058 = _T_9005 + _T_9006; // @[Bitwise.scala 48:55:@9109.4]
  assign _T_9059 = _T_9007 + _T_9008; // @[Bitwise.scala 48:55:@9110.4]
  assign _T_9060 = _T_9058 + _T_9059; // @[Bitwise.scala 48:55:@9111.4]
  assign _T_9061 = _T_9057 + _T_9060; // @[Bitwise.scala 48:55:@9112.4]
  assign _T_9062 = _T_9054 + _T_9061; // @[Bitwise.scala 48:55:@9113.4]
  assign _T_9063 = _T_9048 + _T_9062; // @[Bitwise.scala 48:55:@9114.4]
  assign _T_9064 = _T_9035 + _T_9063; // @[Bitwise.scala 48:55:@9115.4]
  assign _T_9128 = _T_2230[57:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@9180.4]
  assign _T_9129 = _T_9128[0]; // @[Bitwise.scala 50:65:@9181.4]
  assign _T_9130 = _T_9128[1]; // @[Bitwise.scala 50:65:@9182.4]
  assign _T_9131 = _T_9128[2]; // @[Bitwise.scala 50:65:@9183.4]
  assign _T_9132 = _T_9128[3]; // @[Bitwise.scala 50:65:@9184.4]
  assign _T_9133 = _T_9128[4]; // @[Bitwise.scala 50:65:@9185.4]
  assign _T_9134 = _T_9128[5]; // @[Bitwise.scala 50:65:@9186.4]
  assign _T_9135 = _T_9128[6]; // @[Bitwise.scala 50:65:@9187.4]
  assign _T_9136 = _T_9128[7]; // @[Bitwise.scala 50:65:@9188.4]
  assign _T_9137 = _T_9128[8]; // @[Bitwise.scala 50:65:@9189.4]
  assign _T_9138 = _T_9128[9]; // @[Bitwise.scala 50:65:@9190.4]
  assign _T_9139 = _T_9128[10]; // @[Bitwise.scala 50:65:@9191.4]
  assign _T_9140 = _T_9128[11]; // @[Bitwise.scala 50:65:@9192.4]
  assign _T_9141 = _T_9128[12]; // @[Bitwise.scala 50:65:@9193.4]
  assign _T_9142 = _T_9128[13]; // @[Bitwise.scala 50:65:@9194.4]
  assign _T_9143 = _T_9128[14]; // @[Bitwise.scala 50:65:@9195.4]
  assign _T_9144 = _T_9128[15]; // @[Bitwise.scala 50:65:@9196.4]
  assign _T_9145 = _T_9128[16]; // @[Bitwise.scala 50:65:@9197.4]
  assign _T_9146 = _T_9128[17]; // @[Bitwise.scala 50:65:@9198.4]
  assign _T_9147 = _T_9128[18]; // @[Bitwise.scala 50:65:@9199.4]
  assign _T_9148 = _T_9128[19]; // @[Bitwise.scala 50:65:@9200.4]
  assign _T_9149 = _T_9128[20]; // @[Bitwise.scala 50:65:@9201.4]
  assign _T_9150 = _T_9128[21]; // @[Bitwise.scala 50:65:@9202.4]
  assign _T_9151 = _T_9128[22]; // @[Bitwise.scala 50:65:@9203.4]
  assign _T_9152 = _T_9128[23]; // @[Bitwise.scala 50:65:@9204.4]
  assign _T_9153 = _T_9128[24]; // @[Bitwise.scala 50:65:@9205.4]
  assign _T_9154 = _T_9128[25]; // @[Bitwise.scala 50:65:@9206.4]
  assign _T_9155 = _T_9128[26]; // @[Bitwise.scala 50:65:@9207.4]
  assign _T_9156 = _T_9128[27]; // @[Bitwise.scala 50:65:@9208.4]
  assign _T_9157 = _T_9128[28]; // @[Bitwise.scala 50:65:@9209.4]
  assign _T_9158 = _T_9128[29]; // @[Bitwise.scala 50:65:@9210.4]
  assign _T_9159 = _T_9128[30]; // @[Bitwise.scala 50:65:@9211.4]
  assign _T_9160 = _T_9128[31]; // @[Bitwise.scala 50:65:@9212.4]
  assign _T_9161 = _T_9128[32]; // @[Bitwise.scala 50:65:@9213.4]
  assign _T_9162 = _T_9128[33]; // @[Bitwise.scala 50:65:@9214.4]
  assign _T_9163 = _T_9128[34]; // @[Bitwise.scala 50:65:@9215.4]
  assign _T_9164 = _T_9128[35]; // @[Bitwise.scala 50:65:@9216.4]
  assign _T_9165 = _T_9128[36]; // @[Bitwise.scala 50:65:@9217.4]
  assign _T_9166 = _T_9128[37]; // @[Bitwise.scala 50:65:@9218.4]
  assign _T_9167 = _T_9128[38]; // @[Bitwise.scala 50:65:@9219.4]
  assign _T_9168 = _T_9128[39]; // @[Bitwise.scala 50:65:@9220.4]
  assign _T_9169 = _T_9128[40]; // @[Bitwise.scala 50:65:@9221.4]
  assign _T_9170 = _T_9128[41]; // @[Bitwise.scala 50:65:@9222.4]
  assign _T_9171 = _T_9128[42]; // @[Bitwise.scala 50:65:@9223.4]
  assign _T_9172 = _T_9128[43]; // @[Bitwise.scala 50:65:@9224.4]
  assign _T_9173 = _T_9128[44]; // @[Bitwise.scala 50:65:@9225.4]
  assign _T_9174 = _T_9128[45]; // @[Bitwise.scala 50:65:@9226.4]
  assign _T_9175 = _T_9128[46]; // @[Bitwise.scala 50:65:@9227.4]
  assign _T_9176 = _T_9128[47]; // @[Bitwise.scala 50:65:@9228.4]
  assign _T_9177 = _T_9128[48]; // @[Bitwise.scala 50:65:@9229.4]
  assign _T_9178 = _T_9128[49]; // @[Bitwise.scala 50:65:@9230.4]
  assign _T_9179 = _T_9128[50]; // @[Bitwise.scala 50:65:@9231.4]
  assign _T_9180 = _T_9128[51]; // @[Bitwise.scala 50:65:@9232.4]
  assign _T_9181 = _T_9128[52]; // @[Bitwise.scala 50:65:@9233.4]
  assign _T_9182 = _T_9128[53]; // @[Bitwise.scala 50:65:@9234.4]
  assign _T_9183 = _T_9128[54]; // @[Bitwise.scala 50:65:@9235.4]
  assign _T_9184 = _T_9128[55]; // @[Bitwise.scala 50:65:@9236.4]
  assign _T_9185 = _T_9128[56]; // @[Bitwise.scala 50:65:@9237.4]
  assign _T_9186 = _T_9128[57]; // @[Bitwise.scala 50:65:@9238.4]
  assign _T_9187 = _T_9130 + _T_9131; // @[Bitwise.scala 48:55:@9239.4]
  assign _GEN_976 = {{1'd0}, _T_9129}; // @[Bitwise.scala 48:55:@9240.4]
  assign _T_9188 = _GEN_976 + _T_9187; // @[Bitwise.scala 48:55:@9240.4]
  assign _T_9189 = _T_9132 + _T_9133; // @[Bitwise.scala 48:55:@9241.4]
  assign _T_9190 = _T_9134 + _T_9135; // @[Bitwise.scala 48:55:@9242.4]
  assign _T_9191 = _T_9189 + _T_9190; // @[Bitwise.scala 48:55:@9243.4]
  assign _T_9192 = _T_9188 + _T_9191; // @[Bitwise.scala 48:55:@9244.4]
  assign _T_9193 = _T_9137 + _T_9138; // @[Bitwise.scala 48:55:@9245.4]
  assign _GEN_977 = {{1'd0}, _T_9136}; // @[Bitwise.scala 48:55:@9246.4]
  assign _T_9194 = _GEN_977 + _T_9193; // @[Bitwise.scala 48:55:@9246.4]
  assign _T_9195 = _T_9139 + _T_9140; // @[Bitwise.scala 48:55:@9247.4]
  assign _T_9196 = _T_9141 + _T_9142; // @[Bitwise.scala 48:55:@9248.4]
  assign _T_9197 = _T_9195 + _T_9196; // @[Bitwise.scala 48:55:@9249.4]
  assign _T_9198 = _T_9194 + _T_9197; // @[Bitwise.scala 48:55:@9250.4]
  assign _T_9199 = _T_9192 + _T_9198; // @[Bitwise.scala 48:55:@9251.4]
  assign _T_9200 = _T_9144 + _T_9145; // @[Bitwise.scala 48:55:@9252.4]
  assign _GEN_978 = {{1'd0}, _T_9143}; // @[Bitwise.scala 48:55:@9253.4]
  assign _T_9201 = _GEN_978 + _T_9200; // @[Bitwise.scala 48:55:@9253.4]
  assign _T_9202 = _T_9146 + _T_9147; // @[Bitwise.scala 48:55:@9254.4]
  assign _T_9203 = _T_9148 + _T_9149; // @[Bitwise.scala 48:55:@9255.4]
  assign _T_9204 = _T_9202 + _T_9203; // @[Bitwise.scala 48:55:@9256.4]
  assign _T_9205 = _T_9201 + _T_9204; // @[Bitwise.scala 48:55:@9257.4]
  assign _T_9206 = _T_9150 + _T_9151; // @[Bitwise.scala 48:55:@9258.4]
  assign _T_9207 = _T_9152 + _T_9153; // @[Bitwise.scala 48:55:@9259.4]
  assign _T_9208 = _T_9206 + _T_9207; // @[Bitwise.scala 48:55:@9260.4]
  assign _T_9209 = _T_9154 + _T_9155; // @[Bitwise.scala 48:55:@9261.4]
  assign _T_9210 = _T_9156 + _T_9157; // @[Bitwise.scala 48:55:@9262.4]
  assign _T_9211 = _T_9209 + _T_9210; // @[Bitwise.scala 48:55:@9263.4]
  assign _T_9212 = _T_9208 + _T_9211; // @[Bitwise.scala 48:55:@9264.4]
  assign _T_9213 = _T_9205 + _T_9212; // @[Bitwise.scala 48:55:@9265.4]
  assign _T_9214 = _T_9199 + _T_9213; // @[Bitwise.scala 48:55:@9266.4]
  assign _T_9215 = _T_9159 + _T_9160; // @[Bitwise.scala 48:55:@9267.4]
  assign _GEN_979 = {{1'd0}, _T_9158}; // @[Bitwise.scala 48:55:@9268.4]
  assign _T_9216 = _GEN_979 + _T_9215; // @[Bitwise.scala 48:55:@9268.4]
  assign _T_9217 = _T_9161 + _T_9162; // @[Bitwise.scala 48:55:@9269.4]
  assign _T_9218 = _T_9163 + _T_9164; // @[Bitwise.scala 48:55:@9270.4]
  assign _T_9219 = _T_9217 + _T_9218; // @[Bitwise.scala 48:55:@9271.4]
  assign _T_9220 = _T_9216 + _T_9219; // @[Bitwise.scala 48:55:@9272.4]
  assign _T_9221 = _T_9166 + _T_9167; // @[Bitwise.scala 48:55:@9273.4]
  assign _GEN_980 = {{1'd0}, _T_9165}; // @[Bitwise.scala 48:55:@9274.4]
  assign _T_9222 = _GEN_980 + _T_9221; // @[Bitwise.scala 48:55:@9274.4]
  assign _T_9223 = _T_9168 + _T_9169; // @[Bitwise.scala 48:55:@9275.4]
  assign _T_9224 = _T_9170 + _T_9171; // @[Bitwise.scala 48:55:@9276.4]
  assign _T_9225 = _T_9223 + _T_9224; // @[Bitwise.scala 48:55:@9277.4]
  assign _T_9226 = _T_9222 + _T_9225; // @[Bitwise.scala 48:55:@9278.4]
  assign _T_9227 = _T_9220 + _T_9226; // @[Bitwise.scala 48:55:@9279.4]
  assign _T_9228 = _T_9173 + _T_9174; // @[Bitwise.scala 48:55:@9280.4]
  assign _GEN_981 = {{1'd0}, _T_9172}; // @[Bitwise.scala 48:55:@9281.4]
  assign _T_9229 = _GEN_981 + _T_9228; // @[Bitwise.scala 48:55:@9281.4]
  assign _T_9230 = _T_9175 + _T_9176; // @[Bitwise.scala 48:55:@9282.4]
  assign _T_9231 = _T_9177 + _T_9178; // @[Bitwise.scala 48:55:@9283.4]
  assign _T_9232 = _T_9230 + _T_9231; // @[Bitwise.scala 48:55:@9284.4]
  assign _T_9233 = _T_9229 + _T_9232; // @[Bitwise.scala 48:55:@9285.4]
  assign _T_9234 = _T_9179 + _T_9180; // @[Bitwise.scala 48:55:@9286.4]
  assign _T_9235 = _T_9181 + _T_9182; // @[Bitwise.scala 48:55:@9287.4]
  assign _T_9236 = _T_9234 + _T_9235; // @[Bitwise.scala 48:55:@9288.4]
  assign _T_9237 = _T_9183 + _T_9184; // @[Bitwise.scala 48:55:@9289.4]
  assign _T_9238 = _T_9185 + _T_9186; // @[Bitwise.scala 48:55:@9290.4]
  assign _T_9239 = _T_9237 + _T_9238; // @[Bitwise.scala 48:55:@9291.4]
  assign _T_9240 = _T_9236 + _T_9239; // @[Bitwise.scala 48:55:@9292.4]
  assign _T_9241 = _T_9233 + _T_9240; // @[Bitwise.scala 48:55:@9293.4]
  assign _T_9242 = _T_9227 + _T_9241; // @[Bitwise.scala 48:55:@9294.4]
  assign _T_9243 = _T_9214 + _T_9242; // @[Bitwise.scala 48:55:@9295.4]
  assign _T_9307 = _T_2230[58:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@9360.4]
  assign _T_9308 = _T_9307[0]; // @[Bitwise.scala 50:65:@9361.4]
  assign _T_9309 = _T_9307[1]; // @[Bitwise.scala 50:65:@9362.4]
  assign _T_9310 = _T_9307[2]; // @[Bitwise.scala 50:65:@9363.4]
  assign _T_9311 = _T_9307[3]; // @[Bitwise.scala 50:65:@9364.4]
  assign _T_9312 = _T_9307[4]; // @[Bitwise.scala 50:65:@9365.4]
  assign _T_9313 = _T_9307[5]; // @[Bitwise.scala 50:65:@9366.4]
  assign _T_9314 = _T_9307[6]; // @[Bitwise.scala 50:65:@9367.4]
  assign _T_9315 = _T_9307[7]; // @[Bitwise.scala 50:65:@9368.4]
  assign _T_9316 = _T_9307[8]; // @[Bitwise.scala 50:65:@9369.4]
  assign _T_9317 = _T_9307[9]; // @[Bitwise.scala 50:65:@9370.4]
  assign _T_9318 = _T_9307[10]; // @[Bitwise.scala 50:65:@9371.4]
  assign _T_9319 = _T_9307[11]; // @[Bitwise.scala 50:65:@9372.4]
  assign _T_9320 = _T_9307[12]; // @[Bitwise.scala 50:65:@9373.4]
  assign _T_9321 = _T_9307[13]; // @[Bitwise.scala 50:65:@9374.4]
  assign _T_9322 = _T_9307[14]; // @[Bitwise.scala 50:65:@9375.4]
  assign _T_9323 = _T_9307[15]; // @[Bitwise.scala 50:65:@9376.4]
  assign _T_9324 = _T_9307[16]; // @[Bitwise.scala 50:65:@9377.4]
  assign _T_9325 = _T_9307[17]; // @[Bitwise.scala 50:65:@9378.4]
  assign _T_9326 = _T_9307[18]; // @[Bitwise.scala 50:65:@9379.4]
  assign _T_9327 = _T_9307[19]; // @[Bitwise.scala 50:65:@9380.4]
  assign _T_9328 = _T_9307[20]; // @[Bitwise.scala 50:65:@9381.4]
  assign _T_9329 = _T_9307[21]; // @[Bitwise.scala 50:65:@9382.4]
  assign _T_9330 = _T_9307[22]; // @[Bitwise.scala 50:65:@9383.4]
  assign _T_9331 = _T_9307[23]; // @[Bitwise.scala 50:65:@9384.4]
  assign _T_9332 = _T_9307[24]; // @[Bitwise.scala 50:65:@9385.4]
  assign _T_9333 = _T_9307[25]; // @[Bitwise.scala 50:65:@9386.4]
  assign _T_9334 = _T_9307[26]; // @[Bitwise.scala 50:65:@9387.4]
  assign _T_9335 = _T_9307[27]; // @[Bitwise.scala 50:65:@9388.4]
  assign _T_9336 = _T_9307[28]; // @[Bitwise.scala 50:65:@9389.4]
  assign _T_9337 = _T_9307[29]; // @[Bitwise.scala 50:65:@9390.4]
  assign _T_9338 = _T_9307[30]; // @[Bitwise.scala 50:65:@9391.4]
  assign _T_9339 = _T_9307[31]; // @[Bitwise.scala 50:65:@9392.4]
  assign _T_9340 = _T_9307[32]; // @[Bitwise.scala 50:65:@9393.4]
  assign _T_9341 = _T_9307[33]; // @[Bitwise.scala 50:65:@9394.4]
  assign _T_9342 = _T_9307[34]; // @[Bitwise.scala 50:65:@9395.4]
  assign _T_9343 = _T_9307[35]; // @[Bitwise.scala 50:65:@9396.4]
  assign _T_9344 = _T_9307[36]; // @[Bitwise.scala 50:65:@9397.4]
  assign _T_9345 = _T_9307[37]; // @[Bitwise.scala 50:65:@9398.4]
  assign _T_9346 = _T_9307[38]; // @[Bitwise.scala 50:65:@9399.4]
  assign _T_9347 = _T_9307[39]; // @[Bitwise.scala 50:65:@9400.4]
  assign _T_9348 = _T_9307[40]; // @[Bitwise.scala 50:65:@9401.4]
  assign _T_9349 = _T_9307[41]; // @[Bitwise.scala 50:65:@9402.4]
  assign _T_9350 = _T_9307[42]; // @[Bitwise.scala 50:65:@9403.4]
  assign _T_9351 = _T_9307[43]; // @[Bitwise.scala 50:65:@9404.4]
  assign _T_9352 = _T_9307[44]; // @[Bitwise.scala 50:65:@9405.4]
  assign _T_9353 = _T_9307[45]; // @[Bitwise.scala 50:65:@9406.4]
  assign _T_9354 = _T_9307[46]; // @[Bitwise.scala 50:65:@9407.4]
  assign _T_9355 = _T_9307[47]; // @[Bitwise.scala 50:65:@9408.4]
  assign _T_9356 = _T_9307[48]; // @[Bitwise.scala 50:65:@9409.4]
  assign _T_9357 = _T_9307[49]; // @[Bitwise.scala 50:65:@9410.4]
  assign _T_9358 = _T_9307[50]; // @[Bitwise.scala 50:65:@9411.4]
  assign _T_9359 = _T_9307[51]; // @[Bitwise.scala 50:65:@9412.4]
  assign _T_9360 = _T_9307[52]; // @[Bitwise.scala 50:65:@9413.4]
  assign _T_9361 = _T_9307[53]; // @[Bitwise.scala 50:65:@9414.4]
  assign _T_9362 = _T_9307[54]; // @[Bitwise.scala 50:65:@9415.4]
  assign _T_9363 = _T_9307[55]; // @[Bitwise.scala 50:65:@9416.4]
  assign _T_9364 = _T_9307[56]; // @[Bitwise.scala 50:65:@9417.4]
  assign _T_9365 = _T_9307[57]; // @[Bitwise.scala 50:65:@9418.4]
  assign _T_9366 = _T_9307[58]; // @[Bitwise.scala 50:65:@9419.4]
  assign _T_9367 = _T_9309 + _T_9310; // @[Bitwise.scala 48:55:@9420.4]
  assign _GEN_982 = {{1'd0}, _T_9308}; // @[Bitwise.scala 48:55:@9421.4]
  assign _T_9368 = _GEN_982 + _T_9367; // @[Bitwise.scala 48:55:@9421.4]
  assign _T_9369 = _T_9311 + _T_9312; // @[Bitwise.scala 48:55:@9422.4]
  assign _T_9370 = _T_9313 + _T_9314; // @[Bitwise.scala 48:55:@9423.4]
  assign _T_9371 = _T_9369 + _T_9370; // @[Bitwise.scala 48:55:@9424.4]
  assign _T_9372 = _T_9368 + _T_9371; // @[Bitwise.scala 48:55:@9425.4]
  assign _T_9373 = _T_9316 + _T_9317; // @[Bitwise.scala 48:55:@9426.4]
  assign _GEN_983 = {{1'd0}, _T_9315}; // @[Bitwise.scala 48:55:@9427.4]
  assign _T_9374 = _GEN_983 + _T_9373; // @[Bitwise.scala 48:55:@9427.4]
  assign _T_9375 = _T_9318 + _T_9319; // @[Bitwise.scala 48:55:@9428.4]
  assign _T_9376 = _T_9320 + _T_9321; // @[Bitwise.scala 48:55:@9429.4]
  assign _T_9377 = _T_9375 + _T_9376; // @[Bitwise.scala 48:55:@9430.4]
  assign _T_9378 = _T_9374 + _T_9377; // @[Bitwise.scala 48:55:@9431.4]
  assign _T_9379 = _T_9372 + _T_9378; // @[Bitwise.scala 48:55:@9432.4]
  assign _T_9380 = _T_9323 + _T_9324; // @[Bitwise.scala 48:55:@9433.4]
  assign _GEN_984 = {{1'd0}, _T_9322}; // @[Bitwise.scala 48:55:@9434.4]
  assign _T_9381 = _GEN_984 + _T_9380; // @[Bitwise.scala 48:55:@9434.4]
  assign _T_9382 = _T_9325 + _T_9326; // @[Bitwise.scala 48:55:@9435.4]
  assign _T_9383 = _T_9327 + _T_9328; // @[Bitwise.scala 48:55:@9436.4]
  assign _T_9384 = _T_9382 + _T_9383; // @[Bitwise.scala 48:55:@9437.4]
  assign _T_9385 = _T_9381 + _T_9384; // @[Bitwise.scala 48:55:@9438.4]
  assign _T_9386 = _T_9329 + _T_9330; // @[Bitwise.scala 48:55:@9439.4]
  assign _T_9387 = _T_9331 + _T_9332; // @[Bitwise.scala 48:55:@9440.4]
  assign _T_9388 = _T_9386 + _T_9387; // @[Bitwise.scala 48:55:@9441.4]
  assign _T_9389 = _T_9333 + _T_9334; // @[Bitwise.scala 48:55:@9442.4]
  assign _T_9390 = _T_9335 + _T_9336; // @[Bitwise.scala 48:55:@9443.4]
  assign _T_9391 = _T_9389 + _T_9390; // @[Bitwise.scala 48:55:@9444.4]
  assign _T_9392 = _T_9388 + _T_9391; // @[Bitwise.scala 48:55:@9445.4]
  assign _T_9393 = _T_9385 + _T_9392; // @[Bitwise.scala 48:55:@9446.4]
  assign _T_9394 = _T_9379 + _T_9393; // @[Bitwise.scala 48:55:@9447.4]
  assign _T_9395 = _T_9338 + _T_9339; // @[Bitwise.scala 48:55:@9448.4]
  assign _GEN_985 = {{1'd0}, _T_9337}; // @[Bitwise.scala 48:55:@9449.4]
  assign _T_9396 = _GEN_985 + _T_9395; // @[Bitwise.scala 48:55:@9449.4]
  assign _T_9397 = _T_9340 + _T_9341; // @[Bitwise.scala 48:55:@9450.4]
  assign _T_9398 = _T_9342 + _T_9343; // @[Bitwise.scala 48:55:@9451.4]
  assign _T_9399 = _T_9397 + _T_9398; // @[Bitwise.scala 48:55:@9452.4]
  assign _T_9400 = _T_9396 + _T_9399; // @[Bitwise.scala 48:55:@9453.4]
  assign _T_9401 = _T_9344 + _T_9345; // @[Bitwise.scala 48:55:@9454.4]
  assign _T_9402 = _T_9346 + _T_9347; // @[Bitwise.scala 48:55:@9455.4]
  assign _T_9403 = _T_9401 + _T_9402; // @[Bitwise.scala 48:55:@9456.4]
  assign _T_9404 = _T_9348 + _T_9349; // @[Bitwise.scala 48:55:@9457.4]
  assign _T_9405 = _T_9350 + _T_9351; // @[Bitwise.scala 48:55:@9458.4]
  assign _T_9406 = _T_9404 + _T_9405; // @[Bitwise.scala 48:55:@9459.4]
  assign _T_9407 = _T_9403 + _T_9406; // @[Bitwise.scala 48:55:@9460.4]
  assign _T_9408 = _T_9400 + _T_9407; // @[Bitwise.scala 48:55:@9461.4]
  assign _T_9409 = _T_9353 + _T_9354; // @[Bitwise.scala 48:55:@9462.4]
  assign _GEN_986 = {{1'd0}, _T_9352}; // @[Bitwise.scala 48:55:@9463.4]
  assign _T_9410 = _GEN_986 + _T_9409; // @[Bitwise.scala 48:55:@9463.4]
  assign _T_9411 = _T_9355 + _T_9356; // @[Bitwise.scala 48:55:@9464.4]
  assign _T_9412 = _T_9357 + _T_9358; // @[Bitwise.scala 48:55:@9465.4]
  assign _T_9413 = _T_9411 + _T_9412; // @[Bitwise.scala 48:55:@9466.4]
  assign _T_9414 = _T_9410 + _T_9413; // @[Bitwise.scala 48:55:@9467.4]
  assign _T_9415 = _T_9359 + _T_9360; // @[Bitwise.scala 48:55:@9468.4]
  assign _T_9416 = _T_9361 + _T_9362; // @[Bitwise.scala 48:55:@9469.4]
  assign _T_9417 = _T_9415 + _T_9416; // @[Bitwise.scala 48:55:@9470.4]
  assign _T_9418 = _T_9363 + _T_9364; // @[Bitwise.scala 48:55:@9471.4]
  assign _T_9419 = _T_9365 + _T_9366; // @[Bitwise.scala 48:55:@9472.4]
  assign _T_9420 = _T_9418 + _T_9419; // @[Bitwise.scala 48:55:@9473.4]
  assign _T_9421 = _T_9417 + _T_9420; // @[Bitwise.scala 48:55:@9474.4]
  assign _T_9422 = _T_9414 + _T_9421; // @[Bitwise.scala 48:55:@9475.4]
  assign _T_9423 = _T_9408 + _T_9422; // @[Bitwise.scala 48:55:@9476.4]
  assign _T_9424 = _T_9394 + _T_9423; // @[Bitwise.scala 48:55:@9477.4]
  assign _T_9488 = _T_2230[59:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@9542.4]
  assign _T_9489 = _T_9488[0]; // @[Bitwise.scala 50:65:@9543.4]
  assign _T_9490 = _T_9488[1]; // @[Bitwise.scala 50:65:@9544.4]
  assign _T_9491 = _T_9488[2]; // @[Bitwise.scala 50:65:@9545.4]
  assign _T_9492 = _T_9488[3]; // @[Bitwise.scala 50:65:@9546.4]
  assign _T_9493 = _T_9488[4]; // @[Bitwise.scala 50:65:@9547.4]
  assign _T_9494 = _T_9488[5]; // @[Bitwise.scala 50:65:@9548.4]
  assign _T_9495 = _T_9488[6]; // @[Bitwise.scala 50:65:@9549.4]
  assign _T_9496 = _T_9488[7]; // @[Bitwise.scala 50:65:@9550.4]
  assign _T_9497 = _T_9488[8]; // @[Bitwise.scala 50:65:@9551.4]
  assign _T_9498 = _T_9488[9]; // @[Bitwise.scala 50:65:@9552.4]
  assign _T_9499 = _T_9488[10]; // @[Bitwise.scala 50:65:@9553.4]
  assign _T_9500 = _T_9488[11]; // @[Bitwise.scala 50:65:@9554.4]
  assign _T_9501 = _T_9488[12]; // @[Bitwise.scala 50:65:@9555.4]
  assign _T_9502 = _T_9488[13]; // @[Bitwise.scala 50:65:@9556.4]
  assign _T_9503 = _T_9488[14]; // @[Bitwise.scala 50:65:@9557.4]
  assign _T_9504 = _T_9488[15]; // @[Bitwise.scala 50:65:@9558.4]
  assign _T_9505 = _T_9488[16]; // @[Bitwise.scala 50:65:@9559.4]
  assign _T_9506 = _T_9488[17]; // @[Bitwise.scala 50:65:@9560.4]
  assign _T_9507 = _T_9488[18]; // @[Bitwise.scala 50:65:@9561.4]
  assign _T_9508 = _T_9488[19]; // @[Bitwise.scala 50:65:@9562.4]
  assign _T_9509 = _T_9488[20]; // @[Bitwise.scala 50:65:@9563.4]
  assign _T_9510 = _T_9488[21]; // @[Bitwise.scala 50:65:@9564.4]
  assign _T_9511 = _T_9488[22]; // @[Bitwise.scala 50:65:@9565.4]
  assign _T_9512 = _T_9488[23]; // @[Bitwise.scala 50:65:@9566.4]
  assign _T_9513 = _T_9488[24]; // @[Bitwise.scala 50:65:@9567.4]
  assign _T_9514 = _T_9488[25]; // @[Bitwise.scala 50:65:@9568.4]
  assign _T_9515 = _T_9488[26]; // @[Bitwise.scala 50:65:@9569.4]
  assign _T_9516 = _T_9488[27]; // @[Bitwise.scala 50:65:@9570.4]
  assign _T_9517 = _T_9488[28]; // @[Bitwise.scala 50:65:@9571.4]
  assign _T_9518 = _T_9488[29]; // @[Bitwise.scala 50:65:@9572.4]
  assign _T_9519 = _T_9488[30]; // @[Bitwise.scala 50:65:@9573.4]
  assign _T_9520 = _T_9488[31]; // @[Bitwise.scala 50:65:@9574.4]
  assign _T_9521 = _T_9488[32]; // @[Bitwise.scala 50:65:@9575.4]
  assign _T_9522 = _T_9488[33]; // @[Bitwise.scala 50:65:@9576.4]
  assign _T_9523 = _T_9488[34]; // @[Bitwise.scala 50:65:@9577.4]
  assign _T_9524 = _T_9488[35]; // @[Bitwise.scala 50:65:@9578.4]
  assign _T_9525 = _T_9488[36]; // @[Bitwise.scala 50:65:@9579.4]
  assign _T_9526 = _T_9488[37]; // @[Bitwise.scala 50:65:@9580.4]
  assign _T_9527 = _T_9488[38]; // @[Bitwise.scala 50:65:@9581.4]
  assign _T_9528 = _T_9488[39]; // @[Bitwise.scala 50:65:@9582.4]
  assign _T_9529 = _T_9488[40]; // @[Bitwise.scala 50:65:@9583.4]
  assign _T_9530 = _T_9488[41]; // @[Bitwise.scala 50:65:@9584.4]
  assign _T_9531 = _T_9488[42]; // @[Bitwise.scala 50:65:@9585.4]
  assign _T_9532 = _T_9488[43]; // @[Bitwise.scala 50:65:@9586.4]
  assign _T_9533 = _T_9488[44]; // @[Bitwise.scala 50:65:@9587.4]
  assign _T_9534 = _T_9488[45]; // @[Bitwise.scala 50:65:@9588.4]
  assign _T_9535 = _T_9488[46]; // @[Bitwise.scala 50:65:@9589.4]
  assign _T_9536 = _T_9488[47]; // @[Bitwise.scala 50:65:@9590.4]
  assign _T_9537 = _T_9488[48]; // @[Bitwise.scala 50:65:@9591.4]
  assign _T_9538 = _T_9488[49]; // @[Bitwise.scala 50:65:@9592.4]
  assign _T_9539 = _T_9488[50]; // @[Bitwise.scala 50:65:@9593.4]
  assign _T_9540 = _T_9488[51]; // @[Bitwise.scala 50:65:@9594.4]
  assign _T_9541 = _T_9488[52]; // @[Bitwise.scala 50:65:@9595.4]
  assign _T_9542 = _T_9488[53]; // @[Bitwise.scala 50:65:@9596.4]
  assign _T_9543 = _T_9488[54]; // @[Bitwise.scala 50:65:@9597.4]
  assign _T_9544 = _T_9488[55]; // @[Bitwise.scala 50:65:@9598.4]
  assign _T_9545 = _T_9488[56]; // @[Bitwise.scala 50:65:@9599.4]
  assign _T_9546 = _T_9488[57]; // @[Bitwise.scala 50:65:@9600.4]
  assign _T_9547 = _T_9488[58]; // @[Bitwise.scala 50:65:@9601.4]
  assign _T_9548 = _T_9488[59]; // @[Bitwise.scala 50:65:@9602.4]
  assign _T_9549 = _T_9490 + _T_9491; // @[Bitwise.scala 48:55:@9603.4]
  assign _GEN_987 = {{1'd0}, _T_9489}; // @[Bitwise.scala 48:55:@9604.4]
  assign _T_9550 = _GEN_987 + _T_9549; // @[Bitwise.scala 48:55:@9604.4]
  assign _T_9551 = _T_9492 + _T_9493; // @[Bitwise.scala 48:55:@9605.4]
  assign _T_9552 = _T_9494 + _T_9495; // @[Bitwise.scala 48:55:@9606.4]
  assign _T_9553 = _T_9551 + _T_9552; // @[Bitwise.scala 48:55:@9607.4]
  assign _T_9554 = _T_9550 + _T_9553; // @[Bitwise.scala 48:55:@9608.4]
  assign _T_9555 = _T_9496 + _T_9497; // @[Bitwise.scala 48:55:@9609.4]
  assign _T_9556 = _T_9498 + _T_9499; // @[Bitwise.scala 48:55:@9610.4]
  assign _T_9557 = _T_9555 + _T_9556; // @[Bitwise.scala 48:55:@9611.4]
  assign _T_9558 = _T_9500 + _T_9501; // @[Bitwise.scala 48:55:@9612.4]
  assign _T_9559 = _T_9502 + _T_9503; // @[Bitwise.scala 48:55:@9613.4]
  assign _T_9560 = _T_9558 + _T_9559; // @[Bitwise.scala 48:55:@9614.4]
  assign _T_9561 = _T_9557 + _T_9560; // @[Bitwise.scala 48:55:@9615.4]
  assign _T_9562 = _T_9554 + _T_9561; // @[Bitwise.scala 48:55:@9616.4]
  assign _T_9563 = _T_9505 + _T_9506; // @[Bitwise.scala 48:55:@9617.4]
  assign _GEN_988 = {{1'd0}, _T_9504}; // @[Bitwise.scala 48:55:@9618.4]
  assign _T_9564 = _GEN_988 + _T_9563; // @[Bitwise.scala 48:55:@9618.4]
  assign _T_9565 = _T_9507 + _T_9508; // @[Bitwise.scala 48:55:@9619.4]
  assign _T_9566 = _T_9509 + _T_9510; // @[Bitwise.scala 48:55:@9620.4]
  assign _T_9567 = _T_9565 + _T_9566; // @[Bitwise.scala 48:55:@9621.4]
  assign _T_9568 = _T_9564 + _T_9567; // @[Bitwise.scala 48:55:@9622.4]
  assign _T_9569 = _T_9511 + _T_9512; // @[Bitwise.scala 48:55:@9623.4]
  assign _T_9570 = _T_9513 + _T_9514; // @[Bitwise.scala 48:55:@9624.4]
  assign _T_9571 = _T_9569 + _T_9570; // @[Bitwise.scala 48:55:@9625.4]
  assign _T_9572 = _T_9515 + _T_9516; // @[Bitwise.scala 48:55:@9626.4]
  assign _T_9573 = _T_9517 + _T_9518; // @[Bitwise.scala 48:55:@9627.4]
  assign _T_9574 = _T_9572 + _T_9573; // @[Bitwise.scala 48:55:@9628.4]
  assign _T_9575 = _T_9571 + _T_9574; // @[Bitwise.scala 48:55:@9629.4]
  assign _T_9576 = _T_9568 + _T_9575; // @[Bitwise.scala 48:55:@9630.4]
  assign _T_9577 = _T_9562 + _T_9576; // @[Bitwise.scala 48:55:@9631.4]
  assign _T_9578 = _T_9520 + _T_9521; // @[Bitwise.scala 48:55:@9632.4]
  assign _GEN_989 = {{1'd0}, _T_9519}; // @[Bitwise.scala 48:55:@9633.4]
  assign _T_9579 = _GEN_989 + _T_9578; // @[Bitwise.scala 48:55:@9633.4]
  assign _T_9580 = _T_9522 + _T_9523; // @[Bitwise.scala 48:55:@9634.4]
  assign _T_9581 = _T_9524 + _T_9525; // @[Bitwise.scala 48:55:@9635.4]
  assign _T_9582 = _T_9580 + _T_9581; // @[Bitwise.scala 48:55:@9636.4]
  assign _T_9583 = _T_9579 + _T_9582; // @[Bitwise.scala 48:55:@9637.4]
  assign _T_9584 = _T_9526 + _T_9527; // @[Bitwise.scala 48:55:@9638.4]
  assign _T_9585 = _T_9528 + _T_9529; // @[Bitwise.scala 48:55:@9639.4]
  assign _T_9586 = _T_9584 + _T_9585; // @[Bitwise.scala 48:55:@9640.4]
  assign _T_9587 = _T_9530 + _T_9531; // @[Bitwise.scala 48:55:@9641.4]
  assign _T_9588 = _T_9532 + _T_9533; // @[Bitwise.scala 48:55:@9642.4]
  assign _T_9589 = _T_9587 + _T_9588; // @[Bitwise.scala 48:55:@9643.4]
  assign _T_9590 = _T_9586 + _T_9589; // @[Bitwise.scala 48:55:@9644.4]
  assign _T_9591 = _T_9583 + _T_9590; // @[Bitwise.scala 48:55:@9645.4]
  assign _T_9592 = _T_9535 + _T_9536; // @[Bitwise.scala 48:55:@9646.4]
  assign _GEN_990 = {{1'd0}, _T_9534}; // @[Bitwise.scala 48:55:@9647.4]
  assign _T_9593 = _GEN_990 + _T_9592; // @[Bitwise.scala 48:55:@9647.4]
  assign _T_9594 = _T_9537 + _T_9538; // @[Bitwise.scala 48:55:@9648.4]
  assign _T_9595 = _T_9539 + _T_9540; // @[Bitwise.scala 48:55:@9649.4]
  assign _T_9596 = _T_9594 + _T_9595; // @[Bitwise.scala 48:55:@9650.4]
  assign _T_9597 = _T_9593 + _T_9596; // @[Bitwise.scala 48:55:@9651.4]
  assign _T_9598 = _T_9541 + _T_9542; // @[Bitwise.scala 48:55:@9652.4]
  assign _T_9599 = _T_9543 + _T_9544; // @[Bitwise.scala 48:55:@9653.4]
  assign _T_9600 = _T_9598 + _T_9599; // @[Bitwise.scala 48:55:@9654.4]
  assign _T_9601 = _T_9545 + _T_9546; // @[Bitwise.scala 48:55:@9655.4]
  assign _T_9602 = _T_9547 + _T_9548; // @[Bitwise.scala 48:55:@9656.4]
  assign _T_9603 = _T_9601 + _T_9602; // @[Bitwise.scala 48:55:@9657.4]
  assign _T_9604 = _T_9600 + _T_9603; // @[Bitwise.scala 48:55:@9658.4]
  assign _T_9605 = _T_9597 + _T_9604; // @[Bitwise.scala 48:55:@9659.4]
  assign _T_9606 = _T_9591 + _T_9605; // @[Bitwise.scala 48:55:@9660.4]
  assign _T_9607 = _T_9577 + _T_9606; // @[Bitwise.scala 48:55:@9661.4]
  assign _T_9671 = _T_2230[60:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@9726.4]
  assign _T_9672 = _T_9671[0]; // @[Bitwise.scala 50:65:@9727.4]
  assign _T_9673 = _T_9671[1]; // @[Bitwise.scala 50:65:@9728.4]
  assign _T_9674 = _T_9671[2]; // @[Bitwise.scala 50:65:@9729.4]
  assign _T_9675 = _T_9671[3]; // @[Bitwise.scala 50:65:@9730.4]
  assign _T_9676 = _T_9671[4]; // @[Bitwise.scala 50:65:@9731.4]
  assign _T_9677 = _T_9671[5]; // @[Bitwise.scala 50:65:@9732.4]
  assign _T_9678 = _T_9671[6]; // @[Bitwise.scala 50:65:@9733.4]
  assign _T_9679 = _T_9671[7]; // @[Bitwise.scala 50:65:@9734.4]
  assign _T_9680 = _T_9671[8]; // @[Bitwise.scala 50:65:@9735.4]
  assign _T_9681 = _T_9671[9]; // @[Bitwise.scala 50:65:@9736.4]
  assign _T_9682 = _T_9671[10]; // @[Bitwise.scala 50:65:@9737.4]
  assign _T_9683 = _T_9671[11]; // @[Bitwise.scala 50:65:@9738.4]
  assign _T_9684 = _T_9671[12]; // @[Bitwise.scala 50:65:@9739.4]
  assign _T_9685 = _T_9671[13]; // @[Bitwise.scala 50:65:@9740.4]
  assign _T_9686 = _T_9671[14]; // @[Bitwise.scala 50:65:@9741.4]
  assign _T_9687 = _T_9671[15]; // @[Bitwise.scala 50:65:@9742.4]
  assign _T_9688 = _T_9671[16]; // @[Bitwise.scala 50:65:@9743.4]
  assign _T_9689 = _T_9671[17]; // @[Bitwise.scala 50:65:@9744.4]
  assign _T_9690 = _T_9671[18]; // @[Bitwise.scala 50:65:@9745.4]
  assign _T_9691 = _T_9671[19]; // @[Bitwise.scala 50:65:@9746.4]
  assign _T_9692 = _T_9671[20]; // @[Bitwise.scala 50:65:@9747.4]
  assign _T_9693 = _T_9671[21]; // @[Bitwise.scala 50:65:@9748.4]
  assign _T_9694 = _T_9671[22]; // @[Bitwise.scala 50:65:@9749.4]
  assign _T_9695 = _T_9671[23]; // @[Bitwise.scala 50:65:@9750.4]
  assign _T_9696 = _T_9671[24]; // @[Bitwise.scala 50:65:@9751.4]
  assign _T_9697 = _T_9671[25]; // @[Bitwise.scala 50:65:@9752.4]
  assign _T_9698 = _T_9671[26]; // @[Bitwise.scala 50:65:@9753.4]
  assign _T_9699 = _T_9671[27]; // @[Bitwise.scala 50:65:@9754.4]
  assign _T_9700 = _T_9671[28]; // @[Bitwise.scala 50:65:@9755.4]
  assign _T_9701 = _T_9671[29]; // @[Bitwise.scala 50:65:@9756.4]
  assign _T_9702 = _T_9671[30]; // @[Bitwise.scala 50:65:@9757.4]
  assign _T_9703 = _T_9671[31]; // @[Bitwise.scala 50:65:@9758.4]
  assign _T_9704 = _T_9671[32]; // @[Bitwise.scala 50:65:@9759.4]
  assign _T_9705 = _T_9671[33]; // @[Bitwise.scala 50:65:@9760.4]
  assign _T_9706 = _T_9671[34]; // @[Bitwise.scala 50:65:@9761.4]
  assign _T_9707 = _T_9671[35]; // @[Bitwise.scala 50:65:@9762.4]
  assign _T_9708 = _T_9671[36]; // @[Bitwise.scala 50:65:@9763.4]
  assign _T_9709 = _T_9671[37]; // @[Bitwise.scala 50:65:@9764.4]
  assign _T_9710 = _T_9671[38]; // @[Bitwise.scala 50:65:@9765.4]
  assign _T_9711 = _T_9671[39]; // @[Bitwise.scala 50:65:@9766.4]
  assign _T_9712 = _T_9671[40]; // @[Bitwise.scala 50:65:@9767.4]
  assign _T_9713 = _T_9671[41]; // @[Bitwise.scala 50:65:@9768.4]
  assign _T_9714 = _T_9671[42]; // @[Bitwise.scala 50:65:@9769.4]
  assign _T_9715 = _T_9671[43]; // @[Bitwise.scala 50:65:@9770.4]
  assign _T_9716 = _T_9671[44]; // @[Bitwise.scala 50:65:@9771.4]
  assign _T_9717 = _T_9671[45]; // @[Bitwise.scala 50:65:@9772.4]
  assign _T_9718 = _T_9671[46]; // @[Bitwise.scala 50:65:@9773.4]
  assign _T_9719 = _T_9671[47]; // @[Bitwise.scala 50:65:@9774.4]
  assign _T_9720 = _T_9671[48]; // @[Bitwise.scala 50:65:@9775.4]
  assign _T_9721 = _T_9671[49]; // @[Bitwise.scala 50:65:@9776.4]
  assign _T_9722 = _T_9671[50]; // @[Bitwise.scala 50:65:@9777.4]
  assign _T_9723 = _T_9671[51]; // @[Bitwise.scala 50:65:@9778.4]
  assign _T_9724 = _T_9671[52]; // @[Bitwise.scala 50:65:@9779.4]
  assign _T_9725 = _T_9671[53]; // @[Bitwise.scala 50:65:@9780.4]
  assign _T_9726 = _T_9671[54]; // @[Bitwise.scala 50:65:@9781.4]
  assign _T_9727 = _T_9671[55]; // @[Bitwise.scala 50:65:@9782.4]
  assign _T_9728 = _T_9671[56]; // @[Bitwise.scala 50:65:@9783.4]
  assign _T_9729 = _T_9671[57]; // @[Bitwise.scala 50:65:@9784.4]
  assign _T_9730 = _T_9671[58]; // @[Bitwise.scala 50:65:@9785.4]
  assign _T_9731 = _T_9671[59]; // @[Bitwise.scala 50:65:@9786.4]
  assign _T_9732 = _T_9671[60]; // @[Bitwise.scala 50:65:@9787.4]
  assign _T_9733 = _T_9673 + _T_9674; // @[Bitwise.scala 48:55:@9788.4]
  assign _GEN_991 = {{1'd0}, _T_9672}; // @[Bitwise.scala 48:55:@9789.4]
  assign _T_9734 = _GEN_991 + _T_9733; // @[Bitwise.scala 48:55:@9789.4]
  assign _T_9735 = _T_9675 + _T_9676; // @[Bitwise.scala 48:55:@9790.4]
  assign _T_9736 = _T_9677 + _T_9678; // @[Bitwise.scala 48:55:@9791.4]
  assign _T_9737 = _T_9735 + _T_9736; // @[Bitwise.scala 48:55:@9792.4]
  assign _T_9738 = _T_9734 + _T_9737; // @[Bitwise.scala 48:55:@9793.4]
  assign _T_9739 = _T_9679 + _T_9680; // @[Bitwise.scala 48:55:@9794.4]
  assign _T_9740 = _T_9681 + _T_9682; // @[Bitwise.scala 48:55:@9795.4]
  assign _T_9741 = _T_9739 + _T_9740; // @[Bitwise.scala 48:55:@9796.4]
  assign _T_9742 = _T_9683 + _T_9684; // @[Bitwise.scala 48:55:@9797.4]
  assign _T_9743 = _T_9685 + _T_9686; // @[Bitwise.scala 48:55:@9798.4]
  assign _T_9744 = _T_9742 + _T_9743; // @[Bitwise.scala 48:55:@9799.4]
  assign _T_9745 = _T_9741 + _T_9744; // @[Bitwise.scala 48:55:@9800.4]
  assign _T_9746 = _T_9738 + _T_9745; // @[Bitwise.scala 48:55:@9801.4]
  assign _T_9747 = _T_9688 + _T_9689; // @[Bitwise.scala 48:55:@9802.4]
  assign _GEN_992 = {{1'd0}, _T_9687}; // @[Bitwise.scala 48:55:@9803.4]
  assign _T_9748 = _GEN_992 + _T_9747; // @[Bitwise.scala 48:55:@9803.4]
  assign _T_9749 = _T_9690 + _T_9691; // @[Bitwise.scala 48:55:@9804.4]
  assign _T_9750 = _T_9692 + _T_9693; // @[Bitwise.scala 48:55:@9805.4]
  assign _T_9751 = _T_9749 + _T_9750; // @[Bitwise.scala 48:55:@9806.4]
  assign _T_9752 = _T_9748 + _T_9751; // @[Bitwise.scala 48:55:@9807.4]
  assign _T_9753 = _T_9694 + _T_9695; // @[Bitwise.scala 48:55:@9808.4]
  assign _T_9754 = _T_9696 + _T_9697; // @[Bitwise.scala 48:55:@9809.4]
  assign _T_9755 = _T_9753 + _T_9754; // @[Bitwise.scala 48:55:@9810.4]
  assign _T_9756 = _T_9698 + _T_9699; // @[Bitwise.scala 48:55:@9811.4]
  assign _T_9757 = _T_9700 + _T_9701; // @[Bitwise.scala 48:55:@9812.4]
  assign _T_9758 = _T_9756 + _T_9757; // @[Bitwise.scala 48:55:@9813.4]
  assign _T_9759 = _T_9755 + _T_9758; // @[Bitwise.scala 48:55:@9814.4]
  assign _T_9760 = _T_9752 + _T_9759; // @[Bitwise.scala 48:55:@9815.4]
  assign _T_9761 = _T_9746 + _T_9760; // @[Bitwise.scala 48:55:@9816.4]
  assign _T_9762 = _T_9703 + _T_9704; // @[Bitwise.scala 48:55:@9817.4]
  assign _GEN_993 = {{1'd0}, _T_9702}; // @[Bitwise.scala 48:55:@9818.4]
  assign _T_9763 = _GEN_993 + _T_9762; // @[Bitwise.scala 48:55:@9818.4]
  assign _T_9764 = _T_9705 + _T_9706; // @[Bitwise.scala 48:55:@9819.4]
  assign _T_9765 = _T_9707 + _T_9708; // @[Bitwise.scala 48:55:@9820.4]
  assign _T_9766 = _T_9764 + _T_9765; // @[Bitwise.scala 48:55:@9821.4]
  assign _T_9767 = _T_9763 + _T_9766; // @[Bitwise.scala 48:55:@9822.4]
  assign _T_9768 = _T_9709 + _T_9710; // @[Bitwise.scala 48:55:@9823.4]
  assign _T_9769 = _T_9711 + _T_9712; // @[Bitwise.scala 48:55:@9824.4]
  assign _T_9770 = _T_9768 + _T_9769; // @[Bitwise.scala 48:55:@9825.4]
  assign _T_9771 = _T_9713 + _T_9714; // @[Bitwise.scala 48:55:@9826.4]
  assign _T_9772 = _T_9715 + _T_9716; // @[Bitwise.scala 48:55:@9827.4]
  assign _T_9773 = _T_9771 + _T_9772; // @[Bitwise.scala 48:55:@9828.4]
  assign _T_9774 = _T_9770 + _T_9773; // @[Bitwise.scala 48:55:@9829.4]
  assign _T_9775 = _T_9767 + _T_9774; // @[Bitwise.scala 48:55:@9830.4]
  assign _T_9776 = _T_9717 + _T_9718; // @[Bitwise.scala 48:55:@9831.4]
  assign _T_9777 = _T_9719 + _T_9720; // @[Bitwise.scala 48:55:@9832.4]
  assign _T_9778 = _T_9776 + _T_9777; // @[Bitwise.scala 48:55:@9833.4]
  assign _T_9779 = _T_9721 + _T_9722; // @[Bitwise.scala 48:55:@9834.4]
  assign _T_9780 = _T_9723 + _T_9724; // @[Bitwise.scala 48:55:@9835.4]
  assign _T_9781 = _T_9779 + _T_9780; // @[Bitwise.scala 48:55:@9836.4]
  assign _T_9782 = _T_9778 + _T_9781; // @[Bitwise.scala 48:55:@9837.4]
  assign _T_9783 = _T_9725 + _T_9726; // @[Bitwise.scala 48:55:@9838.4]
  assign _T_9784 = _T_9727 + _T_9728; // @[Bitwise.scala 48:55:@9839.4]
  assign _T_9785 = _T_9783 + _T_9784; // @[Bitwise.scala 48:55:@9840.4]
  assign _T_9786 = _T_9729 + _T_9730; // @[Bitwise.scala 48:55:@9841.4]
  assign _T_9787 = _T_9731 + _T_9732; // @[Bitwise.scala 48:55:@9842.4]
  assign _T_9788 = _T_9786 + _T_9787; // @[Bitwise.scala 48:55:@9843.4]
  assign _T_9789 = _T_9785 + _T_9788; // @[Bitwise.scala 48:55:@9844.4]
  assign _T_9790 = _T_9782 + _T_9789; // @[Bitwise.scala 48:55:@9845.4]
  assign _T_9791 = _T_9775 + _T_9790; // @[Bitwise.scala 48:55:@9846.4]
  assign _T_9792 = _T_9761 + _T_9791; // @[Bitwise.scala 48:55:@9847.4]
  assign _T_9856 = _T_2230[61:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@9912.4]
  assign _T_9857 = _T_9856[0]; // @[Bitwise.scala 50:65:@9913.4]
  assign _T_9858 = _T_9856[1]; // @[Bitwise.scala 50:65:@9914.4]
  assign _T_9859 = _T_9856[2]; // @[Bitwise.scala 50:65:@9915.4]
  assign _T_9860 = _T_9856[3]; // @[Bitwise.scala 50:65:@9916.4]
  assign _T_9861 = _T_9856[4]; // @[Bitwise.scala 50:65:@9917.4]
  assign _T_9862 = _T_9856[5]; // @[Bitwise.scala 50:65:@9918.4]
  assign _T_9863 = _T_9856[6]; // @[Bitwise.scala 50:65:@9919.4]
  assign _T_9864 = _T_9856[7]; // @[Bitwise.scala 50:65:@9920.4]
  assign _T_9865 = _T_9856[8]; // @[Bitwise.scala 50:65:@9921.4]
  assign _T_9866 = _T_9856[9]; // @[Bitwise.scala 50:65:@9922.4]
  assign _T_9867 = _T_9856[10]; // @[Bitwise.scala 50:65:@9923.4]
  assign _T_9868 = _T_9856[11]; // @[Bitwise.scala 50:65:@9924.4]
  assign _T_9869 = _T_9856[12]; // @[Bitwise.scala 50:65:@9925.4]
  assign _T_9870 = _T_9856[13]; // @[Bitwise.scala 50:65:@9926.4]
  assign _T_9871 = _T_9856[14]; // @[Bitwise.scala 50:65:@9927.4]
  assign _T_9872 = _T_9856[15]; // @[Bitwise.scala 50:65:@9928.4]
  assign _T_9873 = _T_9856[16]; // @[Bitwise.scala 50:65:@9929.4]
  assign _T_9874 = _T_9856[17]; // @[Bitwise.scala 50:65:@9930.4]
  assign _T_9875 = _T_9856[18]; // @[Bitwise.scala 50:65:@9931.4]
  assign _T_9876 = _T_9856[19]; // @[Bitwise.scala 50:65:@9932.4]
  assign _T_9877 = _T_9856[20]; // @[Bitwise.scala 50:65:@9933.4]
  assign _T_9878 = _T_9856[21]; // @[Bitwise.scala 50:65:@9934.4]
  assign _T_9879 = _T_9856[22]; // @[Bitwise.scala 50:65:@9935.4]
  assign _T_9880 = _T_9856[23]; // @[Bitwise.scala 50:65:@9936.4]
  assign _T_9881 = _T_9856[24]; // @[Bitwise.scala 50:65:@9937.4]
  assign _T_9882 = _T_9856[25]; // @[Bitwise.scala 50:65:@9938.4]
  assign _T_9883 = _T_9856[26]; // @[Bitwise.scala 50:65:@9939.4]
  assign _T_9884 = _T_9856[27]; // @[Bitwise.scala 50:65:@9940.4]
  assign _T_9885 = _T_9856[28]; // @[Bitwise.scala 50:65:@9941.4]
  assign _T_9886 = _T_9856[29]; // @[Bitwise.scala 50:65:@9942.4]
  assign _T_9887 = _T_9856[30]; // @[Bitwise.scala 50:65:@9943.4]
  assign _T_9888 = _T_9856[31]; // @[Bitwise.scala 50:65:@9944.4]
  assign _T_9889 = _T_9856[32]; // @[Bitwise.scala 50:65:@9945.4]
  assign _T_9890 = _T_9856[33]; // @[Bitwise.scala 50:65:@9946.4]
  assign _T_9891 = _T_9856[34]; // @[Bitwise.scala 50:65:@9947.4]
  assign _T_9892 = _T_9856[35]; // @[Bitwise.scala 50:65:@9948.4]
  assign _T_9893 = _T_9856[36]; // @[Bitwise.scala 50:65:@9949.4]
  assign _T_9894 = _T_9856[37]; // @[Bitwise.scala 50:65:@9950.4]
  assign _T_9895 = _T_9856[38]; // @[Bitwise.scala 50:65:@9951.4]
  assign _T_9896 = _T_9856[39]; // @[Bitwise.scala 50:65:@9952.4]
  assign _T_9897 = _T_9856[40]; // @[Bitwise.scala 50:65:@9953.4]
  assign _T_9898 = _T_9856[41]; // @[Bitwise.scala 50:65:@9954.4]
  assign _T_9899 = _T_9856[42]; // @[Bitwise.scala 50:65:@9955.4]
  assign _T_9900 = _T_9856[43]; // @[Bitwise.scala 50:65:@9956.4]
  assign _T_9901 = _T_9856[44]; // @[Bitwise.scala 50:65:@9957.4]
  assign _T_9902 = _T_9856[45]; // @[Bitwise.scala 50:65:@9958.4]
  assign _T_9903 = _T_9856[46]; // @[Bitwise.scala 50:65:@9959.4]
  assign _T_9904 = _T_9856[47]; // @[Bitwise.scala 50:65:@9960.4]
  assign _T_9905 = _T_9856[48]; // @[Bitwise.scala 50:65:@9961.4]
  assign _T_9906 = _T_9856[49]; // @[Bitwise.scala 50:65:@9962.4]
  assign _T_9907 = _T_9856[50]; // @[Bitwise.scala 50:65:@9963.4]
  assign _T_9908 = _T_9856[51]; // @[Bitwise.scala 50:65:@9964.4]
  assign _T_9909 = _T_9856[52]; // @[Bitwise.scala 50:65:@9965.4]
  assign _T_9910 = _T_9856[53]; // @[Bitwise.scala 50:65:@9966.4]
  assign _T_9911 = _T_9856[54]; // @[Bitwise.scala 50:65:@9967.4]
  assign _T_9912 = _T_9856[55]; // @[Bitwise.scala 50:65:@9968.4]
  assign _T_9913 = _T_9856[56]; // @[Bitwise.scala 50:65:@9969.4]
  assign _T_9914 = _T_9856[57]; // @[Bitwise.scala 50:65:@9970.4]
  assign _T_9915 = _T_9856[58]; // @[Bitwise.scala 50:65:@9971.4]
  assign _T_9916 = _T_9856[59]; // @[Bitwise.scala 50:65:@9972.4]
  assign _T_9917 = _T_9856[60]; // @[Bitwise.scala 50:65:@9973.4]
  assign _T_9918 = _T_9856[61]; // @[Bitwise.scala 50:65:@9974.4]
  assign _T_9919 = _T_9858 + _T_9859; // @[Bitwise.scala 48:55:@9975.4]
  assign _GEN_994 = {{1'd0}, _T_9857}; // @[Bitwise.scala 48:55:@9976.4]
  assign _T_9920 = _GEN_994 + _T_9919; // @[Bitwise.scala 48:55:@9976.4]
  assign _T_9921 = _T_9860 + _T_9861; // @[Bitwise.scala 48:55:@9977.4]
  assign _T_9922 = _T_9862 + _T_9863; // @[Bitwise.scala 48:55:@9978.4]
  assign _T_9923 = _T_9921 + _T_9922; // @[Bitwise.scala 48:55:@9979.4]
  assign _T_9924 = _T_9920 + _T_9923; // @[Bitwise.scala 48:55:@9980.4]
  assign _T_9925 = _T_9864 + _T_9865; // @[Bitwise.scala 48:55:@9981.4]
  assign _T_9926 = _T_9866 + _T_9867; // @[Bitwise.scala 48:55:@9982.4]
  assign _T_9927 = _T_9925 + _T_9926; // @[Bitwise.scala 48:55:@9983.4]
  assign _T_9928 = _T_9868 + _T_9869; // @[Bitwise.scala 48:55:@9984.4]
  assign _T_9929 = _T_9870 + _T_9871; // @[Bitwise.scala 48:55:@9985.4]
  assign _T_9930 = _T_9928 + _T_9929; // @[Bitwise.scala 48:55:@9986.4]
  assign _T_9931 = _T_9927 + _T_9930; // @[Bitwise.scala 48:55:@9987.4]
  assign _T_9932 = _T_9924 + _T_9931; // @[Bitwise.scala 48:55:@9988.4]
  assign _T_9933 = _T_9872 + _T_9873; // @[Bitwise.scala 48:55:@9989.4]
  assign _T_9934 = _T_9874 + _T_9875; // @[Bitwise.scala 48:55:@9990.4]
  assign _T_9935 = _T_9933 + _T_9934; // @[Bitwise.scala 48:55:@9991.4]
  assign _T_9936 = _T_9876 + _T_9877; // @[Bitwise.scala 48:55:@9992.4]
  assign _T_9937 = _T_9878 + _T_9879; // @[Bitwise.scala 48:55:@9993.4]
  assign _T_9938 = _T_9936 + _T_9937; // @[Bitwise.scala 48:55:@9994.4]
  assign _T_9939 = _T_9935 + _T_9938; // @[Bitwise.scala 48:55:@9995.4]
  assign _T_9940 = _T_9880 + _T_9881; // @[Bitwise.scala 48:55:@9996.4]
  assign _T_9941 = _T_9882 + _T_9883; // @[Bitwise.scala 48:55:@9997.4]
  assign _T_9942 = _T_9940 + _T_9941; // @[Bitwise.scala 48:55:@9998.4]
  assign _T_9943 = _T_9884 + _T_9885; // @[Bitwise.scala 48:55:@9999.4]
  assign _T_9944 = _T_9886 + _T_9887; // @[Bitwise.scala 48:55:@10000.4]
  assign _T_9945 = _T_9943 + _T_9944; // @[Bitwise.scala 48:55:@10001.4]
  assign _T_9946 = _T_9942 + _T_9945; // @[Bitwise.scala 48:55:@10002.4]
  assign _T_9947 = _T_9939 + _T_9946; // @[Bitwise.scala 48:55:@10003.4]
  assign _T_9948 = _T_9932 + _T_9947; // @[Bitwise.scala 48:55:@10004.4]
  assign _T_9949 = _T_9889 + _T_9890; // @[Bitwise.scala 48:55:@10005.4]
  assign _GEN_995 = {{1'd0}, _T_9888}; // @[Bitwise.scala 48:55:@10006.4]
  assign _T_9950 = _GEN_995 + _T_9949; // @[Bitwise.scala 48:55:@10006.4]
  assign _T_9951 = _T_9891 + _T_9892; // @[Bitwise.scala 48:55:@10007.4]
  assign _T_9952 = _T_9893 + _T_9894; // @[Bitwise.scala 48:55:@10008.4]
  assign _T_9953 = _T_9951 + _T_9952; // @[Bitwise.scala 48:55:@10009.4]
  assign _T_9954 = _T_9950 + _T_9953; // @[Bitwise.scala 48:55:@10010.4]
  assign _T_9955 = _T_9895 + _T_9896; // @[Bitwise.scala 48:55:@10011.4]
  assign _T_9956 = _T_9897 + _T_9898; // @[Bitwise.scala 48:55:@10012.4]
  assign _T_9957 = _T_9955 + _T_9956; // @[Bitwise.scala 48:55:@10013.4]
  assign _T_9958 = _T_9899 + _T_9900; // @[Bitwise.scala 48:55:@10014.4]
  assign _T_9959 = _T_9901 + _T_9902; // @[Bitwise.scala 48:55:@10015.4]
  assign _T_9960 = _T_9958 + _T_9959; // @[Bitwise.scala 48:55:@10016.4]
  assign _T_9961 = _T_9957 + _T_9960; // @[Bitwise.scala 48:55:@10017.4]
  assign _T_9962 = _T_9954 + _T_9961; // @[Bitwise.scala 48:55:@10018.4]
  assign _T_9963 = _T_9903 + _T_9904; // @[Bitwise.scala 48:55:@10019.4]
  assign _T_9964 = _T_9905 + _T_9906; // @[Bitwise.scala 48:55:@10020.4]
  assign _T_9965 = _T_9963 + _T_9964; // @[Bitwise.scala 48:55:@10021.4]
  assign _T_9966 = _T_9907 + _T_9908; // @[Bitwise.scala 48:55:@10022.4]
  assign _T_9967 = _T_9909 + _T_9910; // @[Bitwise.scala 48:55:@10023.4]
  assign _T_9968 = _T_9966 + _T_9967; // @[Bitwise.scala 48:55:@10024.4]
  assign _T_9969 = _T_9965 + _T_9968; // @[Bitwise.scala 48:55:@10025.4]
  assign _T_9970 = _T_9911 + _T_9912; // @[Bitwise.scala 48:55:@10026.4]
  assign _T_9971 = _T_9913 + _T_9914; // @[Bitwise.scala 48:55:@10027.4]
  assign _T_9972 = _T_9970 + _T_9971; // @[Bitwise.scala 48:55:@10028.4]
  assign _T_9973 = _T_9915 + _T_9916; // @[Bitwise.scala 48:55:@10029.4]
  assign _T_9974 = _T_9917 + _T_9918; // @[Bitwise.scala 48:55:@10030.4]
  assign _T_9975 = _T_9973 + _T_9974; // @[Bitwise.scala 48:55:@10031.4]
  assign _T_9976 = _T_9972 + _T_9975; // @[Bitwise.scala 48:55:@10032.4]
  assign _T_9977 = _T_9969 + _T_9976; // @[Bitwise.scala 48:55:@10033.4]
  assign _T_9978 = _T_9962 + _T_9977; // @[Bitwise.scala 48:55:@10034.4]
  assign _T_9979 = _T_9948 + _T_9978; // @[Bitwise.scala 48:55:@10035.4]
  assign _T_10043 = _T_2230[62:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@10100.4]
  assign _T_10044 = _T_10043[0]; // @[Bitwise.scala 50:65:@10101.4]
  assign _T_10045 = _T_10043[1]; // @[Bitwise.scala 50:65:@10102.4]
  assign _T_10046 = _T_10043[2]; // @[Bitwise.scala 50:65:@10103.4]
  assign _T_10047 = _T_10043[3]; // @[Bitwise.scala 50:65:@10104.4]
  assign _T_10048 = _T_10043[4]; // @[Bitwise.scala 50:65:@10105.4]
  assign _T_10049 = _T_10043[5]; // @[Bitwise.scala 50:65:@10106.4]
  assign _T_10050 = _T_10043[6]; // @[Bitwise.scala 50:65:@10107.4]
  assign _T_10051 = _T_10043[7]; // @[Bitwise.scala 50:65:@10108.4]
  assign _T_10052 = _T_10043[8]; // @[Bitwise.scala 50:65:@10109.4]
  assign _T_10053 = _T_10043[9]; // @[Bitwise.scala 50:65:@10110.4]
  assign _T_10054 = _T_10043[10]; // @[Bitwise.scala 50:65:@10111.4]
  assign _T_10055 = _T_10043[11]; // @[Bitwise.scala 50:65:@10112.4]
  assign _T_10056 = _T_10043[12]; // @[Bitwise.scala 50:65:@10113.4]
  assign _T_10057 = _T_10043[13]; // @[Bitwise.scala 50:65:@10114.4]
  assign _T_10058 = _T_10043[14]; // @[Bitwise.scala 50:65:@10115.4]
  assign _T_10059 = _T_10043[15]; // @[Bitwise.scala 50:65:@10116.4]
  assign _T_10060 = _T_10043[16]; // @[Bitwise.scala 50:65:@10117.4]
  assign _T_10061 = _T_10043[17]; // @[Bitwise.scala 50:65:@10118.4]
  assign _T_10062 = _T_10043[18]; // @[Bitwise.scala 50:65:@10119.4]
  assign _T_10063 = _T_10043[19]; // @[Bitwise.scala 50:65:@10120.4]
  assign _T_10064 = _T_10043[20]; // @[Bitwise.scala 50:65:@10121.4]
  assign _T_10065 = _T_10043[21]; // @[Bitwise.scala 50:65:@10122.4]
  assign _T_10066 = _T_10043[22]; // @[Bitwise.scala 50:65:@10123.4]
  assign _T_10067 = _T_10043[23]; // @[Bitwise.scala 50:65:@10124.4]
  assign _T_10068 = _T_10043[24]; // @[Bitwise.scala 50:65:@10125.4]
  assign _T_10069 = _T_10043[25]; // @[Bitwise.scala 50:65:@10126.4]
  assign _T_10070 = _T_10043[26]; // @[Bitwise.scala 50:65:@10127.4]
  assign _T_10071 = _T_10043[27]; // @[Bitwise.scala 50:65:@10128.4]
  assign _T_10072 = _T_10043[28]; // @[Bitwise.scala 50:65:@10129.4]
  assign _T_10073 = _T_10043[29]; // @[Bitwise.scala 50:65:@10130.4]
  assign _T_10074 = _T_10043[30]; // @[Bitwise.scala 50:65:@10131.4]
  assign _T_10075 = _T_10043[31]; // @[Bitwise.scala 50:65:@10132.4]
  assign _T_10076 = _T_10043[32]; // @[Bitwise.scala 50:65:@10133.4]
  assign _T_10077 = _T_10043[33]; // @[Bitwise.scala 50:65:@10134.4]
  assign _T_10078 = _T_10043[34]; // @[Bitwise.scala 50:65:@10135.4]
  assign _T_10079 = _T_10043[35]; // @[Bitwise.scala 50:65:@10136.4]
  assign _T_10080 = _T_10043[36]; // @[Bitwise.scala 50:65:@10137.4]
  assign _T_10081 = _T_10043[37]; // @[Bitwise.scala 50:65:@10138.4]
  assign _T_10082 = _T_10043[38]; // @[Bitwise.scala 50:65:@10139.4]
  assign _T_10083 = _T_10043[39]; // @[Bitwise.scala 50:65:@10140.4]
  assign _T_10084 = _T_10043[40]; // @[Bitwise.scala 50:65:@10141.4]
  assign _T_10085 = _T_10043[41]; // @[Bitwise.scala 50:65:@10142.4]
  assign _T_10086 = _T_10043[42]; // @[Bitwise.scala 50:65:@10143.4]
  assign _T_10087 = _T_10043[43]; // @[Bitwise.scala 50:65:@10144.4]
  assign _T_10088 = _T_10043[44]; // @[Bitwise.scala 50:65:@10145.4]
  assign _T_10089 = _T_10043[45]; // @[Bitwise.scala 50:65:@10146.4]
  assign _T_10090 = _T_10043[46]; // @[Bitwise.scala 50:65:@10147.4]
  assign _T_10091 = _T_10043[47]; // @[Bitwise.scala 50:65:@10148.4]
  assign _T_10092 = _T_10043[48]; // @[Bitwise.scala 50:65:@10149.4]
  assign _T_10093 = _T_10043[49]; // @[Bitwise.scala 50:65:@10150.4]
  assign _T_10094 = _T_10043[50]; // @[Bitwise.scala 50:65:@10151.4]
  assign _T_10095 = _T_10043[51]; // @[Bitwise.scala 50:65:@10152.4]
  assign _T_10096 = _T_10043[52]; // @[Bitwise.scala 50:65:@10153.4]
  assign _T_10097 = _T_10043[53]; // @[Bitwise.scala 50:65:@10154.4]
  assign _T_10098 = _T_10043[54]; // @[Bitwise.scala 50:65:@10155.4]
  assign _T_10099 = _T_10043[55]; // @[Bitwise.scala 50:65:@10156.4]
  assign _T_10100 = _T_10043[56]; // @[Bitwise.scala 50:65:@10157.4]
  assign _T_10101 = _T_10043[57]; // @[Bitwise.scala 50:65:@10158.4]
  assign _T_10102 = _T_10043[58]; // @[Bitwise.scala 50:65:@10159.4]
  assign _T_10103 = _T_10043[59]; // @[Bitwise.scala 50:65:@10160.4]
  assign _T_10104 = _T_10043[60]; // @[Bitwise.scala 50:65:@10161.4]
  assign _T_10105 = _T_10043[61]; // @[Bitwise.scala 50:65:@10162.4]
  assign _T_10106 = _T_10043[62]; // @[Bitwise.scala 50:65:@10163.4]
  assign _T_10107 = _T_10045 + _T_10046; // @[Bitwise.scala 48:55:@10164.4]
  assign _GEN_996 = {{1'd0}, _T_10044}; // @[Bitwise.scala 48:55:@10165.4]
  assign _T_10108 = _GEN_996 + _T_10107; // @[Bitwise.scala 48:55:@10165.4]
  assign _T_10109 = _T_10047 + _T_10048; // @[Bitwise.scala 48:55:@10166.4]
  assign _T_10110 = _T_10049 + _T_10050; // @[Bitwise.scala 48:55:@10167.4]
  assign _T_10111 = _T_10109 + _T_10110; // @[Bitwise.scala 48:55:@10168.4]
  assign _T_10112 = _T_10108 + _T_10111; // @[Bitwise.scala 48:55:@10169.4]
  assign _T_10113 = _T_10051 + _T_10052; // @[Bitwise.scala 48:55:@10170.4]
  assign _T_10114 = _T_10053 + _T_10054; // @[Bitwise.scala 48:55:@10171.4]
  assign _T_10115 = _T_10113 + _T_10114; // @[Bitwise.scala 48:55:@10172.4]
  assign _T_10116 = _T_10055 + _T_10056; // @[Bitwise.scala 48:55:@10173.4]
  assign _T_10117 = _T_10057 + _T_10058; // @[Bitwise.scala 48:55:@10174.4]
  assign _T_10118 = _T_10116 + _T_10117; // @[Bitwise.scala 48:55:@10175.4]
  assign _T_10119 = _T_10115 + _T_10118; // @[Bitwise.scala 48:55:@10176.4]
  assign _T_10120 = _T_10112 + _T_10119; // @[Bitwise.scala 48:55:@10177.4]
  assign _T_10121 = _T_10059 + _T_10060; // @[Bitwise.scala 48:55:@10178.4]
  assign _T_10122 = _T_10061 + _T_10062; // @[Bitwise.scala 48:55:@10179.4]
  assign _T_10123 = _T_10121 + _T_10122; // @[Bitwise.scala 48:55:@10180.4]
  assign _T_10124 = _T_10063 + _T_10064; // @[Bitwise.scala 48:55:@10181.4]
  assign _T_10125 = _T_10065 + _T_10066; // @[Bitwise.scala 48:55:@10182.4]
  assign _T_10126 = _T_10124 + _T_10125; // @[Bitwise.scala 48:55:@10183.4]
  assign _T_10127 = _T_10123 + _T_10126; // @[Bitwise.scala 48:55:@10184.4]
  assign _T_10128 = _T_10067 + _T_10068; // @[Bitwise.scala 48:55:@10185.4]
  assign _T_10129 = _T_10069 + _T_10070; // @[Bitwise.scala 48:55:@10186.4]
  assign _T_10130 = _T_10128 + _T_10129; // @[Bitwise.scala 48:55:@10187.4]
  assign _T_10131 = _T_10071 + _T_10072; // @[Bitwise.scala 48:55:@10188.4]
  assign _T_10132 = _T_10073 + _T_10074; // @[Bitwise.scala 48:55:@10189.4]
  assign _T_10133 = _T_10131 + _T_10132; // @[Bitwise.scala 48:55:@10190.4]
  assign _T_10134 = _T_10130 + _T_10133; // @[Bitwise.scala 48:55:@10191.4]
  assign _T_10135 = _T_10127 + _T_10134; // @[Bitwise.scala 48:55:@10192.4]
  assign _T_10136 = _T_10120 + _T_10135; // @[Bitwise.scala 48:55:@10193.4]
  assign _T_10137 = _T_10075 + _T_10076; // @[Bitwise.scala 48:55:@10194.4]
  assign _T_10138 = _T_10077 + _T_10078; // @[Bitwise.scala 48:55:@10195.4]
  assign _T_10139 = _T_10137 + _T_10138; // @[Bitwise.scala 48:55:@10196.4]
  assign _T_10140 = _T_10079 + _T_10080; // @[Bitwise.scala 48:55:@10197.4]
  assign _T_10141 = _T_10081 + _T_10082; // @[Bitwise.scala 48:55:@10198.4]
  assign _T_10142 = _T_10140 + _T_10141; // @[Bitwise.scala 48:55:@10199.4]
  assign _T_10143 = _T_10139 + _T_10142; // @[Bitwise.scala 48:55:@10200.4]
  assign _T_10144 = _T_10083 + _T_10084; // @[Bitwise.scala 48:55:@10201.4]
  assign _T_10145 = _T_10085 + _T_10086; // @[Bitwise.scala 48:55:@10202.4]
  assign _T_10146 = _T_10144 + _T_10145; // @[Bitwise.scala 48:55:@10203.4]
  assign _T_10147 = _T_10087 + _T_10088; // @[Bitwise.scala 48:55:@10204.4]
  assign _T_10148 = _T_10089 + _T_10090; // @[Bitwise.scala 48:55:@10205.4]
  assign _T_10149 = _T_10147 + _T_10148; // @[Bitwise.scala 48:55:@10206.4]
  assign _T_10150 = _T_10146 + _T_10149; // @[Bitwise.scala 48:55:@10207.4]
  assign _T_10151 = _T_10143 + _T_10150; // @[Bitwise.scala 48:55:@10208.4]
  assign _T_10152 = _T_10091 + _T_10092; // @[Bitwise.scala 48:55:@10209.4]
  assign _T_10153 = _T_10093 + _T_10094; // @[Bitwise.scala 48:55:@10210.4]
  assign _T_10154 = _T_10152 + _T_10153; // @[Bitwise.scala 48:55:@10211.4]
  assign _T_10155 = _T_10095 + _T_10096; // @[Bitwise.scala 48:55:@10212.4]
  assign _T_10156 = _T_10097 + _T_10098; // @[Bitwise.scala 48:55:@10213.4]
  assign _T_10157 = _T_10155 + _T_10156; // @[Bitwise.scala 48:55:@10214.4]
  assign _T_10158 = _T_10154 + _T_10157; // @[Bitwise.scala 48:55:@10215.4]
  assign _T_10159 = _T_10099 + _T_10100; // @[Bitwise.scala 48:55:@10216.4]
  assign _T_10160 = _T_10101 + _T_10102; // @[Bitwise.scala 48:55:@10217.4]
  assign _T_10161 = _T_10159 + _T_10160; // @[Bitwise.scala 48:55:@10218.4]
  assign _T_10162 = _T_10103 + _T_10104; // @[Bitwise.scala 48:55:@10219.4]
  assign _T_10163 = _T_10105 + _T_10106; // @[Bitwise.scala 48:55:@10220.4]
  assign _T_10164 = _T_10162 + _T_10163; // @[Bitwise.scala 48:55:@10221.4]
  assign _T_10165 = _T_10161 + _T_10164; // @[Bitwise.scala 48:55:@10222.4]
  assign _T_10166 = _T_10158 + _T_10165; // @[Bitwise.scala 48:55:@10223.4]
  assign _T_10167 = _T_10151 + _T_10166; // @[Bitwise.scala 48:55:@10224.4]
  assign _T_10168 = _T_10136 + _T_10167; // @[Bitwise.scala 48:55:@10225.4]
  assign _T_10234 = _T_2230[1]; // @[Bitwise.scala 50:65:@10292.4]
  assign _T_10235 = _T_2230[2]; // @[Bitwise.scala 50:65:@10293.4]
  assign _T_10236 = _T_2230[3]; // @[Bitwise.scala 50:65:@10294.4]
  assign _T_10237 = _T_2230[4]; // @[Bitwise.scala 50:65:@10295.4]
  assign _T_10238 = _T_2230[5]; // @[Bitwise.scala 50:65:@10296.4]
  assign _T_10239 = _T_2230[6]; // @[Bitwise.scala 50:65:@10297.4]
  assign _T_10240 = _T_2230[7]; // @[Bitwise.scala 50:65:@10298.4]
  assign _T_10241 = _T_2230[8]; // @[Bitwise.scala 50:65:@10299.4]
  assign _T_10242 = _T_2230[9]; // @[Bitwise.scala 50:65:@10300.4]
  assign _T_10243 = _T_2230[10]; // @[Bitwise.scala 50:65:@10301.4]
  assign _T_10244 = _T_2230[11]; // @[Bitwise.scala 50:65:@10302.4]
  assign _T_10245 = _T_2230[12]; // @[Bitwise.scala 50:65:@10303.4]
  assign _T_10246 = _T_2230[13]; // @[Bitwise.scala 50:65:@10304.4]
  assign _T_10247 = _T_2230[14]; // @[Bitwise.scala 50:65:@10305.4]
  assign _T_10248 = _T_2230[15]; // @[Bitwise.scala 50:65:@10306.4]
  assign _T_10249 = _T_2230[16]; // @[Bitwise.scala 50:65:@10307.4]
  assign _T_10250 = _T_2230[17]; // @[Bitwise.scala 50:65:@10308.4]
  assign _T_10251 = _T_2230[18]; // @[Bitwise.scala 50:65:@10309.4]
  assign _T_10252 = _T_2230[19]; // @[Bitwise.scala 50:65:@10310.4]
  assign _T_10253 = _T_2230[20]; // @[Bitwise.scala 50:65:@10311.4]
  assign _T_10254 = _T_2230[21]; // @[Bitwise.scala 50:65:@10312.4]
  assign _T_10255 = _T_2230[22]; // @[Bitwise.scala 50:65:@10313.4]
  assign _T_10256 = _T_2230[23]; // @[Bitwise.scala 50:65:@10314.4]
  assign _T_10257 = _T_2230[24]; // @[Bitwise.scala 50:65:@10315.4]
  assign _T_10258 = _T_2230[25]; // @[Bitwise.scala 50:65:@10316.4]
  assign _T_10259 = _T_2230[26]; // @[Bitwise.scala 50:65:@10317.4]
  assign _T_10260 = _T_2230[27]; // @[Bitwise.scala 50:65:@10318.4]
  assign _T_10261 = _T_2230[28]; // @[Bitwise.scala 50:65:@10319.4]
  assign _T_10262 = _T_2230[29]; // @[Bitwise.scala 50:65:@10320.4]
  assign _T_10263 = _T_2230[30]; // @[Bitwise.scala 50:65:@10321.4]
  assign _T_10264 = _T_2230[31]; // @[Bitwise.scala 50:65:@10322.4]
  assign _T_10265 = _T_2230[32]; // @[Bitwise.scala 50:65:@10323.4]
  assign _T_10266 = _T_2230[33]; // @[Bitwise.scala 50:65:@10324.4]
  assign _T_10267 = _T_2230[34]; // @[Bitwise.scala 50:65:@10325.4]
  assign _T_10268 = _T_2230[35]; // @[Bitwise.scala 50:65:@10326.4]
  assign _T_10269 = _T_2230[36]; // @[Bitwise.scala 50:65:@10327.4]
  assign _T_10270 = _T_2230[37]; // @[Bitwise.scala 50:65:@10328.4]
  assign _T_10271 = _T_2230[38]; // @[Bitwise.scala 50:65:@10329.4]
  assign _T_10272 = _T_2230[39]; // @[Bitwise.scala 50:65:@10330.4]
  assign _T_10273 = _T_2230[40]; // @[Bitwise.scala 50:65:@10331.4]
  assign _T_10274 = _T_2230[41]; // @[Bitwise.scala 50:65:@10332.4]
  assign _T_10275 = _T_2230[42]; // @[Bitwise.scala 50:65:@10333.4]
  assign _T_10276 = _T_2230[43]; // @[Bitwise.scala 50:65:@10334.4]
  assign _T_10277 = _T_2230[44]; // @[Bitwise.scala 50:65:@10335.4]
  assign _T_10278 = _T_2230[45]; // @[Bitwise.scala 50:65:@10336.4]
  assign _T_10279 = _T_2230[46]; // @[Bitwise.scala 50:65:@10337.4]
  assign _T_10280 = _T_2230[47]; // @[Bitwise.scala 50:65:@10338.4]
  assign _T_10281 = _T_2230[48]; // @[Bitwise.scala 50:65:@10339.4]
  assign _T_10282 = _T_2230[49]; // @[Bitwise.scala 50:65:@10340.4]
  assign _T_10283 = _T_2230[50]; // @[Bitwise.scala 50:65:@10341.4]
  assign _T_10284 = _T_2230[51]; // @[Bitwise.scala 50:65:@10342.4]
  assign _T_10285 = _T_2230[52]; // @[Bitwise.scala 50:65:@10343.4]
  assign _T_10286 = _T_2230[53]; // @[Bitwise.scala 50:65:@10344.4]
  assign _T_10287 = _T_2230[54]; // @[Bitwise.scala 50:65:@10345.4]
  assign _T_10288 = _T_2230[55]; // @[Bitwise.scala 50:65:@10346.4]
  assign _T_10289 = _T_2230[56]; // @[Bitwise.scala 50:65:@10347.4]
  assign _T_10290 = _T_2230[57]; // @[Bitwise.scala 50:65:@10348.4]
  assign _T_10291 = _T_2230[58]; // @[Bitwise.scala 50:65:@10349.4]
  assign _T_10292 = _T_2230[59]; // @[Bitwise.scala 50:65:@10350.4]
  assign _T_10293 = _T_2230[60]; // @[Bitwise.scala 50:65:@10351.4]
  assign _T_10294 = _T_2230[61]; // @[Bitwise.scala 50:65:@10352.4]
  assign _T_10295 = _T_2230[62]; // @[Bitwise.scala 50:65:@10353.4]
  assign _T_10296 = _T_2230[63]; // @[Bitwise.scala 50:65:@10354.4]
  assign _T_10297 = _T_2231 + _T_10234; // @[Bitwise.scala 48:55:@10355.4]
  assign _T_10298 = _T_10235 + _T_10236; // @[Bitwise.scala 48:55:@10356.4]
  assign _T_10299 = _T_10297 + _T_10298; // @[Bitwise.scala 48:55:@10357.4]
  assign _T_10300 = _T_10237 + _T_10238; // @[Bitwise.scala 48:55:@10358.4]
  assign _T_10301 = _T_10239 + _T_10240; // @[Bitwise.scala 48:55:@10359.4]
  assign _T_10302 = _T_10300 + _T_10301; // @[Bitwise.scala 48:55:@10360.4]
  assign _T_10303 = _T_10299 + _T_10302; // @[Bitwise.scala 48:55:@10361.4]
  assign _T_10304 = _T_10241 + _T_10242; // @[Bitwise.scala 48:55:@10362.4]
  assign _T_10305 = _T_10243 + _T_10244; // @[Bitwise.scala 48:55:@10363.4]
  assign _T_10306 = _T_10304 + _T_10305; // @[Bitwise.scala 48:55:@10364.4]
  assign _T_10307 = _T_10245 + _T_10246; // @[Bitwise.scala 48:55:@10365.4]
  assign _T_10308 = _T_10247 + _T_10248; // @[Bitwise.scala 48:55:@10366.4]
  assign _T_10309 = _T_10307 + _T_10308; // @[Bitwise.scala 48:55:@10367.4]
  assign _T_10310 = _T_10306 + _T_10309; // @[Bitwise.scala 48:55:@10368.4]
  assign _T_10311 = _T_10303 + _T_10310; // @[Bitwise.scala 48:55:@10369.4]
  assign _T_10312 = _T_10249 + _T_10250; // @[Bitwise.scala 48:55:@10370.4]
  assign _T_10313 = _T_10251 + _T_10252; // @[Bitwise.scala 48:55:@10371.4]
  assign _T_10314 = _T_10312 + _T_10313; // @[Bitwise.scala 48:55:@10372.4]
  assign _T_10315 = _T_10253 + _T_10254; // @[Bitwise.scala 48:55:@10373.4]
  assign _T_10316 = _T_10255 + _T_10256; // @[Bitwise.scala 48:55:@10374.4]
  assign _T_10317 = _T_10315 + _T_10316; // @[Bitwise.scala 48:55:@10375.4]
  assign _T_10318 = _T_10314 + _T_10317; // @[Bitwise.scala 48:55:@10376.4]
  assign _T_10319 = _T_10257 + _T_10258; // @[Bitwise.scala 48:55:@10377.4]
  assign _T_10320 = _T_10259 + _T_10260; // @[Bitwise.scala 48:55:@10378.4]
  assign _T_10321 = _T_10319 + _T_10320; // @[Bitwise.scala 48:55:@10379.4]
  assign _T_10322 = _T_10261 + _T_10262; // @[Bitwise.scala 48:55:@10380.4]
  assign _T_10323 = _T_10263 + _T_10264; // @[Bitwise.scala 48:55:@10381.4]
  assign _T_10324 = _T_10322 + _T_10323; // @[Bitwise.scala 48:55:@10382.4]
  assign _T_10325 = _T_10321 + _T_10324; // @[Bitwise.scala 48:55:@10383.4]
  assign _T_10326 = _T_10318 + _T_10325; // @[Bitwise.scala 48:55:@10384.4]
  assign _T_10327 = _T_10311 + _T_10326; // @[Bitwise.scala 48:55:@10385.4]
  assign _T_10328 = _T_10265 + _T_10266; // @[Bitwise.scala 48:55:@10386.4]
  assign _T_10329 = _T_10267 + _T_10268; // @[Bitwise.scala 48:55:@10387.4]
  assign _T_10330 = _T_10328 + _T_10329; // @[Bitwise.scala 48:55:@10388.4]
  assign _T_10331 = _T_10269 + _T_10270; // @[Bitwise.scala 48:55:@10389.4]
  assign _T_10332 = _T_10271 + _T_10272; // @[Bitwise.scala 48:55:@10390.4]
  assign _T_10333 = _T_10331 + _T_10332; // @[Bitwise.scala 48:55:@10391.4]
  assign _T_10334 = _T_10330 + _T_10333; // @[Bitwise.scala 48:55:@10392.4]
  assign _T_10335 = _T_10273 + _T_10274; // @[Bitwise.scala 48:55:@10393.4]
  assign _T_10336 = _T_10275 + _T_10276; // @[Bitwise.scala 48:55:@10394.4]
  assign _T_10337 = _T_10335 + _T_10336; // @[Bitwise.scala 48:55:@10395.4]
  assign _T_10338 = _T_10277 + _T_10278; // @[Bitwise.scala 48:55:@10396.4]
  assign _T_10339 = _T_10279 + _T_10280; // @[Bitwise.scala 48:55:@10397.4]
  assign _T_10340 = _T_10338 + _T_10339; // @[Bitwise.scala 48:55:@10398.4]
  assign _T_10341 = _T_10337 + _T_10340; // @[Bitwise.scala 48:55:@10399.4]
  assign _T_10342 = _T_10334 + _T_10341; // @[Bitwise.scala 48:55:@10400.4]
  assign _T_10343 = _T_10281 + _T_10282; // @[Bitwise.scala 48:55:@10401.4]
  assign _T_10344 = _T_10283 + _T_10284; // @[Bitwise.scala 48:55:@10402.4]
  assign _T_10345 = _T_10343 + _T_10344; // @[Bitwise.scala 48:55:@10403.4]
  assign _T_10346 = _T_10285 + _T_10286; // @[Bitwise.scala 48:55:@10404.4]
  assign _T_10347 = _T_10287 + _T_10288; // @[Bitwise.scala 48:55:@10405.4]
  assign _T_10348 = _T_10346 + _T_10347; // @[Bitwise.scala 48:55:@10406.4]
  assign _T_10349 = _T_10345 + _T_10348; // @[Bitwise.scala 48:55:@10407.4]
  assign _T_10350 = _T_10289 + _T_10290; // @[Bitwise.scala 48:55:@10408.4]
  assign _T_10351 = _T_10291 + _T_10292; // @[Bitwise.scala 48:55:@10409.4]
  assign _T_10352 = _T_10350 + _T_10351; // @[Bitwise.scala 48:55:@10410.4]
  assign _T_10353 = _T_10293 + _T_10294; // @[Bitwise.scala 48:55:@10411.4]
  assign _T_10354 = _T_10295 + _T_10296; // @[Bitwise.scala 48:55:@10412.4]
  assign _T_10355 = _T_10353 + _T_10354; // @[Bitwise.scala 48:55:@10413.4]
  assign _T_10356 = _T_10352 + _T_10355; // @[Bitwise.scala 48:55:@10414.4]
  assign _T_10357 = _T_10349 + _T_10356; // @[Bitwise.scala 48:55:@10415.4]
  assign _T_10358 = _T_10342 + _T_10357; // @[Bitwise.scala 48:55:@10416.4]
  assign _T_10359 = _T_10327 + _T_10358; // @[Bitwise.scala 48:55:@10417.4]
  assign _GEN_128 = io_input_valid ? io_input_bits_sel_0 : _T_10641_0; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_129 = io_input_valid ? io_input_bits_sel_1 : _T_10641_1; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_130 = io_input_valid ? io_input_bits_sel_2 : _T_10641_2; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_131 = io_input_valid ? io_input_bits_sel_3 : _T_10641_3; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_132 = io_input_valid ? io_input_bits_sel_4 : _T_10641_4; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_133 = io_input_valid ? io_input_bits_sel_5 : _T_10641_5; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_134 = io_input_valid ? io_input_bits_sel_6 : _T_10641_6; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_135 = io_input_valid ? io_input_bits_sel_7 : _T_10641_7; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_136 = io_input_valid ? io_input_bits_sel_8 : _T_10641_8; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_137 = io_input_valid ? io_input_bits_sel_9 : _T_10641_9; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_138 = io_input_valid ? io_input_bits_sel_10 : _T_10641_10; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_139 = io_input_valid ? io_input_bits_sel_11 : _T_10641_11; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_140 = io_input_valid ? io_input_bits_sel_12 : _T_10641_12; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_141 = io_input_valid ? io_input_bits_sel_13 : _T_10641_13; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_142 = io_input_valid ? io_input_bits_sel_14 : _T_10641_14; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_143 = io_input_valid ? io_input_bits_sel_15 : _T_10641_15; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_144 = io_input_valid ? io_input_bits_sel_16 : _T_10641_16; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_145 = io_input_valid ? io_input_bits_sel_17 : _T_10641_17; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_146 = io_input_valid ? io_input_bits_sel_18 : _T_10641_18; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_147 = io_input_valid ? io_input_bits_sel_19 : _T_10641_19; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_148 = io_input_valid ? io_input_bits_sel_20 : _T_10641_20; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_149 = io_input_valid ? io_input_bits_sel_21 : _T_10641_21; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_150 = io_input_valid ? io_input_bits_sel_22 : _T_10641_22; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_151 = io_input_valid ? io_input_bits_sel_23 : _T_10641_23; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_152 = io_input_valid ? io_input_bits_sel_24 : _T_10641_24; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_153 = io_input_valid ? io_input_bits_sel_25 : _T_10641_25; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_154 = io_input_valid ? io_input_bits_sel_26 : _T_10641_26; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_155 = io_input_valid ? io_input_bits_sel_27 : _T_10641_27; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_156 = io_input_valid ? io_input_bits_sel_28 : _T_10641_28; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_157 = io_input_valid ? io_input_bits_sel_29 : _T_10641_29; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_158 = io_input_valid ? io_input_bits_sel_30 : _T_10641_30; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _GEN_159 = io_input_valid ? io_input_bits_sel_31 : _T_10641_31; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@10586.4]
  assign _T_11318 = io_input_mask_en[0]; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@10748.4]
  assign _T_11319 = io_input_valid & _T_11318; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@10749.4]
  assign _GEN_160 = _T_11319 ? _T_2231 : _T_11317_0; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10750.4]
  assign _GEN_161 = _T_11319 ? _T_2299 : _T_11317_1; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10755.4]
  assign _T_2167_2 = _T_2368[1:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2366.4]
  assign _GEN_162 = _T_11319 ? _T_2167_2 : _T_11317_2; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10760.4]
  assign _GEN_163 = _T_11319 ? _T_2439 : _T_11317_3; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10765.4]
  assign _T_2167_4 = _T_2512[2:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2512.4]
  assign _GEN_164 = _T_11319 ? _T_2167_4 : _T_11317_4; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10770.4]
  assign _T_2167_5 = _T_2587[2:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2588.4]
  assign _GEN_165 = _T_11319 ? _T_2167_5 : _T_11317_5; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10775.4]
  assign _T_2167_6 = _T_2664[2:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2666.4]
  assign _GEN_166 = _T_11319 ? _T_2167_6 : _T_11317_6; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10780.4]
  assign _GEN_167 = _T_11319 ? _T_2743 : _T_11317_7; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10785.4]
  assign _T_11334 = io_input_mask_en[1]; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@10788.4]
  assign _T_11335 = io_input_valid & _T_11334; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@10789.4]
  assign _T_2167_8 = _T_2824[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2828.4]
  assign _GEN_168 = _T_11335 ? _T_2167_8 : _T_11317_8; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10790.4]
  assign _T_2167_9 = _T_2907[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2912.4]
  assign _GEN_169 = _T_11335 ? _T_2167_9 : _T_11317_9; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10795.4]
  assign _T_2167_10 = _T_2992[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2998.4]
  assign _GEN_170 = _T_11335 ? _T_2167_10 : _T_11317_10; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10800.4]
  assign _T_2167_11 = _T_3079[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3086.4]
  assign _GEN_171 = _T_11335 ? _T_2167_11 : _T_11317_11; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10805.4]
  assign _T_2167_12 = _T_3168[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3176.4]
  assign _GEN_172 = _T_11335 ? _T_2167_12 : _T_11317_12; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10810.4]
  assign _T_2167_13 = _T_3259[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3268.4]
  assign _GEN_173 = _T_11335 ? _T_2167_13 : _T_11317_13; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10815.4]
  assign _T_2167_14 = _T_3352[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3362.4]
  assign _GEN_174 = _T_11335 ? _T_2167_14 : _T_11317_14; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10820.4]
  assign _GEN_175 = _T_11335 ? _T_3447 : _T_11317_15; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10825.4]
  assign _T_11350 = io_input_mask_en[2]; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@10828.4]
  assign _T_11351 = io_input_valid & _T_11350; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@10829.4]
  assign _T_2167_16 = _T_3544[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3556.4]
  assign _GEN_176 = _T_11351 ? _T_2167_16 : _T_11317_16; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10830.4]
  assign _T_2167_17 = _T_3643[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3656.4]
  assign _GEN_177 = _T_11351 ? _T_2167_17 : _T_11317_17; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10835.4]
  assign _T_2167_18 = _T_3744[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3758.4]
  assign _GEN_178 = _T_11351 ? _T_2167_18 : _T_11317_18; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10840.4]
  assign _T_2167_19 = _T_3847[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3862.4]
  assign _GEN_179 = _T_11351 ? _T_2167_19 : _T_11317_19; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10845.4]
  assign _T_2167_20 = _T_3952[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3968.4]
  assign _GEN_180 = _T_11351 ? _T_2167_20 : _T_11317_20; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10850.4]
  assign _T_2167_21 = _T_4059[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4076.4]
  assign _GEN_181 = _T_11351 ? _T_2167_21 : _T_11317_21; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10855.4]
  assign _T_2167_22 = _T_4168[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4186.4]
  assign _GEN_182 = _T_11351 ? _T_2167_22 : _T_11317_22; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10860.4]
  assign _T_2167_23 = _T_4279[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4298.4]
  assign _GEN_183 = _T_11351 ? _T_2167_23 : _T_11317_23; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10865.4]
  assign _T_11366 = io_input_mask_en[3]; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@10868.4]
  assign _T_11367 = io_input_valid & _T_11366; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@10869.4]
  assign _T_2167_24 = _T_4392[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4412.4]
  assign _GEN_184 = _T_11367 ? _T_2167_24 : _T_11317_24; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10870.4]
  assign _T_2167_25 = _T_4507[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4528.4]
  assign _GEN_185 = _T_11367 ? _T_2167_25 : _T_11317_25; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10875.4]
  assign _T_2167_26 = _T_4624[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4646.4]
  assign _GEN_186 = _T_11367 ? _T_2167_26 : _T_11317_26; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10880.4]
  assign _T_2167_27 = _T_4743[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4766.4]
  assign _GEN_187 = _T_11367 ? _T_2167_27 : _T_11317_27; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10885.4]
  assign _T_2167_28 = _T_4864[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4888.4]
  assign _GEN_188 = _T_11367 ? _T_2167_28 : _T_11317_28; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10890.4]
  assign _T_2167_29 = _T_4987[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5012.4]
  assign _GEN_189 = _T_11367 ? _T_2167_29 : _T_11317_29; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10895.4]
  assign _T_2167_30 = _T_5112[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5138.4]
  assign _GEN_190 = _T_11367 ? _T_2167_30 : _T_11317_30; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10900.4]
  assign _GEN_191 = _T_11367 ? _T_5239 : _T_11317_31; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10905.4]
  assign _T_11382 = io_input_mask_en[4]; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@10908.4]
  assign _T_11383 = io_input_valid & _T_11382; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@10909.4]
  assign _T_2167_32 = _T_5368[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5396.4]
  assign _GEN_192 = _T_11383 ? _T_2167_32 : _T_11317_32; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10910.4]
  assign _T_2167_33 = _T_5499[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5528.4]
  assign _GEN_193 = _T_11383 ? _T_2167_33 : _T_11317_33; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10915.4]
  assign _T_2167_34 = _T_5632[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5662.4]
  assign _GEN_194 = _T_11383 ? _T_2167_34 : _T_11317_34; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10920.4]
  assign _T_2167_35 = _T_5767[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5798.4]
  assign _GEN_195 = _T_11383 ? _T_2167_35 : _T_11317_35; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10925.4]
  assign _T_2167_36 = _T_5904[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5936.4]
  assign _GEN_196 = _T_11383 ? _T_2167_36 : _T_11317_36; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10930.4]
  assign _T_2167_37 = _T_6043[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6076.4]
  assign _GEN_197 = _T_11383 ? _T_2167_37 : _T_11317_37; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10935.4]
  assign _T_2167_38 = _T_6184[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6218.4]
  assign _GEN_198 = _T_11383 ? _T_2167_38 : _T_11317_38; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10940.4]
  assign _T_2167_39 = _T_6327[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6362.4]
  assign _GEN_199 = _T_11383 ? _T_2167_39 : _T_11317_39; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10945.4]
  assign _T_11398 = io_input_mask_en[5]; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@10948.4]
  assign _T_11399 = io_input_valid & _T_11398; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@10949.4]
  assign _T_2167_40 = _T_6472[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6508.4]
  assign _GEN_200 = _T_11399 ? _T_2167_40 : _T_11317_40; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10950.4]
  assign _T_2167_41 = _T_6619[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6656.4]
  assign _GEN_201 = _T_11399 ? _T_2167_41 : _T_11317_41; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10955.4]
  assign _T_2167_42 = _T_6768[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6806.4]
  assign _GEN_202 = _T_11399 ? _T_2167_42 : _T_11317_42; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10960.4]
  assign _T_2167_43 = _T_6919[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6958.4]
  assign _GEN_203 = _T_11399 ? _T_2167_43 : _T_11317_43; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10965.4]
  assign _T_2167_44 = _T_7072[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7112.4]
  assign _GEN_204 = _T_11399 ? _T_2167_44 : _T_11317_44; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10970.4]
  assign _T_2167_45 = _T_7227[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7268.4]
  assign _GEN_205 = _T_11399 ? _T_2167_45 : _T_11317_45; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10975.4]
  assign _T_2167_46 = _T_7384[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7426.4]
  assign _GEN_206 = _T_11399 ? _T_2167_46 : _T_11317_46; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10980.4]
  assign _T_2167_47 = _T_7543[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7586.4]
  assign _GEN_207 = _T_11399 ? _T_2167_47 : _T_11317_47; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10985.4]
  assign _T_11414 = io_input_mask_en[6]; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@10988.4]
  assign _T_11415 = io_input_valid & _T_11414; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@10989.4]
  assign _T_2167_48 = _T_7704[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7748.4]
  assign _GEN_208 = _T_11415 ? _T_2167_48 : _T_11317_48; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10990.4]
  assign _T_2167_49 = _T_7867[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7912.4]
  assign _GEN_209 = _T_11415 ? _T_2167_49 : _T_11317_49; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@10995.4]
  assign _T_2167_50 = _T_8032[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@8078.4]
  assign _GEN_210 = _T_11415 ? _T_2167_50 : _T_11317_50; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11000.4]
  assign _T_2167_51 = _T_8199[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@8246.4]
  assign _GEN_211 = _T_11415 ? _T_2167_51 : _T_11317_51; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11005.4]
  assign _T_2167_52 = _T_8368[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@8416.4]
  assign _GEN_212 = _T_11415 ? _T_2167_52 : _T_11317_52; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11010.4]
  assign _T_2167_53 = _T_8539[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@8588.4]
  assign _GEN_213 = _T_11415 ? _T_2167_53 : _T_11317_53; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11015.4]
  assign _T_2167_54 = _T_8712[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@8762.4]
  assign _GEN_214 = _T_11415 ? _T_2167_54 : _T_11317_54; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11020.4]
  assign _T_2167_55 = _T_8887[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@8938.4]
  assign _GEN_215 = _T_11415 ? _T_2167_55 : _T_11317_55; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11025.4]
  assign _T_11430 = io_input_mask_en[7]; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@11028.4]
  assign _T_11431 = io_input_valid & _T_11430; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@11029.4]
  assign _T_2167_56 = _T_9064[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@9116.4]
  assign _GEN_216 = _T_11431 ? _T_2167_56 : _T_11317_56; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11030.4]
  assign _T_2167_57 = _T_9243[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@9296.4]
  assign _GEN_217 = _T_11431 ? _T_2167_57 : _T_11317_57; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11035.4]
  assign _T_2167_58 = _T_9424[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@9478.4]
  assign _GEN_218 = _T_11431 ? _T_2167_58 : _T_11317_58; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11040.4]
  assign _T_2167_59 = _T_9607[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@9662.4]
  assign _GEN_219 = _T_11431 ? _T_2167_59 : _T_11317_59; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11045.4]
  assign _T_2167_60 = _T_9792[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@9848.4]
  assign _GEN_220 = _T_11431 ? _T_2167_60 : _T_11317_60; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11050.4]
  assign _T_2167_61 = _T_9979[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@10036.4]
  assign _GEN_221 = _T_11431 ? _T_2167_61 : _T_11317_61; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11055.4]
  assign _T_2167_62 = _T_10168[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@2162.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@10226.4]
  assign _GEN_222 = _T_11431 ? _T_2167_62 : _T_11317_62; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11060.4]
  assign _GEN_223 = _T_11431 ? _T_10359 : _T_11317_63; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@11065.4]
  assign _T_11519 = _T_11317_0 ? _T_10366_0 : 8'h0; // @[Mux.scala 46:16:@11070.4]
  assign _T_11523 = 2'h2 == _T_11317_1; // @[Mux.scala 46:19:@11072.4]
  assign _T_11524 = _T_11523 ? _T_10366_1 : 8'h0; // @[Mux.scala 46:16:@11073.4]
  assign _T_11525 = 2'h1 == _T_11317_1; // @[Mux.scala 46:19:@11074.4]
  assign _T_11526 = _T_11525 ? _T_10366_0 : _T_11524; // @[Mux.scala 46:16:@11075.4]
  assign _T_11531 = 2'h3 == _T_11317_2; // @[Mux.scala 46:19:@11077.4]
  assign _T_11532 = _T_11531 ? _T_10366_2 : 8'h0; // @[Mux.scala 46:16:@11078.4]
  assign _T_11533 = 2'h2 == _T_11317_2; // @[Mux.scala 46:19:@11079.4]
  assign _T_11534 = _T_11533 ? _T_10366_1 : _T_11532; // @[Mux.scala 46:16:@11080.4]
  assign _T_11535 = 2'h1 == _T_11317_2; // @[Mux.scala 46:19:@11081.4]
  assign _T_11536 = _T_11535 ? _T_10366_0 : _T_11534; // @[Mux.scala 46:16:@11082.4]
  assign _T_11542 = 3'h4 == _T_11317_3; // @[Mux.scala 46:19:@11084.4]
  assign _T_11543 = _T_11542 ? _T_10366_3 : 8'h0; // @[Mux.scala 46:16:@11085.4]
  assign _T_11544 = 3'h3 == _T_11317_3; // @[Mux.scala 46:19:@11086.4]
  assign _T_11545 = _T_11544 ? _T_10366_2 : _T_11543; // @[Mux.scala 46:16:@11087.4]
  assign _T_11546 = 3'h2 == _T_11317_3; // @[Mux.scala 46:19:@11088.4]
  assign _T_11547 = _T_11546 ? _T_10366_1 : _T_11545; // @[Mux.scala 46:16:@11089.4]
  assign _T_11548 = 3'h1 == _T_11317_3; // @[Mux.scala 46:19:@11090.4]
  assign _T_11549 = _T_11548 ? _T_10366_0 : _T_11547; // @[Mux.scala 46:16:@11091.4]
  assign _T_11556 = 3'h5 == _T_11317_4; // @[Mux.scala 46:19:@11093.4]
  assign _T_11557 = _T_11556 ? _T_10366_4 : 8'h0; // @[Mux.scala 46:16:@11094.4]
  assign _T_11558 = 3'h4 == _T_11317_4; // @[Mux.scala 46:19:@11095.4]
  assign _T_11559 = _T_11558 ? _T_10366_3 : _T_11557; // @[Mux.scala 46:16:@11096.4]
  assign _T_11560 = 3'h3 == _T_11317_4; // @[Mux.scala 46:19:@11097.4]
  assign _T_11561 = _T_11560 ? _T_10366_2 : _T_11559; // @[Mux.scala 46:16:@11098.4]
  assign _T_11562 = 3'h2 == _T_11317_4; // @[Mux.scala 46:19:@11099.4]
  assign _T_11563 = _T_11562 ? _T_10366_1 : _T_11561; // @[Mux.scala 46:16:@11100.4]
  assign _T_11564 = 3'h1 == _T_11317_4; // @[Mux.scala 46:19:@11101.4]
  assign _T_11565 = _T_11564 ? _T_10366_0 : _T_11563; // @[Mux.scala 46:16:@11102.4]
  assign _T_11573 = 3'h6 == _T_11317_5; // @[Mux.scala 46:19:@11104.4]
  assign _T_11574 = _T_11573 ? _T_10366_5 : 8'h0; // @[Mux.scala 46:16:@11105.4]
  assign _T_11575 = 3'h5 == _T_11317_5; // @[Mux.scala 46:19:@11106.4]
  assign _T_11576 = _T_11575 ? _T_10366_4 : _T_11574; // @[Mux.scala 46:16:@11107.4]
  assign _T_11577 = 3'h4 == _T_11317_5; // @[Mux.scala 46:19:@11108.4]
  assign _T_11578 = _T_11577 ? _T_10366_3 : _T_11576; // @[Mux.scala 46:16:@11109.4]
  assign _T_11579 = 3'h3 == _T_11317_5; // @[Mux.scala 46:19:@11110.4]
  assign _T_11580 = _T_11579 ? _T_10366_2 : _T_11578; // @[Mux.scala 46:16:@11111.4]
  assign _T_11581 = 3'h2 == _T_11317_5; // @[Mux.scala 46:19:@11112.4]
  assign _T_11582 = _T_11581 ? _T_10366_1 : _T_11580; // @[Mux.scala 46:16:@11113.4]
  assign _T_11583 = 3'h1 == _T_11317_5; // @[Mux.scala 46:19:@11114.4]
  assign _T_11584 = _T_11583 ? _T_10366_0 : _T_11582; // @[Mux.scala 46:16:@11115.4]
  assign _T_11593 = 3'h7 == _T_11317_6; // @[Mux.scala 46:19:@11117.4]
  assign _T_11594 = _T_11593 ? _T_10366_6 : 8'h0; // @[Mux.scala 46:16:@11118.4]
  assign _T_11595 = 3'h6 == _T_11317_6; // @[Mux.scala 46:19:@11119.4]
  assign _T_11596 = _T_11595 ? _T_10366_5 : _T_11594; // @[Mux.scala 46:16:@11120.4]
  assign _T_11597 = 3'h5 == _T_11317_6; // @[Mux.scala 46:19:@11121.4]
  assign _T_11598 = _T_11597 ? _T_10366_4 : _T_11596; // @[Mux.scala 46:16:@11122.4]
  assign _T_11599 = 3'h4 == _T_11317_6; // @[Mux.scala 46:19:@11123.4]
  assign _T_11600 = _T_11599 ? _T_10366_3 : _T_11598; // @[Mux.scala 46:16:@11124.4]
  assign _T_11601 = 3'h3 == _T_11317_6; // @[Mux.scala 46:19:@11125.4]
  assign _T_11602 = _T_11601 ? _T_10366_2 : _T_11600; // @[Mux.scala 46:16:@11126.4]
  assign _T_11603 = 3'h2 == _T_11317_6; // @[Mux.scala 46:19:@11127.4]
  assign _T_11604 = _T_11603 ? _T_10366_1 : _T_11602; // @[Mux.scala 46:16:@11128.4]
  assign _T_11605 = 3'h1 == _T_11317_6; // @[Mux.scala 46:19:@11129.4]
  assign _T_11606 = _T_11605 ? _T_10366_0 : _T_11604; // @[Mux.scala 46:16:@11130.4]
  assign _T_11616 = 4'h8 == _T_11317_7; // @[Mux.scala 46:19:@11132.4]
  assign _T_11617 = _T_11616 ? _T_10366_7 : 8'h0; // @[Mux.scala 46:16:@11133.4]
  assign _T_11618 = 4'h7 == _T_11317_7; // @[Mux.scala 46:19:@11134.4]
  assign _T_11619 = _T_11618 ? _T_10366_6 : _T_11617; // @[Mux.scala 46:16:@11135.4]
  assign _T_11620 = 4'h6 == _T_11317_7; // @[Mux.scala 46:19:@11136.4]
  assign _T_11621 = _T_11620 ? _T_10366_5 : _T_11619; // @[Mux.scala 46:16:@11137.4]
  assign _T_11622 = 4'h5 == _T_11317_7; // @[Mux.scala 46:19:@11138.4]
  assign _T_11623 = _T_11622 ? _T_10366_4 : _T_11621; // @[Mux.scala 46:16:@11139.4]
  assign _T_11624 = 4'h4 == _T_11317_7; // @[Mux.scala 46:19:@11140.4]
  assign _T_11625 = _T_11624 ? _T_10366_3 : _T_11623; // @[Mux.scala 46:16:@11141.4]
  assign _T_11626 = 4'h3 == _T_11317_7; // @[Mux.scala 46:19:@11142.4]
  assign _T_11627 = _T_11626 ? _T_10366_2 : _T_11625; // @[Mux.scala 46:16:@11143.4]
  assign _T_11628 = 4'h2 == _T_11317_7; // @[Mux.scala 46:19:@11144.4]
  assign _T_11629 = _T_11628 ? _T_10366_1 : _T_11627; // @[Mux.scala 46:16:@11145.4]
  assign _T_11630 = 4'h1 == _T_11317_7; // @[Mux.scala 46:19:@11146.4]
  assign _T_11631 = _T_11630 ? _T_10366_0 : _T_11629; // @[Mux.scala 46:16:@11147.4]
  assign _T_11642 = 4'h9 == _T_11317_8; // @[Mux.scala 46:19:@11149.4]
  assign _T_11643 = _T_11642 ? _T_10366_8 : 8'h0; // @[Mux.scala 46:16:@11150.4]
  assign _T_11644 = 4'h8 == _T_11317_8; // @[Mux.scala 46:19:@11151.4]
  assign _T_11645 = _T_11644 ? _T_10366_7 : _T_11643; // @[Mux.scala 46:16:@11152.4]
  assign _T_11646 = 4'h7 == _T_11317_8; // @[Mux.scala 46:19:@11153.4]
  assign _T_11647 = _T_11646 ? _T_10366_6 : _T_11645; // @[Mux.scala 46:16:@11154.4]
  assign _T_11648 = 4'h6 == _T_11317_8; // @[Mux.scala 46:19:@11155.4]
  assign _T_11649 = _T_11648 ? _T_10366_5 : _T_11647; // @[Mux.scala 46:16:@11156.4]
  assign _T_11650 = 4'h5 == _T_11317_8; // @[Mux.scala 46:19:@11157.4]
  assign _T_11651 = _T_11650 ? _T_10366_4 : _T_11649; // @[Mux.scala 46:16:@11158.4]
  assign _T_11652 = 4'h4 == _T_11317_8; // @[Mux.scala 46:19:@11159.4]
  assign _T_11653 = _T_11652 ? _T_10366_3 : _T_11651; // @[Mux.scala 46:16:@11160.4]
  assign _T_11654 = 4'h3 == _T_11317_8; // @[Mux.scala 46:19:@11161.4]
  assign _T_11655 = _T_11654 ? _T_10366_2 : _T_11653; // @[Mux.scala 46:16:@11162.4]
  assign _T_11656 = 4'h2 == _T_11317_8; // @[Mux.scala 46:19:@11163.4]
  assign _T_11657 = _T_11656 ? _T_10366_1 : _T_11655; // @[Mux.scala 46:16:@11164.4]
  assign _T_11658 = 4'h1 == _T_11317_8; // @[Mux.scala 46:19:@11165.4]
  assign _T_11659 = _T_11658 ? _T_10366_0 : _T_11657; // @[Mux.scala 46:16:@11166.4]
  assign _T_11671 = 4'ha == _T_11317_9; // @[Mux.scala 46:19:@11168.4]
  assign _T_11672 = _T_11671 ? _T_10366_9 : 8'h0; // @[Mux.scala 46:16:@11169.4]
  assign _T_11673 = 4'h9 == _T_11317_9; // @[Mux.scala 46:19:@11170.4]
  assign _T_11674 = _T_11673 ? _T_10366_8 : _T_11672; // @[Mux.scala 46:16:@11171.4]
  assign _T_11675 = 4'h8 == _T_11317_9; // @[Mux.scala 46:19:@11172.4]
  assign _T_11676 = _T_11675 ? _T_10366_7 : _T_11674; // @[Mux.scala 46:16:@11173.4]
  assign _T_11677 = 4'h7 == _T_11317_9; // @[Mux.scala 46:19:@11174.4]
  assign _T_11678 = _T_11677 ? _T_10366_6 : _T_11676; // @[Mux.scala 46:16:@11175.4]
  assign _T_11679 = 4'h6 == _T_11317_9; // @[Mux.scala 46:19:@11176.4]
  assign _T_11680 = _T_11679 ? _T_10366_5 : _T_11678; // @[Mux.scala 46:16:@11177.4]
  assign _T_11681 = 4'h5 == _T_11317_9; // @[Mux.scala 46:19:@11178.4]
  assign _T_11682 = _T_11681 ? _T_10366_4 : _T_11680; // @[Mux.scala 46:16:@11179.4]
  assign _T_11683 = 4'h4 == _T_11317_9; // @[Mux.scala 46:19:@11180.4]
  assign _T_11684 = _T_11683 ? _T_10366_3 : _T_11682; // @[Mux.scala 46:16:@11181.4]
  assign _T_11685 = 4'h3 == _T_11317_9; // @[Mux.scala 46:19:@11182.4]
  assign _T_11686 = _T_11685 ? _T_10366_2 : _T_11684; // @[Mux.scala 46:16:@11183.4]
  assign _T_11687 = 4'h2 == _T_11317_9; // @[Mux.scala 46:19:@11184.4]
  assign _T_11688 = _T_11687 ? _T_10366_1 : _T_11686; // @[Mux.scala 46:16:@11185.4]
  assign _T_11689 = 4'h1 == _T_11317_9; // @[Mux.scala 46:19:@11186.4]
  assign _T_11690 = _T_11689 ? _T_10366_0 : _T_11688; // @[Mux.scala 46:16:@11187.4]
  assign _T_11703 = 4'hb == _T_11317_10; // @[Mux.scala 46:19:@11189.4]
  assign _T_11704 = _T_11703 ? _T_10366_10 : 8'h0; // @[Mux.scala 46:16:@11190.4]
  assign _T_11705 = 4'ha == _T_11317_10; // @[Mux.scala 46:19:@11191.4]
  assign _T_11706 = _T_11705 ? _T_10366_9 : _T_11704; // @[Mux.scala 46:16:@11192.4]
  assign _T_11707 = 4'h9 == _T_11317_10; // @[Mux.scala 46:19:@11193.4]
  assign _T_11708 = _T_11707 ? _T_10366_8 : _T_11706; // @[Mux.scala 46:16:@11194.4]
  assign _T_11709 = 4'h8 == _T_11317_10; // @[Mux.scala 46:19:@11195.4]
  assign _T_11710 = _T_11709 ? _T_10366_7 : _T_11708; // @[Mux.scala 46:16:@11196.4]
  assign _T_11711 = 4'h7 == _T_11317_10; // @[Mux.scala 46:19:@11197.4]
  assign _T_11712 = _T_11711 ? _T_10366_6 : _T_11710; // @[Mux.scala 46:16:@11198.4]
  assign _T_11713 = 4'h6 == _T_11317_10; // @[Mux.scala 46:19:@11199.4]
  assign _T_11714 = _T_11713 ? _T_10366_5 : _T_11712; // @[Mux.scala 46:16:@11200.4]
  assign _T_11715 = 4'h5 == _T_11317_10; // @[Mux.scala 46:19:@11201.4]
  assign _T_11716 = _T_11715 ? _T_10366_4 : _T_11714; // @[Mux.scala 46:16:@11202.4]
  assign _T_11717 = 4'h4 == _T_11317_10; // @[Mux.scala 46:19:@11203.4]
  assign _T_11718 = _T_11717 ? _T_10366_3 : _T_11716; // @[Mux.scala 46:16:@11204.4]
  assign _T_11719 = 4'h3 == _T_11317_10; // @[Mux.scala 46:19:@11205.4]
  assign _T_11720 = _T_11719 ? _T_10366_2 : _T_11718; // @[Mux.scala 46:16:@11206.4]
  assign _T_11721 = 4'h2 == _T_11317_10; // @[Mux.scala 46:19:@11207.4]
  assign _T_11722 = _T_11721 ? _T_10366_1 : _T_11720; // @[Mux.scala 46:16:@11208.4]
  assign _T_11723 = 4'h1 == _T_11317_10; // @[Mux.scala 46:19:@11209.4]
  assign _T_11724 = _T_11723 ? _T_10366_0 : _T_11722; // @[Mux.scala 46:16:@11210.4]
  assign _T_11738 = 4'hc == _T_11317_11; // @[Mux.scala 46:19:@11212.4]
  assign _T_11739 = _T_11738 ? _T_10366_11 : 8'h0; // @[Mux.scala 46:16:@11213.4]
  assign _T_11740 = 4'hb == _T_11317_11; // @[Mux.scala 46:19:@11214.4]
  assign _T_11741 = _T_11740 ? _T_10366_10 : _T_11739; // @[Mux.scala 46:16:@11215.4]
  assign _T_11742 = 4'ha == _T_11317_11; // @[Mux.scala 46:19:@11216.4]
  assign _T_11743 = _T_11742 ? _T_10366_9 : _T_11741; // @[Mux.scala 46:16:@11217.4]
  assign _T_11744 = 4'h9 == _T_11317_11; // @[Mux.scala 46:19:@11218.4]
  assign _T_11745 = _T_11744 ? _T_10366_8 : _T_11743; // @[Mux.scala 46:16:@11219.4]
  assign _T_11746 = 4'h8 == _T_11317_11; // @[Mux.scala 46:19:@11220.4]
  assign _T_11747 = _T_11746 ? _T_10366_7 : _T_11745; // @[Mux.scala 46:16:@11221.4]
  assign _T_11748 = 4'h7 == _T_11317_11; // @[Mux.scala 46:19:@11222.4]
  assign _T_11749 = _T_11748 ? _T_10366_6 : _T_11747; // @[Mux.scala 46:16:@11223.4]
  assign _T_11750 = 4'h6 == _T_11317_11; // @[Mux.scala 46:19:@11224.4]
  assign _T_11751 = _T_11750 ? _T_10366_5 : _T_11749; // @[Mux.scala 46:16:@11225.4]
  assign _T_11752 = 4'h5 == _T_11317_11; // @[Mux.scala 46:19:@11226.4]
  assign _T_11753 = _T_11752 ? _T_10366_4 : _T_11751; // @[Mux.scala 46:16:@11227.4]
  assign _T_11754 = 4'h4 == _T_11317_11; // @[Mux.scala 46:19:@11228.4]
  assign _T_11755 = _T_11754 ? _T_10366_3 : _T_11753; // @[Mux.scala 46:16:@11229.4]
  assign _T_11756 = 4'h3 == _T_11317_11; // @[Mux.scala 46:19:@11230.4]
  assign _T_11757 = _T_11756 ? _T_10366_2 : _T_11755; // @[Mux.scala 46:16:@11231.4]
  assign _T_11758 = 4'h2 == _T_11317_11; // @[Mux.scala 46:19:@11232.4]
  assign _T_11759 = _T_11758 ? _T_10366_1 : _T_11757; // @[Mux.scala 46:16:@11233.4]
  assign _T_11760 = 4'h1 == _T_11317_11; // @[Mux.scala 46:19:@11234.4]
  assign _T_11761 = _T_11760 ? _T_10366_0 : _T_11759; // @[Mux.scala 46:16:@11235.4]
  assign _T_11776 = 4'hd == _T_11317_12; // @[Mux.scala 46:19:@11237.4]
  assign _T_11777 = _T_11776 ? _T_10366_12 : 8'h0; // @[Mux.scala 46:16:@11238.4]
  assign _T_11778 = 4'hc == _T_11317_12; // @[Mux.scala 46:19:@11239.4]
  assign _T_11779 = _T_11778 ? _T_10366_11 : _T_11777; // @[Mux.scala 46:16:@11240.4]
  assign _T_11780 = 4'hb == _T_11317_12; // @[Mux.scala 46:19:@11241.4]
  assign _T_11781 = _T_11780 ? _T_10366_10 : _T_11779; // @[Mux.scala 46:16:@11242.4]
  assign _T_11782 = 4'ha == _T_11317_12; // @[Mux.scala 46:19:@11243.4]
  assign _T_11783 = _T_11782 ? _T_10366_9 : _T_11781; // @[Mux.scala 46:16:@11244.4]
  assign _T_11784 = 4'h9 == _T_11317_12; // @[Mux.scala 46:19:@11245.4]
  assign _T_11785 = _T_11784 ? _T_10366_8 : _T_11783; // @[Mux.scala 46:16:@11246.4]
  assign _T_11786 = 4'h8 == _T_11317_12; // @[Mux.scala 46:19:@11247.4]
  assign _T_11787 = _T_11786 ? _T_10366_7 : _T_11785; // @[Mux.scala 46:16:@11248.4]
  assign _T_11788 = 4'h7 == _T_11317_12; // @[Mux.scala 46:19:@11249.4]
  assign _T_11789 = _T_11788 ? _T_10366_6 : _T_11787; // @[Mux.scala 46:16:@11250.4]
  assign _T_11790 = 4'h6 == _T_11317_12; // @[Mux.scala 46:19:@11251.4]
  assign _T_11791 = _T_11790 ? _T_10366_5 : _T_11789; // @[Mux.scala 46:16:@11252.4]
  assign _T_11792 = 4'h5 == _T_11317_12; // @[Mux.scala 46:19:@11253.4]
  assign _T_11793 = _T_11792 ? _T_10366_4 : _T_11791; // @[Mux.scala 46:16:@11254.4]
  assign _T_11794 = 4'h4 == _T_11317_12; // @[Mux.scala 46:19:@11255.4]
  assign _T_11795 = _T_11794 ? _T_10366_3 : _T_11793; // @[Mux.scala 46:16:@11256.4]
  assign _T_11796 = 4'h3 == _T_11317_12; // @[Mux.scala 46:19:@11257.4]
  assign _T_11797 = _T_11796 ? _T_10366_2 : _T_11795; // @[Mux.scala 46:16:@11258.4]
  assign _T_11798 = 4'h2 == _T_11317_12; // @[Mux.scala 46:19:@11259.4]
  assign _T_11799 = _T_11798 ? _T_10366_1 : _T_11797; // @[Mux.scala 46:16:@11260.4]
  assign _T_11800 = 4'h1 == _T_11317_12; // @[Mux.scala 46:19:@11261.4]
  assign _T_11801 = _T_11800 ? _T_10366_0 : _T_11799; // @[Mux.scala 46:16:@11262.4]
  assign _T_11817 = 4'he == _T_11317_13; // @[Mux.scala 46:19:@11264.4]
  assign _T_11818 = _T_11817 ? _T_10366_13 : 8'h0; // @[Mux.scala 46:16:@11265.4]
  assign _T_11819 = 4'hd == _T_11317_13; // @[Mux.scala 46:19:@11266.4]
  assign _T_11820 = _T_11819 ? _T_10366_12 : _T_11818; // @[Mux.scala 46:16:@11267.4]
  assign _T_11821 = 4'hc == _T_11317_13; // @[Mux.scala 46:19:@11268.4]
  assign _T_11822 = _T_11821 ? _T_10366_11 : _T_11820; // @[Mux.scala 46:16:@11269.4]
  assign _T_11823 = 4'hb == _T_11317_13; // @[Mux.scala 46:19:@11270.4]
  assign _T_11824 = _T_11823 ? _T_10366_10 : _T_11822; // @[Mux.scala 46:16:@11271.4]
  assign _T_11825 = 4'ha == _T_11317_13; // @[Mux.scala 46:19:@11272.4]
  assign _T_11826 = _T_11825 ? _T_10366_9 : _T_11824; // @[Mux.scala 46:16:@11273.4]
  assign _T_11827 = 4'h9 == _T_11317_13; // @[Mux.scala 46:19:@11274.4]
  assign _T_11828 = _T_11827 ? _T_10366_8 : _T_11826; // @[Mux.scala 46:16:@11275.4]
  assign _T_11829 = 4'h8 == _T_11317_13; // @[Mux.scala 46:19:@11276.4]
  assign _T_11830 = _T_11829 ? _T_10366_7 : _T_11828; // @[Mux.scala 46:16:@11277.4]
  assign _T_11831 = 4'h7 == _T_11317_13; // @[Mux.scala 46:19:@11278.4]
  assign _T_11832 = _T_11831 ? _T_10366_6 : _T_11830; // @[Mux.scala 46:16:@11279.4]
  assign _T_11833 = 4'h6 == _T_11317_13; // @[Mux.scala 46:19:@11280.4]
  assign _T_11834 = _T_11833 ? _T_10366_5 : _T_11832; // @[Mux.scala 46:16:@11281.4]
  assign _T_11835 = 4'h5 == _T_11317_13; // @[Mux.scala 46:19:@11282.4]
  assign _T_11836 = _T_11835 ? _T_10366_4 : _T_11834; // @[Mux.scala 46:16:@11283.4]
  assign _T_11837 = 4'h4 == _T_11317_13; // @[Mux.scala 46:19:@11284.4]
  assign _T_11838 = _T_11837 ? _T_10366_3 : _T_11836; // @[Mux.scala 46:16:@11285.4]
  assign _T_11839 = 4'h3 == _T_11317_13; // @[Mux.scala 46:19:@11286.4]
  assign _T_11840 = _T_11839 ? _T_10366_2 : _T_11838; // @[Mux.scala 46:16:@11287.4]
  assign _T_11841 = 4'h2 == _T_11317_13; // @[Mux.scala 46:19:@11288.4]
  assign _T_11842 = _T_11841 ? _T_10366_1 : _T_11840; // @[Mux.scala 46:16:@11289.4]
  assign _T_11843 = 4'h1 == _T_11317_13; // @[Mux.scala 46:19:@11290.4]
  assign _T_11844 = _T_11843 ? _T_10366_0 : _T_11842; // @[Mux.scala 46:16:@11291.4]
  assign _T_11861 = 4'hf == _T_11317_14; // @[Mux.scala 46:19:@11293.4]
  assign _T_11862 = _T_11861 ? _T_10366_14 : 8'h0; // @[Mux.scala 46:16:@11294.4]
  assign _T_11863 = 4'he == _T_11317_14; // @[Mux.scala 46:19:@11295.4]
  assign _T_11864 = _T_11863 ? _T_10366_13 : _T_11862; // @[Mux.scala 46:16:@11296.4]
  assign _T_11865 = 4'hd == _T_11317_14; // @[Mux.scala 46:19:@11297.4]
  assign _T_11866 = _T_11865 ? _T_10366_12 : _T_11864; // @[Mux.scala 46:16:@11298.4]
  assign _T_11867 = 4'hc == _T_11317_14; // @[Mux.scala 46:19:@11299.4]
  assign _T_11868 = _T_11867 ? _T_10366_11 : _T_11866; // @[Mux.scala 46:16:@11300.4]
  assign _T_11869 = 4'hb == _T_11317_14; // @[Mux.scala 46:19:@11301.4]
  assign _T_11870 = _T_11869 ? _T_10366_10 : _T_11868; // @[Mux.scala 46:16:@11302.4]
  assign _T_11871 = 4'ha == _T_11317_14; // @[Mux.scala 46:19:@11303.4]
  assign _T_11872 = _T_11871 ? _T_10366_9 : _T_11870; // @[Mux.scala 46:16:@11304.4]
  assign _T_11873 = 4'h9 == _T_11317_14; // @[Mux.scala 46:19:@11305.4]
  assign _T_11874 = _T_11873 ? _T_10366_8 : _T_11872; // @[Mux.scala 46:16:@11306.4]
  assign _T_11875 = 4'h8 == _T_11317_14; // @[Mux.scala 46:19:@11307.4]
  assign _T_11876 = _T_11875 ? _T_10366_7 : _T_11874; // @[Mux.scala 46:16:@11308.4]
  assign _T_11877 = 4'h7 == _T_11317_14; // @[Mux.scala 46:19:@11309.4]
  assign _T_11878 = _T_11877 ? _T_10366_6 : _T_11876; // @[Mux.scala 46:16:@11310.4]
  assign _T_11879 = 4'h6 == _T_11317_14; // @[Mux.scala 46:19:@11311.4]
  assign _T_11880 = _T_11879 ? _T_10366_5 : _T_11878; // @[Mux.scala 46:16:@11312.4]
  assign _T_11881 = 4'h5 == _T_11317_14; // @[Mux.scala 46:19:@11313.4]
  assign _T_11882 = _T_11881 ? _T_10366_4 : _T_11880; // @[Mux.scala 46:16:@11314.4]
  assign _T_11883 = 4'h4 == _T_11317_14; // @[Mux.scala 46:19:@11315.4]
  assign _T_11884 = _T_11883 ? _T_10366_3 : _T_11882; // @[Mux.scala 46:16:@11316.4]
  assign _T_11885 = 4'h3 == _T_11317_14; // @[Mux.scala 46:19:@11317.4]
  assign _T_11886 = _T_11885 ? _T_10366_2 : _T_11884; // @[Mux.scala 46:16:@11318.4]
  assign _T_11887 = 4'h2 == _T_11317_14; // @[Mux.scala 46:19:@11319.4]
  assign _T_11888 = _T_11887 ? _T_10366_1 : _T_11886; // @[Mux.scala 46:16:@11320.4]
  assign _T_11889 = 4'h1 == _T_11317_14; // @[Mux.scala 46:19:@11321.4]
  assign _T_11890 = _T_11889 ? _T_10366_0 : _T_11888; // @[Mux.scala 46:16:@11322.4]
  assign _T_11908 = 5'h10 == _T_11317_15; // @[Mux.scala 46:19:@11324.4]
  assign _T_11909 = _T_11908 ? _T_10366_15 : 8'h0; // @[Mux.scala 46:16:@11325.4]
  assign _T_11910 = 5'hf == _T_11317_15; // @[Mux.scala 46:19:@11326.4]
  assign _T_11911 = _T_11910 ? _T_10366_14 : _T_11909; // @[Mux.scala 46:16:@11327.4]
  assign _T_11912 = 5'he == _T_11317_15; // @[Mux.scala 46:19:@11328.4]
  assign _T_11913 = _T_11912 ? _T_10366_13 : _T_11911; // @[Mux.scala 46:16:@11329.4]
  assign _T_11914 = 5'hd == _T_11317_15; // @[Mux.scala 46:19:@11330.4]
  assign _T_11915 = _T_11914 ? _T_10366_12 : _T_11913; // @[Mux.scala 46:16:@11331.4]
  assign _T_11916 = 5'hc == _T_11317_15; // @[Mux.scala 46:19:@11332.4]
  assign _T_11917 = _T_11916 ? _T_10366_11 : _T_11915; // @[Mux.scala 46:16:@11333.4]
  assign _T_11918 = 5'hb == _T_11317_15; // @[Mux.scala 46:19:@11334.4]
  assign _T_11919 = _T_11918 ? _T_10366_10 : _T_11917; // @[Mux.scala 46:16:@11335.4]
  assign _T_11920 = 5'ha == _T_11317_15; // @[Mux.scala 46:19:@11336.4]
  assign _T_11921 = _T_11920 ? _T_10366_9 : _T_11919; // @[Mux.scala 46:16:@11337.4]
  assign _T_11922 = 5'h9 == _T_11317_15; // @[Mux.scala 46:19:@11338.4]
  assign _T_11923 = _T_11922 ? _T_10366_8 : _T_11921; // @[Mux.scala 46:16:@11339.4]
  assign _T_11924 = 5'h8 == _T_11317_15; // @[Mux.scala 46:19:@11340.4]
  assign _T_11925 = _T_11924 ? _T_10366_7 : _T_11923; // @[Mux.scala 46:16:@11341.4]
  assign _T_11926 = 5'h7 == _T_11317_15; // @[Mux.scala 46:19:@11342.4]
  assign _T_11927 = _T_11926 ? _T_10366_6 : _T_11925; // @[Mux.scala 46:16:@11343.4]
  assign _T_11928 = 5'h6 == _T_11317_15; // @[Mux.scala 46:19:@11344.4]
  assign _T_11929 = _T_11928 ? _T_10366_5 : _T_11927; // @[Mux.scala 46:16:@11345.4]
  assign _T_11930 = 5'h5 == _T_11317_15; // @[Mux.scala 46:19:@11346.4]
  assign _T_11931 = _T_11930 ? _T_10366_4 : _T_11929; // @[Mux.scala 46:16:@11347.4]
  assign _T_11932 = 5'h4 == _T_11317_15; // @[Mux.scala 46:19:@11348.4]
  assign _T_11933 = _T_11932 ? _T_10366_3 : _T_11931; // @[Mux.scala 46:16:@11349.4]
  assign _T_11934 = 5'h3 == _T_11317_15; // @[Mux.scala 46:19:@11350.4]
  assign _T_11935 = _T_11934 ? _T_10366_2 : _T_11933; // @[Mux.scala 46:16:@11351.4]
  assign _T_11936 = 5'h2 == _T_11317_15; // @[Mux.scala 46:19:@11352.4]
  assign _T_11937 = _T_11936 ? _T_10366_1 : _T_11935; // @[Mux.scala 46:16:@11353.4]
  assign _T_11938 = 5'h1 == _T_11317_15; // @[Mux.scala 46:19:@11354.4]
  assign _T_11939 = _T_11938 ? _T_10366_0 : _T_11937; // @[Mux.scala 46:16:@11355.4]
  assign _T_11958 = 5'h11 == _T_11317_16; // @[Mux.scala 46:19:@11357.4]
  assign _T_11959 = _T_11958 ? _T_10366_16 : 8'h0; // @[Mux.scala 46:16:@11358.4]
  assign _T_11960 = 5'h10 == _T_11317_16; // @[Mux.scala 46:19:@11359.4]
  assign _T_11961 = _T_11960 ? _T_10366_15 : _T_11959; // @[Mux.scala 46:16:@11360.4]
  assign _T_11962 = 5'hf == _T_11317_16; // @[Mux.scala 46:19:@11361.4]
  assign _T_11963 = _T_11962 ? _T_10366_14 : _T_11961; // @[Mux.scala 46:16:@11362.4]
  assign _T_11964 = 5'he == _T_11317_16; // @[Mux.scala 46:19:@11363.4]
  assign _T_11965 = _T_11964 ? _T_10366_13 : _T_11963; // @[Mux.scala 46:16:@11364.4]
  assign _T_11966 = 5'hd == _T_11317_16; // @[Mux.scala 46:19:@11365.4]
  assign _T_11967 = _T_11966 ? _T_10366_12 : _T_11965; // @[Mux.scala 46:16:@11366.4]
  assign _T_11968 = 5'hc == _T_11317_16; // @[Mux.scala 46:19:@11367.4]
  assign _T_11969 = _T_11968 ? _T_10366_11 : _T_11967; // @[Mux.scala 46:16:@11368.4]
  assign _T_11970 = 5'hb == _T_11317_16; // @[Mux.scala 46:19:@11369.4]
  assign _T_11971 = _T_11970 ? _T_10366_10 : _T_11969; // @[Mux.scala 46:16:@11370.4]
  assign _T_11972 = 5'ha == _T_11317_16; // @[Mux.scala 46:19:@11371.4]
  assign _T_11973 = _T_11972 ? _T_10366_9 : _T_11971; // @[Mux.scala 46:16:@11372.4]
  assign _T_11974 = 5'h9 == _T_11317_16; // @[Mux.scala 46:19:@11373.4]
  assign _T_11975 = _T_11974 ? _T_10366_8 : _T_11973; // @[Mux.scala 46:16:@11374.4]
  assign _T_11976 = 5'h8 == _T_11317_16; // @[Mux.scala 46:19:@11375.4]
  assign _T_11977 = _T_11976 ? _T_10366_7 : _T_11975; // @[Mux.scala 46:16:@11376.4]
  assign _T_11978 = 5'h7 == _T_11317_16; // @[Mux.scala 46:19:@11377.4]
  assign _T_11979 = _T_11978 ? _T_10366_6 : _T_11977; // @[Mux.scala 46:16:@11378.4]
  assign _T_11980 = 5'h6 == _T_11317_16; // @[Mux.scala 46:19:@11379.4]
  assign _T_11981 = _T_11980 ? _T_10366_5 : _T_11979; // @[Mux.scala 46:16:@11380.4]
  assign _T_11982 = 5'h5 == _T_11317_16; // @[Mux.scala 46:19:@11381.4]
  assign _T_11983 = _T_11982 ? _T_10366_4 : _T_11981; // @[Mux.scala 46:16:@11382.4]
  assign _T_11984 = 5'h4 == _T_11317_16; // @[Mux.scala 46:19:@11383.4]
  assign _T_11985 = _T_11984 ? _T_10366_3 : _T_11983; // @[Mux.scala 46:16:@11384.4]
  assign _T_11986 = 5'h3 == _T_11317_16; // @[Mux.scala 46:19:@11385.4]
  assign _T_11987 = _T_11986 ? _T_10366_2 : _T_11985; // @[Mux.scala 46:16:@11386.4]
  assign _T_11988 = 5'h2 == _T_11317_16; // @[Mux.scala 46:19:@11387.4]
  assign _T_11989 = _T_11988 ? _T_10366_1 : _T_11987; // @[Mux.scala 46:16:@11388.4]
  assign _T_11990 = 5'h1 == _T_11317_16; // @[Mux.scala 46:19:@11389.4]
  assign _T_11991 = _T_11990 ? _T_10366_0 : _T_11989; // @[Mux.scala 46:16:@11390.4]
  assign _T_12011 = 5'h12 == _T_11317_17; // @[Mux.scala 46:19:@11392.4]
  assign _T_12012 = _T_12011 ? _T_10366_17 : 8'h0; // @[Mux.scala 46:16:@11393.4]
  assign _T_12013 = 5'h11 == _T_11317_17; // @[Mux.scala 46:19:@11394.4]
  assign _T_12014 = _T_12013 ? _T_10366_16 : _T_12012; // @[Mux.scala 46:16:@11395.4]
  assign _T_12015 = 5'h10 == _T_11317_17; // @[Mux.scala 46:19:@11396.4]
  assign _T_12016 = _T_12015 ? _T_10366_15 : _T_12014; // @[Mux.scala 46:16:@11397.4]
  assign _T_12017 = 5'hf == _T_11317_17; // @[Mux.scala 46:19:@11398.4]
  assign _T_12018 = _T_12017 ? _T_10366_14 : _T_12016; // @[Mux.scala 46:16:@11399.4]
  assign _T_12019 = 5'he == _T_11317_17; // @[Mux.scala 46:19:@11400.4]
  assign _T_12020 = _T_12019 ? _T_10366_13 : _T_12018; // @[Mux.scala 46:16:@11401.4]
  assign _T_12021 = 5'hd == _T_11317_17; // @[Mux.scala 46:19:@11402.4]
  assign _T_12022 = _T_12021 ? _T_10366_12 : _T_12020; // @[Mux.scala 46:16:@11403.4]
  assign _T_12023 = 5'hc == _T_11317_17; // @[Mux.scala 46:19:@11404.4]
  assign _T_12024 = _T_12023 ? _T_10366_11 : _T_12022; // @[Mux.scala 46:16:@11405.4]
  assign _T_12025 = 5'hb == _T_11317_17; // @[Mux.scala 46:19:@11406.4]
  assign _T_12026 = _T_12025 ? _T_10366_10 : _T_12024; // @[Mux.scala 46:16:@11407.4]
  assign _T_12027 = 5'ha == _T_11317_17; // @[Mux.scala 46:19:@11408.4]
  assign _T_12028 = _T_12027 ? _T_10366_9 : _T_12026; // @[Mux.scala 46:16:@11409.4]
  assign _T_12029 = 5'h9 == _T_11317_17; // @[Mux.scala 46:19:@11410.4]
  assign _T_12030 = _T_12029 ? _T_10366_8 : _T_12028; // @[Mux.scala 46:16:@11411.4]
  assign _T_12031 = 5'h8 == _T_11317_17; // @[Mux.scala 46:19:@11412.4]
  assign _T_12032 = _T_12031 ? _T_10366_7 : _T_12030; // @[Mux.scala 46:16:@11413.4]
  assign _T_12033 = 5'h7 == _T_11317_17; // @[Mux.scala 46:19:@11414.4]
  assign _T_12034 = _T_12033 ? _T_10366_6 : _T_12032; // @[Mux.scala 46:16:@11415.4]
  assign _T_12035 = 5'h6 == _T_11317_17; // @[Mux.scala 46:19:@11416.4]
  assign _T_12036 = _T_12035 ? _T_10366_5 : _T_12034; // @[Mux.scala 46:16:@11417.4]
  assign _T_12037 = 5'h5 == _T_11317_17; // @[Mux.scala 46:19:@11418.4]
  assign _T_12038 = _T_12037 ? _T_10366_4 : _T_12036; // @[Mux.scala 46:16:@11419.4]
  assign _T_12039 = 5'h4 == _T_11317_17; // @[Mux.scala 46:19:@11420.4]
  assign _T_12040 = _T_12039 ? _T_10366_3 : _T_12038; // @[Mux.scala 46:16:@11421.4]
  assign _T_12041 = 5'h3 == _T_11317_17; // @[Mux.scala 46:19:@11422.4]
  assign _T_12042 = _T_12041 ? _T_10366_2 : _T_12040; // @[Mux.scala 46:16:@11423.4]
  assign _T_12043 = 5'h2 == _T_11317_17; // @[Mux.scala 46:19:@11424.4]
  assign _T_12044 = _T_12043 ? _T_10366_1 : _T_12042; // @[Mux.scala 46:16:@11425.4]
  assign _T_12045 = 5'h1 == _T_11317_17; // @[Mux.scala 46:19:@11426.4]
  assign _T_12046 = _T_12045 ? _T_10366_0 : _T_12044; // @[Mux.scala 46:16:@11427.4]
  assign _T_12067 = 5'h13 == _T_11317_18; // @[Mux.scala 46:19:@11429.4]
  assign _T_12068 = _T_12067 ? _T_10366_18 : 8'h0; // @[Mux.scala 46:16:@11430.4]
  assign _T_12069 = 5'h12 == _T_11317_18; // @[Mux.scala 46:19:@11431.4]
  assign _T_12070 = _T_12069 ? _T_10366_17 : _T_12068; // @[Mux.scala 46:16:@11432.4]
  assign _T_12071 = 5'h11 == _T_11317_18; // @[Mux.scala 46:19:@11433.4]
  assign _T_12072 = _T_12071 ? _T_10366_16 : _T_12070; // @[Mux.scala 46:16:@11434.4]
  assign _T_12073 = 5'h10 == _T_11317_18; // @[Mux.scala 46:19:@11435.4]
  assign _T_12074 = _T_12073 ? _T_10366_15 : _T_12072; // @[Mux.scala 46:16:@11436.4]
  assign _T_12075 = 5'hf == _T_11317_18; // @[Mux.scala 46:19:@11437.4]
  assign _T_12076 = _T_12075 ? _T_10366_14 : _T_12074; // @[Mux.scala 46:16:@11438.4]
  assign _T_12077 = 5'he == _T_11317_18; // @[Mux.scala 46:19:@11439.4]
  assign _T_12078 = _T_12077 ? _T_10366_13 : _T_12076; // @[Mux.scala 46:16:@11440.4]
  assign _T_12079 = 5'hd == _T_11317_18; // @[Mux.scala 46:19:@11441.4]
  assign _T_12080 = _T_12079 ? _T_10366_12 : _T_12078; // @[Mux.scala 46:16:@11442.4]
  assign _T_12081 = 5'hc == _T_11317_18; // @[Mux.scala 46:19:@11443.4]
  assign _T_12082 = _T_12081 ? _T_10366_11 : _T_12080; // @[Mux.scala 46:16:@11444.4]
  assign _T_12083 = 5'hb == _T_11317_18; // @[Mux.scala 46:19:@11445.4]
  assign _T_12084 = _T_12083 ? _T_10366_10 : _T_12082; // @[Mux.scala 46:16:@11446.4]
  assign _T_12085 = 5'ha == _T_11317_18; // @[Mux.scala 46:19:@11447.4]
  assign _T_12086 = _T_12085 ? _T_10366_9 : _T_12084; // @[Mux.scala 46:16:@11448.4]
  assign _T_12087 = 5'h9 == _T_11317_18; // @[Mux.scala 46:19:@11449.4]
  assign _T_12088 = _T_12087 ? _T_10366_8 : _T_12086; // @[Mux.scala 46:16:@11450.4]
  assign _T_12089 = 5'h8 == _T_11317_18; // @[Mux.scala 46:19:@11451.4]
  assign _T_12090 = _T_12089 ? _T_10366_7 : _T_12088; // @[Mux.scala 46:16:@11452.4]
  assign _T_12091 = 5'h7 == _T_11317_18; // @[Mux.scala 46:19:@11453.4]
  assign _T_12092 = _T_12091 ? _T_10366_6 : _T_12090; // @[Mux.scala 46:16:@11454.4]
  assign _T_12093 = 5'h6 == _T_11317_18; // @[Mux.scala 46:19:@11455.4]
  assign _T_12094 = _T_12093 ? _T_10366_5 : _T_12092; // @[Mux.scala 46:16:@11456.4]
  assign _T_12095 = 5'h5 == _T_11317_18; // @[Mux.scala 46:19:@11457.4]
  assign _T_12096 = _T_12095 ? _T_10366_4 : _T_12094; // @[Mux.scala 46:16:@11458.4]
  assign _T_12097 = 5'h4 == _T_11317_18; // @[Mux.scala 46:19:@11459.4]
  assign _T_12098 = _T_12097 ? _T_10366_3 : _T_12096; // @[Mux.scala 46:16:@11460.4]
  assign _T_12099 = 5'h3 == _T_11317_18; // @[Mux.scala 46:19:@11461.4]
  assign _T_12100 = _T_12099 ? _T_10366_2 : _T_12098; // @[Mux.scala 46:16:@11462.4]
  assign _T_12101 = 5'h2 == _T_11317_18; // @[Mux.scala 46:19:@11463.4]
  assign _T_12102 = _T_12101 ? _T_10366_1 : _T_12100; // @[Mux.scala 46:16:@11464.4]
  assign _T_12103 = 5'h1 == _T_11317_18; // @[Mux.scala 46:19:@11465.4]
  assign _T_12104 = _T_12103 ? _T_10366_0 : _T_12102; // @[Mux.scala 46:16:@11466.4]
  assign _T_12126 = 5'h14 == _T_11317_19; // @[Mux.scala 46:19:@11468.4]
  assign _T_12127 = _T_12126 ? _T_10366_19 : 8'h0; // @[Mux.scala 46:16:@11469.4]
  assign _T_12128 = 5'h13 == _T_11317_19; // @[Mux.scala 46:19:@11470.4]
  assign _T_12129 = _T_12128 ? _T_10366_18 : _T_12127; // @[Mux.scala 46:16:@11471.4]
  assign _T_12130 = 5'h12 == _T_11317_19; // @[Mux.scala 46:19:@11472.4]
  assign _T_12131 = _T_12130 ? _T_10366_17 : _T_12129; // @[Mux.scala 46:16:@11473.4]
  assign _T_12132 = 5'h11 == _T_11317_19; // @[Mux.scala 46:19:@11474.4]
  assign _T_12133 = _T_12132 ? _T_10366_16 : _T_12131; // @[Mux.scala 46:16:@11475.4]
  assign _T_12134 = 5'h10 == _T_11317_19; // @[Mux.scala 46:19:@11476.4]
  assign _T_12135 = _T_12134 ? _T_10366_15 : _T_12133; // @[Mux.scala 46:16:@11477.4]
  assign _T_12136 = 5'hf == _T_11317_19; // @[Mux.scala 46:19:@11478.4]
  assign _T_12137 = _T_12136 ? _T_10366_14 : _T_12135; // @[Mux.scala 46:16:@11479.4]
  assign _T_12138 = 5'he == _T_11317_19; // @[Mux.scala 46:19:@11480.4]
  assign _T_12139 = _T_12138 ? _T_10366_13 : _T_12137; // @[Mux.scala 46:16:@11481.4]
  assign _T_12140 = 5'hd == _T_11317_19; // @[Mux.scala 46:19:@11482.4]
  assign _T_12141 = _T_12140 ? _T_10366_12 : _T_12139; // @[Mux.scala 46:16:@11483.4]
  assign _T_12142 = 5'hc == _T_11317_19; // @[Mux.scala 46:19:@11484.4]
  assign _T_12143 = _T_12142 ? _T_10366_11 : _T_12141; // @[Mux.scala 46:16:@11485.4]
  assign _T_12144 = 5'hb == _T_11317_19; // @[Mux.scala 46:19:@11486.4]
  assign _T_12145 = _T_12144 ? _T_10366_10 : _T_12143; // @[Mux.scala 46:16:@11487.4]
  assign _T_12146 = 5'ha == _T_11317_19; // @[Mux.scala 46:19:@11488.4]
  assign _T_12147 = _T_12146 ? _T_10366_9 : _T_12145; // @[Mux.scala 46:16:@11489.4]
  assign _T_12148 = 5'h9 == _T_11317_19; // @[Mux.scala 46:19:@11490.4]
  assign _T_12149 = _T_12148 ? _T_10366_8 : _T_12147; // @[Mux.scala 46:16:@11491.4]
  assign _T_12150 = 5'h8 == _T_11317_19; // @[Mux.scala 46:19:@11492.4]
  assign _T_12151 = _T_12150 ? _T_10366_7 : _T_12149; // @[Mux.scala 46:16:@11493.4]
  assign _T_12152 = 5'h7 == _T_11317_19; // @[Mux.scala 46:19:@11494.4]
  assign _T_12153 = _T_12152 ? _T_10366_6 : _T_12151; // @[Mux.scala 46:16:@11495.4]
  assign _T_12154 = 5'h6 == _T_11317_19; // @[Mux.scala 46:19:@11496.4]
  assign _T_12155 = _T_12154 ? _T_10366_5 : _T_12153; // @[Mux.scala 46:16:@11497.4]
  assign _T_12156 = 5'h5 == _T_11317_19; // @[Mux.scala 46:19:@11498.4]
  assign _T_12157 = _T_12156 ? _T_10366_4 : _T_12155; // @[Mux.scala 46:16:@11499.4]
  assign _T_12158 = 5'h4 == _T_11317_19; // @[Mux.scala 46:19:@11500.4]
  assign _T_12159 = _T_12158 ? _T_10366_3 : _T_12157; // @[Mux.scala 46:16:@11501.4]
  assign _T_12160 = 5'h3 == _T_11317_19; // @[Mux.scala 46:19:@11502.4]
  assign _T_12161 = _T_12160 ? _T_10366_2 : _T_12159; // @[Mux.scala 46:16:@11503.4]
  assign _T_12162 = 5'h2 == _T_11317_19; // @[Mux.scala 46:19:@11504.4]
  assign _T_12163 = _T_12162 ? _T_10366_1 : _T_12161; // @[Mux.scala 46:16:@11505.4]
  assign _T_12164 = 5'h1 == _T_11317_19; // @[Mux.scala 46:19:@11506.4]
  assign _T_12165 = _T_12164 ? _T_10366_0 : _T_12163; // @[Mux.scala 46:16:@11507.4]
  assign _T_12188 = 5'h15 == _T_11317_20; // @[Mux.scala 46:19:@11509.4]
  assign _T_12189 = _T_12188 ? _T_10366_20 : 8'h0; // @[Mux.scala 46:16:@11510.4]
  assign _T_12190 = 5'h14 == _T_11317_20; // @[Mux.scala 46:19:@11511.4]
  assign _T_12191 = _T_12190 ? _T_10366_19 : _T_12189; // @[Mux.scala 46:16:@11512.4]
  assign _T_12192 = 5'h13 == _T_11317_20; // @[Mux.scala 46:19:@11513.4]
  assign _T_12193 = _T_12192 ? _T_10366_18 : _T_12191; // @[Mux.scala 46:16:@11514.4]
  assign _T_12194 = 5'h12 == _T_11317_20; // @[Mux.scala 46:19:@11515.4]
  assign _T_12195 = _T_12194 ? _T_10366_17 : _T_12193; // @[Mux.scala 46:16:@11516.4]
  assign _T_12196 = 5'h11 == _T_11317_20; // @[Mux.scala 46:19:@11517.4]
  assign _T_12197 = _T_12196 ? _T_10366_16 : _T_12195; // @[Mux.scala 46:16:@11518.4]
  assign _T_12198 = 5'h10 == _T_11317_20; // @[Mux.scala 46:19:@11519.4]
  assign _T_12199 = _T_12198 ? _T_10366_15 : _T_12197; // @[Mux.scala 46:16:@11520.4]
  assign _T_12200 = 5'hf == _T_11317_20; // @[Mux.scala 46:19:@11521.4]
  assign _T_12201 = _T_12200 ? _T_10366_14 : _T_12199; // @[Mux.scala 46:16:@11522.4]
  assign _T_12202 = 5'he == _T_11317_20; // @[Mux.scala 46:19:@11523.4]
  assign _T_12203 = _T_12202 ? _T_10366_13 : _T_12201; // @[Mux.scala 46:16:@11524.4]
  assign _T_12204 = 5'hd == _T_11317_20; // @[Mux.scala 46:19:@11525.4]
  assign _T_12205 = _T_12204 ? _T_10366_12 : _T_12203; // @[Mux.scala 46:16:@11526.4]
  assign _T_12206 = 5'hc == _T_11317_20; // @[Mux.scala 46:19:@11527.4]
  assign _T_12207 = _T_12206 ? _T_10366_11 : _T_12205; // @[Mux.scala 46:16:@11528.4]
  assign _T_12208 = 5'hb == _T_11317_20; // @[Mux.scala 46:19:@11529.4]
  assign _T_12209 = _T_12208 ? _T_10366_10 : _T_12207; // @[Mux.scala 46:16:@11530.4]
  assign _T_12210 = 5'ha == _T_11317_20; // @[Mux.scala 46:19:@11531.4]
  assign _T_12211 = _T_12210 ? _T_10366_9 : _T_12209; // @[Mux.scala 46:16:@11532.4]
  assign _T_12212 = 5'h9 == _T_11317_20; // @[Mux.scala 46:19:@11533.4]
  assign _T_12213 = _T_12212 ? _T_10366_8 : _T_12211; // @[Mux.scala 46:16:@11534.4]
  assign _T_12214 = 5'h8 == _T_11317_20; // @[Mux.scala 46:19:@11535.4]
  assign _T_12215 = _T_12214 ? _T_10366_7 : _T_12213; // @[Mux.scala 46:16:@11536.4]
  assign _T_12216 = 5'h7 == _T_11317_20; // @[Mux.scala 46:19:@11537.4]
  assign _T_12217 = _T_12216 ? _T_10366_6 : _T_12215; // @[Mux.scala 46:16:@11538.4]
  assign _T_12218 = 5'h6 == _T_11317_20; // @[Mux.scala 46:19:@11539.4]
  assign _T_12219 = _T_12218 ? _T_10366_5 : _T_12217; // @[Mux.scala 46:16:@11540.4]
  assign _T_12220 = 5'h5 == _T_11317_20; // @[Mux.scala 46:19:@11541.4]
  assign _T_12221 = _T_12220 ? _T_10366_4 : _T_12219; // @[Mux.scala 46:16:@11542.4]
  assign _T_12222 = 5'h4 == _T_11317_20; // @[Mux.scala 46:19:@11543.4]
  assign _T_12223 = _T_12222 ? _T_10366_3 : _T_12221; // @[Mux.scala 46:16:@11544.4]
  assign _T_12224 = 5'h3 == _T_11317_20; // @[Mux.scala 46:19:@11545.4]
  assign _T_12225 = _T_12224 ? _T_10366_2 : _T_12223; // @[Mux.scala 46:16:@11546.4]
  assign _T_12226 = 5'h2 == _T_11317_20; // @[Mux.scala 46:19:@11547.4]
  assign _T_12227 = _T_12226 ? _T_10366_1 : _T_12225; // @[Mux.scala 46:16:@11548.4]
  assign _T_12228 = 5'h1 == _T_11317_20; // @[Mux.scala 46:19:@11549.4]
  assign _T_12229 = _T_12228 ? _T_10366_0 : _T_12227; // @[Mux.scala 46:16:@11550.4]
  assign _T_12253 = 5'h16 == _T_11317_21; // @[Mux.scala 46:19:@11552.4]
  assign _T_12254 = _T_12253 ? _T_10366_21 : 8'h0; // @[Mux.scala 46:16:@11553.4]
  assign _T_12255 = 5'h15 == _T_11317_21; // @[Mux.scala 46:19:@11554.4]
  assign _T_12256 = _T_12255 ? _T_10366_20 : _T_12254; // @[Mux.scala 46:16:@11555.4]
  assign _T_12257 = 5'h14 == _T_11317_21; // @[Mux.scala 46:19:@11556.4]
  assign _T_12258 = _T_12257 ? _T_10366_19 : _T_12256; // @[Mux.scala 46:16:@11557.4]
  assign _T_12259 = 5'h13 == _T_11317_21; // @[Mux.scala 46:19:@11558.4]
  assign _T_12260 = _T_12259 ? _T_10366_18 : _T_12258; // @[Mux.scala 46:16:@11559.4]
  assign _T_12261 = 5'h12 == _T_11317_21; // @[Mux.scala 46:19:@11560.4]
  assign _T_12262 = _T_12261 ? _T_10366_17 : _T_12260; // @[Mux.scala 46:16:@11561.4]
  assign _T_12263 = 5'h11 == _T_11317_21; // @[Mux.scala 46:19:@11562.4]
  assign _T_12264 = _T_12263 ? _T_10366_16 : _T_12262; // @[Mux.scala 46:16:@11563.4]
  assign _T_12265 = 5'h10 == _T_11317_21; // @[Mux.scala 46:19:@11564.4]
  assign _T_12266 = _T_12265 ? _T_10366_15 : _T_12264; // @[Mux.scala 46:16:@11565.4]
  assign _T_12267 = 5'hf == _T_11317_21; // @[Mux.scala 46:19:@11566.4]
  assign _T_12268 = _T_12267 ? _T_10366_14 : _T_12266; // @[Mux.scala 46:16:@11567.4]
  assign _T_12269 = 5'he == _T_11317_21; // @[Mux.scala 46:19:@11568.4]
  assign _T_12270 = _T_12269 ? _T_10366_13 : _T_12268; // @[Mux.scala 46:16:@11569.4]
  assign _T_12271 = 5'hd == _T_11317_21; // @[Mux.scala 46:19:@11570.4]
  assign _T_12272 = _T_12271 ? _T_10366_12 : _T_12270; // @[Mux.scala 46:16:@11571.4]
  assign _T_12273 = 5'hc == _T_11317_21; // @[Mux.scala 46:19:@11572.4]
  assign _T_12274 = _T_12273 ? _T_10366_11 : _T_12272; // @[Mux.scala 46:16:@11573.4]
  assign _T_12275 = 5'hb == _T_11317_21; // @[Mux.scala 46:19:@11574.4]
  assign _T_12276 = _T_12275 ? _T_10366_10 : _T_12274; // @[Mux.scala 46:16:@11575.4]
  assign _T_12277 = 5'ha == _T_11317_21; // @[Mux.scala 46:19:@11576.4]
  assign _T_12278 = _T_12277 ? _T_10366_9 : _T_12276; // @[Mux.scala 46:16:@11577.4]
  assign _T_12279 = 5'h9 == _T_11317_21; // @[Mux.scala 46:19:@11578.4]
  assign _T_12280 = _T_12279 ? _T_10366_8 : _T_12278; // @[Mux.scala 46:16:@11579.4]
  assign _T_12281 = 5'h8 == _T_11317_21; // @[Mux.scala 46:19:@11580.4]
  assign _T_12282 = _T_12281 ? _T_10366_7 : _T_12280; // @[Mux.scala 46:16:@11581.4]
  assign _T_12283 = 5'h7 == _T_11317_21; // @[Mux.scala 46:19:@11582.4]
  assign _T_12284 = _T_12283 ? _T_10366_6 : _T_12282; // @[Mux.scala 46:16:@11583.4]
  assign _T_12285 = 5'h6 == _T_11317_21; // @[Mux.scala 46:19:@11584.4]
  assign _T_12286 = _T_12285 ? _T_10366_5 : _T_12284; // @[Mux.scala 46:16:@11585.4]
  assign _T_12287 = 5'h5 == _T_11317_21; // @[Mux.scala 46:19:@11586.4]
  assign _T_12288 = _T_12287 ? _T_10366_4 : _T_12286; // @[Mux.scala 46:16:@11587.4]
  assign _T_12289 = 5'h4 == _T_11317_21; // @[Mux.scala 46:19:@11588.4]
  assign _T_12290 = _T_12289 ? _T_10366_3 : _T_12288; // @[Mux.scala 46:16:@11589.4]
  assign _T_12291 = 5'h3 == _T_11317_21; // @[Mux.scala 46:19:@11590.4]
  assign _T_12292 = _T_12291 ? _T_10366_2 : _T_12290; // @[Mux.scala 46:16:@11591.4]
  assign _T_12293 = 5'h2 == _T_11317_21; // @[Mux.scala 46:19:@11592.4]
  assign _T_12294 = _T_12293 ? _T_10366_1 : _T_12292; // @[Mux.scala 46:16:@11593.4]
  assign _T_12295 = 5'h1 == _T_11317_21; // @[Mux.scala 46:19:@11594.4]
  assign _T_12296 = _T_12295 ? _T_10366_0 : _T_12294; // @[Mux.scala 46:16:@11595.4]
  assign _T_12321 = 5'h17 == _T_11317_22; // @[Mux.scala 46:19:@11597.4]
  assign _T_12322 = _T_12321 ? _T_10366_22 : 8'h0; // @[Mux.scala 46:16:@11598.4]
  assign _T_12323 = 5'h16 == _T_11317_22; // @[Mux.scala 46:19:@11599.4]
  assign _T_12324 = _T_12323 ? _T_10366_21 : _T_12322; // @[Mux.scala 46:16:@11600.4]
  assign _T_12325 = 5'h15 == _T_11317_22; // @[Mux.scala 46:19:@11601.4]
  assign _T_12326 = _T_12325 ? _T_10366_20 : _T_12324; // @[Mux.scala 46:16:@11602.4]
  assign _T_12327 = 5'h14 == _T_11317_22; // @[Mux.scala 46:19:@11603.4]
  assign _T_12328 = _T_12327 ? _T_10366_19 : _T_12326; // @[Mux.scala 46:16:@11604.4]
  assign _T_12329 = 5'h13 == _T_11317_22; // @[Mux.scala 46:19:@11605.4]
  assign _T_12330 = _T_12329 ? _T_10366_18 : _T_12328; // @[Mux.scala 46:16:@11606.4]
  assign _T_12331 = 5'h12 == _T_11317_22; // @[Mux.scala 46:19:@11607.4]
  assign _T_12332 = _T_12331 ? _T_10366_17 : _T_12330; // @[Mux.scala 46:16:@11608.4]
  assign _T_12333 = 5'h11 == _T_11317_22; // @[Mux.scala 46:19:@11609.4]
  assign _T_12334 = _T_12333 ? _T_10366_16 : _T_12332; // @[Mux.scala 46:16:@11610.4]
  assign _T_12335 = 5'h10 == _T_11317_22; // @[Mux.scala 46:19:@11611.4]
  assign _T_12336 = _T_12335 ? _T_10366_15 : _T_12334; // @[Mux.scala 46:16:@11612.4]
  assign _T_12337 = 5'hf == _T_11317_22; // @[Mux.scala 46:19:@11613.4]
  assign _T_12338 = _T_12337 ? _T_10366_14 : _T_12336; // @[Mux.scala 46:16:@11614.4]
  assign _T_12339 = 5'he == _T_11317_22; // @[Mux.scala 46:19:@11615.4]
  assign _T_12340 = _T_12339 ? _T_10366_13 : _T_12338; // @[Mux.scala 46:16:@11616.4]
  assign _T_12341 = 5'hd == _T_11317_22; // @[Mux.scala 46:19:@11617.4]
  assign _T_12342 = _T_12341 ? _T_10366_12 : _T_12340; // @[Mux.scala 46:16:@11618.4]
  assign _T_12343 = 5'hc == _T_11317_22; // @[Mux.scala 46:19:@11619.4]
  assign _T_12344 = _T_12343 ? _T_10366_11 : _T_12342; // @[Mux.scala 46:16:@11620.4]
  assign _T_12345 = 5'hb == _T_11317_22; // @[Mux.scala 46:19:@11621.4]
  assign _T_12346 = _T_12345 ? _T_10366_10 : _T_12344; // @[Mux.scala 46:16:@11622.4]
  assign _T_12347 = 5'ha == _T_11317_22; // @[Mux.scala 46:19:@11623.4]
  assign _T_12348 = _T_12347 ? _T_10366_9 : _T_12346; // @[Mux.scala 46:16:@11624.4]
  assign _T_12349 = 5'h9 == _T_11317_22; // @[Mux.scala 46:19:@11625.4]
  assign _T_12350 = _T_12349 ? _T_10366_8 : _T_12348; // @[Mux.scala 46:16:@11626.4]
  assign _T_12351 = 5'h8 == _T_11317_22; // @[Mux.scala 46:19:@11627.4]
  assign _T_12352 = _T_12351 ? _T_10366_7 : _T_12350; // @[Mux.scala 46:16:@11628.4]
  assign _T_12353 = 5'h7 == _T_11317_22; // @[Mux.scala 46:19:@11629.4]
  assign _T_12354 = _T_12353 ? _T_10366_6 : _T_12352; // @[Mux.scala 46:16:@11630.4]
  assign _T_12355 = 5'h6 == _T_11317_22; // @[Mux.scala 46:19:@11631.4]
  assign _T_12356 = _T_12355 ? _T_10366_5 : _T_12354; // @[Mux.scala 46:16:@11632.4]
  assign _T_12357 = 5'h5 == _T_11317_22; // @[Mux.scala 46:19:@11633.4]
  assign _T_12358 = _T_12357 ? _T_10366_4 : _T_12356; // @[Mux.scala 46:16:@11634.4]
  assign _T_12359 = 5'h4 == _T_11317_22; // @[Mux.scala 46:19:@11635.4]
  assign _T_12360 = _T_12359 ? _T_10366_3 : _T_12358; // @[Mux.scala 46:16:@11636.4]
  assign _T_12361 = 5'h3 == _T_11317_22; // @[Mux.scala 46:19:@11637.4]
  assign _T_12362 = _T_12361 ? _T_10366_2 : _T_12360; // @[Mux.scala 46:16:@11638.4]
  assign _T_12363 = 5'h2 == _T_11317_22; // @[Mux.scala 46:19:@11639.4]
  assign _T_12364 = _T_12363 ? _T_10366_1 : _T_12362; // @[Mux.scala 46:16:@11640.4]
  assign _T_12365 = 5'h1 == _T_11317_22; // @[Mux.scala 46:19:@11641.4]
  assign _T_12366 = _T_12365 ? _T_10366_0 : _T_12364; // @[Mux.scala 46:16:@11642.4]
  assign _T_12392 = 5'h18 == _T_11317_23; // @[Mux.scala 46:19:@11644.4]
  assign _T_12393 = _T_12392 ? _T_10366_23 : 8'h0; // @[Mux.scala 46:16:@11645.4]
  assign _T_12394 = 5'h17 == _T_11317_23; // @[Mux.scala 46:19:@11646.4]
  assign _T_12395 = _T_12394 ? _T_10366_22 : _T_12393; // @[Mux.scala 46:16:@11647.4]
  assign _T_12396 = 5'h16 == _T_11317_23; // @[Mux.scala 46:19:@11648.4]
  assign _T_12397 = _T_12396 ? _T_10366_21 : _T_12395; // @[Mux.scala 46:16:@11649.4]
  assign _T_12398 = 5'h15 == _T_11317_23; // @[Mux.scala 46:19:@11650.4]
  assign _T_12399 = _T_12398 ? _T_10366_20 : _T_12397; // @[Mux.scala 46:16:@11651.4]
  assign _T_12400 = 5'h14 == _T_11317_23; // @[Mux.scala 46:19:@11652.4]
  assign _T_12401 = _T_12400 ? _T_10366_19 : _T_12399; // @[Mux.scala 46:16:@11653.4]
  assign _T_12402 = 5'h13 == _T_11317_23; // @[Mux.scala 46:19:@11654.4]
  assign _T_12403 = _T_12402 ? _T_10366_18 : _T_12401; // @[Mux.scala 46:16:@11655.4]
  assign _T_12404 = 5'h12 == _T_11317_23; // @[Mux.scala 46:19:@11656.4]
  assign _T_12405 = _T_12404 ? _T_10366_17 : _T_12403; // @[Mux.scala 46:16:@11657.4]
  assign _T_12406 = 5'h11 == _T_11317_23; // @[Mux.scala 46:19:@11658.4]
  assign _T_12407 = _T_12406 ? _T_10366_16 : _T_12405; // @[Mux.scala 46:16:@11659.4]
  assign _T_12408 = 5'h10 == _T_11317_23; // @[Mux.scala 46:19:@11660.4]
  assign _T_12409 = _T_12408 ? _T_10366_15 : _T_12407; // @[Mux.scala 46:16:@11661.4]
  assign _T_12410 = 5'hf == _T_11317_23; // @[Mux.scala 46:19:@11662.4]
  assign _T_12411 = _T_12410 ? _T_10366_14 : _T_12409; // @[Mux.scala 46:16:@11663.4]
  assign _T_12412 = 5'he == _T_11317_23; // @[Mux.scala 46:19:@11664.4]
  assign _T_12413 = _T_12412 ? _T_10366_13 : _T_12411; // @[Mux.scala 46:16:@11665.4]
  assign _T_12414 = 5'hd == _T_11317_23; // @[Mux.scala 46:19:@11666.4]
  assign _T_12415 = _T_12414 ? _T_10366_12 : _T_12413; // @[Mux.scala 46:16:@11667.4]
  assign _T_12416 = 5'hc == _T_11317_23; // @[Mux.scala 46:19:@11668.4]
  assign _T_12417 = _T_12416 ? _T_10366_11 : _T_12415; // @[Mux.scala 46:16:@11669.4]
  assign _T_12418 = 5'hb == _T_11317_23; // @[Mux.scala 46:19:@11670.4]
  assign _T_12419 = _T_12418 ? _T_10366_10 : _T_12417; // @[Mux.scala 46:16:@11671.4]
  assign _T_12420 = 5'ha == _T_11317_23; // @[Mux.scala 46:19:@11672.4]
  assign _T_12421 = _T_12420 ? _T_10366_9 : _T_12419; // @[Mux.scala 46:16:@11673.4]
  assign _T_12422 = 5'h9 == _T_11317_23; // @[Mux.scala 46:19:@11674.4]
  assign _T_12423 = _T_12422 ? _T_10366_8 : _T_12421; // @[Mux.scala 46:16:@11675.4]
  assign _T_12424 = 5'h8 == _T_11317_23; // @[Mux.scala 46:19:@11676.4]
  assign _T_12425 = _T_12424 ? _T_10366_7 : _T_12423; // @[Mux.scala 46:16:@11677.4]
  assign _T_12426 = 5'h7 == _T_11317_23; // @[Mux.scala 46:19:@11678.4]
  assign _T_12427 = _T_12426 ? _T_10366_6 : _T_12425; // @[Mux.scala 46:16:@11679.4]
  assign _T_12428 = 5'h6 == _T_11317_23; // @[Mux.scala 46:19:@11680.4]
  assign _T_12429 = _T_12428 ? _T_10366_5 : _T_12427; // @[Mux.scala 46:16:@11681.4]
  assign _T_12430 = 5'h5 == _T_11317_23; // @[Mux.scala 46:19:@11682.4]
  assign _T_12431 = _T_12430 ? _T_10366_4 : _T_12429; // @[Mux.scala 46:16:@11683.4]
  assign _T_12432 = 5'h4 == _T_11317_23; // @[Mux.scala 46:19:@11684.4]
  assign _T_12433 = _T_12432 ? _T_10366_3 : _T_12431; // @[Mux.scala 46:16:@11685.4]
  assign _T_12434 = 5'h3 == _T_11317_23; // @[Mux.scala 46:19:@11686.4]
  assign _T_12435 = _T_12434 ? _T_10366_2 : _T_12433; // @[Mux.scala 46:16:@11687.4]
  assign _T_12436 = 5'h2 == _T_11317_23; // @[Mux.scala 46:19:@11688.4]
  assign _T_12437 = _T_12436 ? _T_10366_1 : _T_12435; // @[Mux.scala 46:16:@11689.4]
  assign _T_12438 = 5'h1 == _T_11317_23; // @[Mux.scala 46:19:@11690.4]
  assign _T_12439 = _T_12438 ? _T_10366_0 : _T_12437; // @[Mux.scala 46:16:@11691.4]
  assign _T_12466 = 5'h19 == _T_11317_24; // @[Mux.scala 46:19:@11693.4]
  assign _T_12467 = _T_12466 ? _T_10366_24 : 8'h0; // @[Mux.scala 46:16:@11694.4]
  assign _T_12468 = 5'h18 == _T_11317_24; // @[Mux.scala 46:19:@11695.4]
  assign _T_12469 = _T_12468 ? _T_10366_23 : _T_12467; // @[Mux.scala 46:16:@11696.4]
  assign _T_12470 = 5'h17 == _T_11317_24; // @[Mux.scala 46:19:@11697.4]
  assign _T_12471 = _T_12470 ? _T_10366_22 : _T_12469; // @[Mux.scala 46:16:@11698.4]
  assign _T_12472 = 5'h16 == _T_11317_24; // @[Mux.scala 46:19:@11699.4]
  assign _T_12473 = _T_12472 ? _T_10366_21 : _T_12471; // @[Mux.scala 46:16:@11700.4]
  assign _T_12474 = 5'h15 == _T_11317_24; // @[Mux.scala 46:19:@11701.4]
  assign _T_12475 = _T_12474 ? _T_10366_20 : _T_12473; // @[Mux.scala 46:16:@11702.4]
  assign _T_12476 = 5'h14 == _T_11317_24; // @[Mux.scala 46:19:@11703.4]
  assign _T_12477 = _T_12476 ? _T_10366_19 : _T_12475; // @[Mux.scala 46:16:@11704.4]
  assign _T_12478 = 5'h13 == _T_11317_24; // @[Mux.scala 46:19:@11705.4]
  assign _T_12479 = _T_12478 ? _T_10366_18 : _T_12477; // @[Mux.scala 46:16:@11706.4]
  assign _T_12480 = 5'h12 == _T_11317_24; // @[Mux.scala 46:19:@11707.4]
  assign _T_12481 = _T_12480 ? _T_10366_17 : _T_12479; // @[Mux.scala 46:16:@11708.4]
  assign _T_12482 = 5'h11 == _T_11317_24; // @[Mux.scala 46:19:@11709.4]
  assign _T_12483 = _T_12482 ? _T_10366_16 : _T_12481; // @[Mux.scala 46:16:@11710.4]
  assign _T_12484 = 5'h10 == _T_11317_24; // @[Mux.scala 46:19:@11711.4]
  assign _T_12485 = _T_12484 ? _T_10366_15 : _T_12483; // @[Mux.scala 46:16:@11712.4]
  assign _T_12486 = 5'hf == _T_11317_24; // @[Mux.scala 46:19:@11713.4]
  assign _T_12487 = _T_12486 ? _T_10366_14 : _T_12485; // @[Mux.scala 46:16:@11714.4]
  assign _T_12488 = 5'he == _T_11317_24; // @[Mux.scala 46:19:@11715.4]
  assign _T_12489 = _T_12488 ? _T_10366_13 : _T_12487; // @[Mux.scala 46:16:@11716.4]
  assign _T_12490 = 5'hd == _T_11317_24; // @[Mux.scala 46:19:@11717.4]
  assign _T_12491 = _T_12490 ? _T_10366_12 : _T_12489; // @[Mux.scala 46:16:@11718.4]
  assign _T_12492 = 5'hc == _T_11317_24; // @[Mux.scala 46:19:@11719.4]
  assign _T_12493 = _T_12492 ? _T_10366_11 : _T_12491; // @[Mux.scala 46:16:@11720.4]
  assign _T_12494 = 5'hb == _T_11317_24; // @[Mux.scala 46:19:@11721.4]
  assign _T_12495 = _T_12494 ? _T_10366_10 : _T_12493; // @[Mux.scala 46:16:@11722.4]
  assign _T_12496 = 5'ha == _T_11317_24; // @[Mux.scala 46:19:@11723.4]
  assign _T_12497 = _T_12496 ? _T_10366_9 : _T_12495; // @[Mux.scala 46:16:@11724.4]
  assign _T_12498 = 5'h9 == _T_11317_24; // @[Mux.scala 46:19:@11725.4]
  assign _T_12499 = _T_12498 ? _T_10366_8 : _T_12497; // @[Mux.scala 46:16:@11726.4]
  assign _T_12500 = 5'h8 == _T_11317_24; // @[Mux.scala 46:19:@11727.4]
  assign _T_12501 = _T_12500 ? _T_10366_7 : _T_12499; // @[Mux.scala 46:16:@11728.4]
  assign _T_12502 = 5'h7 == _T_11317_24; // @[Mux.scala 46:19:@11729.4]
  assign _T_12503 = _T_12502 ? _T_10366_6 : _T_12501; // @[Mux.scala 46:16:@11730.4]
  assign _T_12504 = 5'h6 == _T_11317_24; // @[Mux.scala 46:19:@11731.4]
  assign _T_12505 = _T_12504 ? _T_10366_5 : _T_12503; // @[Mux.scala 46:16:@11732.4]
  assign _T_12506 = 5'h5 == _T_11317_24; // @[Mux.scala 46:19:@11733.4]
  assign _T_12507 = _T_12506 ? _T_10366_4 : _T_12505; // @[Mux.scala 46:16:@11734.4]
  assign _T_12508 = 5'h4 == _T_11317_24; // @[Mux.scala 46:19:@11735.4]
  assign _T_12509 = _T_12508 ? _T_10366_3 : _T_12507; // @[Mux.scala 46:16:@11736.4]
  assign _T_12510 = 5'h3 == _T_11317_24; // @[Mux.scala 46:19:@11737.4]
  assign _T_12511 = _T_12510 ? _T_10366_2 : _T_12509; // @[Mux.scala 46:16:@11738.4]
  assign _T_12512 = 5'h2 == _T_11317_24; // @[Mux.scala 46:19:@11739.4]
  assign _T_12513 = _T_12512 ? _T_10366_1 : _T_12511; // @[Mux.scala 46:16:@11740.4]
  assign _T_12514 = 5'h1 == _T_11317_24; // @[Mux.scala 46:19:@11741.4]
  assign _T_12515 = _T_12514 ? _T_10366_0 : _T_12513; // @[Mux.scala 46:16:@11742.4]
  assign _T_12543 = 5'h1a == _T_11317_25; // @[Mux.scala 46:19:@11744.4]
  assign _T_12544 = _T_12543 ? _T_10366_25 : 8'h0; // @[Mux.scala 46:16:@11745.4]
  assign _T_12545 = 5'h19 == _T_11317_25; // @[Mux.scala 46:19:@11746.4]
  assign _T_12546 = _T_12545 ? _T_10366_24 : _T_12544; // @[Mux.scala 46:16:@11747.4]
  assign _T_12547 = 5'h18 == _T_11317_25; // @[Mux.scala 46:19:@11748.4]
  assign _T_12548 = _T_12547 ? _T_10366_23 : _T_12546; // @[Mux.scala 46:16:@11749.4]
  assign _T_12549 = 5'h17 == _T_11317_25; // @[Mux.scala 46:19:@11750.4]
  assign _T_12550 = _T_12549 ? _T_10366_22 : _T_12548; // @[Mux.scala 46:16:@11751.4]
  assign _T_12551 = 5'h16 == _T_11317_25; // @[Mux.scala 46:19:@11752.4]
  assign _T_12552 = _T_12551 ? _T_10366_21 : _T_12550; // @[Mux.scala 46:16:@11753.4]
  assign _T_12553 = 5'h15 == _T_11317_25; // @[Mux.scala 46:19:@11754.4]
  assign _T_12554 = _T_12553 ? _T_10366_20 : _T_12552; // @[Mux.scala 46:16:@11755.4]
  assign _T_12555 = 5'h14 == _T_11317_25; // @[Mux.scala 46:19:@11756.4]
  assign _T_12556 = _T_12555 ? _T_10366_19 : _T_12554; // @[Mux.scala 46:16:@11757.4]
  assign _T_12557 = 5'h13 == _T_11317_25; // @[Mux.scala 46:19:@11758.4]
  assign _T_12558 = _T_12557 ? _T_10366_18 : _T_12556; // @[Mux.scala 46:16:@11759.4]
  assign _T_12559 = 5'h12 == _T_11317_25; // @[Mux.scala 46:19:@11760.4]
  assign _T_12560 = _T_12559 ? _T_10366_17 : _T_12558; // @[Mux.scala 46:16:@11761.4]
  assign _T_12561 = 5'h11 == _T_11317_25; // @[Mux.scala 46:19:@11762.4]
  assign _T_12562 = _T_12561 ? _T_10366_16 : _T_12560; // @[Mux.scala 46:16:@11763.4]
  assign _T_12563 = 5'h10 == _T_11317_25; // @[Mux.scala 46:19:@11764.4]
  assign _T_12564 = _T_12563 ? _T_10366_15 : _T_12562; // @[Mux.scala 46:16:@11765.4]
  assign _T_12565 = 5'hf == _T_11317_25; // @[Mux.scala 46:19:@11766.4]
  assign _T_12566 = _T_12565 ? _T_10366_14 : _T_12564; // @[Mux.scala 46:16:@11767.4]
  assign _T_12567 = 5'he == _T_11317_25; // @[Mux.scala 46:19:@11768.4]
  assign _T_12568 = _T_12567 ? _T_10366_13 : _T_12566; // @[Mux.scala 46:16:@11769.4]
  assign _T_12569 = 5'hd == _T_11317_25; // @[Mux.scala 46:19:@11770.4]
  assign _T_12570 = _T_12569 ? _T_10366_12 : _T_12568; // @[Mux.scala 46:16:@11771.4]
  assign _T_12571 = 5'hc == _T_11317_25; // @[Mux.scala 46:19:@11772.4]
  assign _T_12572 = _T_12571 ? _T_10366_11 : _T_12570; // @[Mux.scala 46:16:@11773.4]
  assign _T_12573 = 5'hb == _T_11317_25; // @[Mux.scala 46:19:@11774.4]
  assign _T_12574 = _T_12573 ? _T_10366_10 : _T_12572; // @[Mux.scala 46:16:@11775.4]
  assign _T_12575 = 5'ha == _T_11317_25; // @[Mux.scala 46:19:@11776.4]
  assign _T_12576 = _T_12575 ? _T_10366_9 : _T_12574; // @[Mux.scala 46:16:@11777.4]
  assign _T_12577 = 5'h9 == _T_11317_25; // @[Mux.scala 46:19:@11778.4]
  assign _T_12578 = _T_12577 ? _T_10366_8 : _T_12576; // @[Mux.scala 46:16:@11779.4]
  assign _T_12579 = 5'h8 == _T_11317_25; // @[Mux.scala 46:19:@11780.4]
  assign _T_12580 = _T_12579 ? _T_10366_7 : _T_12578; // @[Mux.scala 46:16:@11781.4]
  assign _T_12581 = 5'h7 == _T_11317_25; // @[Mux.scala 46:19:@11782.4]
  assign _T_12582 = _T_12581 ? _T_10366_6 : _T_12580; // @[Mux.scala 46:16:@11783.4]
  assign _T_12583 = 5'h6 == _T_11317_25; // @[Mux.scala 46:19:@11784.4]
  assign _T_12584 = _T_12583 ? _T_10366_5 : _T_12582; // @[Mux.scala 46:16:@11785.4]
  assign _T_12585 = 5'h5 == _T_11317_25; // @[Mux.scala 46:19:@11786.4]
  assign _T_12586 = _T_12585 ? _T_10366_4 : _T_12584; // @[Mux.scala 46:16:@11787.4]
  assign _T_12587 = 5'h4 == _T_11317_25; // @[Mux.scala 46:19:@11788.4]
  assign _T_12588 = _T_12587 ? _T_10366_3 : _T_12586; // @[Mux.scala 46:16:@11789.4]
  assign _T_12589 = 5'h3 == _T_11317_25; // @[Mux.scala 46:19:@11790.4]
  assign _T_12590 = _T_12589 ? _T_10366_2 : _T_12588; // @[Mux.scala 46:16:@11791.4]
  assign _T_12591 = 5'h2 == _T_11317_25; // @[Mux.scala 46:19:@11792.4]
  assign _T_12592 = _T_12591 ? _T_10366_1 : _T_12590; // @[Mux.scala 46:16:@11793.4]
  assign _T_12593 = 5'h1 == _T_11317_25; // @[Mux.scala 46:19:@11794.4]
  assign _T_12594 = _T_12593 ? _T_10366_0 : _T_12592; // @[Mux.scala 46:16:@11795.4]
  assign _T_12623 = 5'h1b == _T_11317_26; // @[Mux.scala 46:19:@11797.4]
  assign _T_12624 = _T_12623 ? _T_10366_26 : 8'h0; // @[Mux.scala 46:16:@11798.4]
  assign _T_12625 = 5'h1a == _T_11317_26; // @[Mux.scala 46:19:@11799.4]
  assign _T_12626 = _T_12625 ? _T_10366_25 : _T_12624; // @[Mux.scala 46:16:@11800.4]
  assign _T_12627 = 5'h19 == _T_11317_26; // @[Mux.scala 46:19:@11801.4]
  assign _T_12628 = _T_12627 ? _T_10366_24 : _T_12626; // @[Mux.scala 46:16:@11802.4]
  assign _T_12629 = 5'h18 == _T_11317_26; // @[Mux.scala 46:19:@11803.4]
  assign _T_12630 = _T_12629 ? _T_10366_23 : _T_12628; // @[Mux.scala 46:16:@11804.4]
  assign _T_12631 = 5'h17 == _T_11317_26; // @[Mux.scala 46:19:@11805.4]
  assign _T_12632 = _T_12631 ? _T_10366_22 : _T_12630; // @[Mux.scala 46:16:@11806.4]
  assign _T_12633 = 5'h16 == _T_11317_26; // @[Mux.scala 46:19:@11807.4]
  assign _T_12634 = _T_12633 ? _T_10366_21 : _T_12632; // @[Mux.scala 46:16:@11808.4]
  assign _T_12635 = 5'h15 == _T_11317_26; // @[Mux.scala 46:19:@11809.4]
  assign _T_12636 = _T_12635 ? _T_10366_20 : _T_12634; // @[Mux.scala 46:16:@11810.4]
  assign _T_12637 = 5'h14 == _T_11317_26; // @[Mux.scala 46:19:@11811.4]
  assign _T_12638 = _T_12637 ? _T_10366_19 : _T_12636; // @[Mux.scala 46:16:@11812.4]
  assign _T_12639 = 5'h13 == _T_11317_26; // @[Mux.scala 46:19:@11813.4]
  assign _T_12640 = _T_12639 ? _T_10366_18 : _T_12638; // @[Mux.scala 46:16:@11814.4]
  assign _T_12641 = 5'h12 == _T_11317_26; // @[Mux.scala 46:19:@11815.4]
  assign _T_12642 = _T_12641 ? _T_10366_17 : _T_12640; // @[Mux.scala 46:16:@11816.4]
  assign _T_12643 = 5'h11 == _T_11317_26; // @[Mux.scala 46:19:@11817.4]
  assign _T_12644 = _T_12643 ? _T_10366_16 : _T_12642; // @[Mux.scala 46:16:@11818.4]
  assign _T_12645 = 5'h10 == _T_11317_26; // @[Mux.scala 46:19:@11819.4]
  assign _T_12646 = _T_12645 ? _T_10366_15 : _T_12644; // @[Mux.scala 46:16:@11820.4]
  assign _T_12647 = 5'hf == _T_11317_26; // @[Mux.scala 46:19:@11821.4]
  assign _T_12648 = _T_12647 ? _T_10366_14 : _T_12646; // @[Mux.scala 46:16:@11822.4]
  assign _T_12649 = 5'he == _T_11317_26; // @[Mux.scala 46:19:@11823.4]
  assign _T_12650 = _T_12649 ? _T_10366_13 : _T_12648; // @[Mux.scala 46:16:@11824.4]
  assign _T_12651 = 5'hd == _T_11317_26; // @[Mux.scala 46:19:@11825.4]
  assign _T_12652 = _T_12651 ? _T_10366_12 : _T_12650; // @[Mux.scala 46:16:@11826.4]
  assign _T_12653 = 5'hc == _T_11317_26; // @[Mux.scala 46:19:@11827.4]
  assign _T_12654 = _T_12653 ? _T_10366_11 : _T_12652; // @[Mux.scala 46:16:@11828.4]
  assign _T_12655 = 5'hb == _T_11317_26; // @[Mux.scala 46:19:@11829.4]
  assign _T_12656 = _T_12655 ? _T_10366_10 : _T_12654; // @[Mux.scala 46:16:@11830.4]
  assign _T_12657 = 5'ha == _T_11317_26; // @[Mux.scala 46:19:@11831.4]
  assign _T_12658 = _T_12657 ? _T_10366_9 : _T_12656; // @[Mux.scala 46:16:@11832.4]
  assign _T_12659 = 5'h9 == _T_11317_26; // @[Mux.scala 46:19:@11833.4]
  assign _T_12660 = _T_12659 ? _T_10366_8 : _T_12658; // @[Mux.scala 46:16:@11834.4]
  assign _T_12661 = 5'h8 == _T_11317_26; // @[Mux.scala 46:19:@11835.4]
  assign _T_12662 = _T_12661 ? _T_10366_7 : _T_12660; // @[Mux.scala 46:16:@11836.4]
  assign _T_12663 = 5'h7 == _T_11317_26; // @[Mux.scala 46:19:@11837.4]
  assign _T_12664 = _T_12663 ? _T_10366_6 : _T_12662; // @[Mux.scala 46:16:@11838.4]
  assign _T_12665 = 5'h6 == _T_11317_26; // @[Mux.scala 46:19:@11839.4]
  assign _T_12666 = _T_12665 ? _T_10366_5 : _T_12664; // @[Mux.scala 46:16:@11840.4]
  assign _T_12667 = 5'h5 == _T_11317_26; // @[Mux.scala 46:19:@11841.4]
  assign _T_12668 = _T_12667 ? _T_10366_4 : _T_12666; // @[Mux.scala 46:16:@11842.4]
  assign _T_12669 = 5'h4 == _T_11317_26; // @[Mux.scala 46:19:@11843.4]
  assign _T_12670 = _T_12669 ? _T_10366_3 : _T_12668; // @[Mux.scala 46:16:@11844.4]
  assign _T_12671 = 5'h3 == _T_11317_26; // @[Mux.scala 46:19:@11845.4]
  assign _T_12672 = _T_12671 ? _T_10366_2 : _T_12670; // @[Mux.scala 46:16:@11846.4]
  assign _T_12673 = 5'h2 == _T_11317_26; // @[Mux.scala 46:19:@11847.4]
  assign _T_12674 = _T_12673 ? _T_10366_1 : _T_12672; // @[Mux.scala 46:16:@11848.4]
  assign _T_12675 = 5'h1 == _T_11317_26; // @[Mux.scala 46:19:@11849.4]
  assign _T_12676 = _T_12675 ? _T_10366_0 : _T_12674; // @[Mux.scala 46:16:@11850.4]
  assign _T_12706 = 5'h1c == _T_11317_27; // @[Mux.scala 46:19:@11852.4]
  assign _T_12707 = _T_12706 ? _T_10366_27 : 8'h0; // @[Mux.scala 46:16:@11853.4]
  assign _T_12708 = 5'h1b == _T_11317_27; // @[Mux.scala 46:19:@11854.4]
  assign _T_12709 = _T_12708 ? _T_10366_26 : _T_12707; // @[Mux.scala 46:16:@11855.4]
  assign _T_12710 = 5'h1a == _T_11317_27; // @[Mux.scala 46:19:@11856.4]
  assign _T_12711 = _T_12710 ? _T_10366_25 : _T_12709; // @[Mux.scala 46:16:@11857.4]
  assign _T_12712 = 5'h19 == _T_11317_27; // @[Mux.scala 46:19:@11858.4]
  assign _T_12713 = _T_12712 ? _T_10366_24 : _T_12711; // @[Mux.scala 46:16:@11859.4]
  assign _T_12714 = 5'h18 == _T_11317_27; // @[Mux.scala 46:19:@11860.4]
  assign _T_12715 = _T_12714 ? _T_10366_23 : _T_12713; // @[Mux.scala 46:16:@11861.4]
  assign _T_12716 = 5'h17 == _T_11317_27; // @[Mux.scala 46:19:@11862.4]
  assign _T_12717 = _T_12716 ? _T_10366_22 : _T_12715; // @[Mux.scala 46:16:@11863.4]
  assign _T_12718 = 5'h16 == _T_11317_27; // @[Mux.scala 46:19:@11864.4]
  assign _T_12719 = _T_12718 ? _T_10366_21 : _T_12717; // @[Mux.scala 46:16:@11865.4]
  assign _T_12720 = 5'h15 == _T_11317_27; // @[Mux.scala 46:19:@11866.4]
  assign _T_12721 = _T_12720 ? _T_10366_20 : _T_12719; // @[Mux.scala 46:16:@11867.4]
  assign _T_12722 = 5'h14 == _T_11317_27; // @[Mux.scala 46:19:@11868.4]
  assign _T_12723 = _T_12722 ? _T_10366_19 : _T_12721; // @[Mux.scala 46:16:@11869.4]
  assign _T_12724 = 5'h13 == _T_11317_27; // @[Mux.scala 46:19:@11870.4]
  assign _T_12725 = _T_12724 ? _T_10366_18 : _T_12723; // @[Mux.scala 46:16:@11871.4]
  assign _T_12726 = 5'h12 == _T_11317_27; // @[Mux.scala 46:19:@11872.4]
  assign _T_12727 = _T_12726 ? _T_10366_17 : _T_12725; // @[Mux.scala 46:16:@11873.4]
  assign _T_12728 = 5'h11 == _T_11317_27; // @[Mux.scala 46:19:@11874.4]
  assign _T_12729 = _T_12728 ? _T_10366_16 : _T_12727; // @[Mux.scala 46:16:@11875.4]
  assign _T_12730 = 5'h10 == _T_11317_27; // @[Mux.scala 46:19:@11876.4]
  assign _T_12731 = _T_12730 ? _T_10366_15 : _T_12729; // @[Mux.scala 46:16:@11877.4]
  assign _T_12732 = 5'hf == _T_11317_27; // @[Mux.scala 46:19:@11878.4]
  assign _T_12733 = _T_12732 ? _T_10366_14 : _T_12731; // @[Mux.scala 46:16:@11879.4]
  assign _T_12734 = 5'he == _T_11317_27; // @[Mux.scala 46:19:@11880.4]
  assign _T_12735 = _T_12734 ? _T_10366_13 : _T_12733; // @[Mux.scala 46:16:@11881.4]
  assign _T_12736 = 5'hd == _T_11317_27; // @[Mux.scala 46:19:@11882.4]
  assign _T_12737 = _T_12736 ? _T_10366_12 : _T_12735; // @[Mux.scala 46:16:@11883.4]
  assign _T_12738 = 5'hc == _T_11317_27; // @[Mux.scala 46:19:@11884.4]
  assign _T_12739 = _T_12738 ? _T_10366_11 : _T_12737; // @[Mux.scala 46:16:@11885.4]
  assign _T_12740 = 5'hb == _T_11317_27; // @[Mux.scala 46:19:@11886.4]
  assign _T_12741 = _T_12740 ? _T_10366_10 : _T_12739; // @[Mux.scala 46:16:@11887.4]
  assign _T_12742 = 5'ha == _T_11317_27; // @[Mux.scala 46:19:@11888.4]
  assign _T_12743 = _T_12742 ? _T_10366_9 : _T_12741; // @[Mux.scala 46:16:@11889.4]
  assign _T_12744 = 5'h9 == _T_11317_27; // @[Mux.scala 46:19:@11890.4]
  assign _T_12745 = _T_12744 ? _T_10366_8 : _T_12743; // @[Mux.scala 46:16:@11891.4]
  assign _T_12746 = 5'h8 == _T_11317_27; // @[Mux.scala 46:19:@11892.4]
  assign _T_12747 = _T_12746 ? _T_10366_7 : _T_12745; // @[Mux.scala 46:16:@11893.4]
  assign _T_12748 = 5'h7 == _T_11317_27; // @[Mux.scala 46:19:@11894.4]
  assign _T_12749 = _T_12748 ? _T_10366_6 : _T_12747; // @[Mux.scala 46:16:@11895.4]
  assign _T_12750 = 5'h6 == _T_11317_27; // @[Mux.scala 46:19:@11896.4]
  assign _T_12751 = _T_12750 ? _T_10366_5 : _T_12749; // @[Mux.scala 46:16:@11897.4]
  assign _T_12752 = 5'h5 == _T_11317_27; // @[Mux.scala 46:19:@11898.4]
  assign _T_12753 = _T_12752 ? _T_10366_4 : _T_12751; // @[Mux.scala 46:16:@11899.4]
  assign _T_12754 = 5'h4 == _T_11317_27; // @[Mux.scala 46:19:@11900.4]
  assign _T_12755 = _T_12754 ? _T_10366_3 : _T_12753; // @[Mux.scala 46:16:@11901.4]
  assign _T_12756 = 5'h3 == _T_11317_27; // @[Mux.scala 46:19:@11902.4]
  assign _T_12757 = _T_12756 ? _T_10366_2 : _T_12755; // @[Mux.scala 46:16:@11903.4]
  assign _T_12758 = 5'h2 == _T_11317_27; // @[Mux.scala 46:19:@11904.4]
  assign _T_12759 = _T_12758 ? _T_10366_1 : _T_12757; // @[Mux.scala 46:16:@11905.4]
  assign _T_12760 = 5'h1 == _T_11317_27; // @[Mux.scala 46:19:@11906.4]
  assign _T_12761 = _T_12760 ? _T_10366_0 : _T_12759; // @[Mux.scala 46:16:@11907.4]
  assign _T_12792 = 5'h1d == _T_11317_28; // @[Mux.scala 46:19:@11909.4]
  assign _T_12793 = _T_12792 ? _T_10366_28 : 8'h0; // @[Mux.scala 46:16:@11910.4]
  assign _T_12794 = 5'h1c == _T_11317_28; // @[Mux.scala 46:19:@11911.4]
  assign _T_12795 = _T_12794 ? _T_10366_27 : _T_12793; // @[Mux.scala 46:16:@11912.4]
  assign _T_12796 = 5'h1b == _T_11317_28; // @[Mux.scala 46:19:@11913.4]
  assign _T_12797 = _T_12796 ? _T_10366_26 : _T_12795; // @[Mux.scala 46:16:@11914.4]
  assign _T_12798 = 5'h1a == _T_11317_28; // @[Mux.scala 46:19:@11915.4]
  assign _T_12799 = _T_12798 ? _T_10366_25 : _T_12797; // @[Mux.scala 46:16:@11916.4]
  assign _T_12800 = 5'h19 == _T_11317_28; // @[Mux.scala 46:19:@11917.4]
  assign _T_12801 = _T_12800 ? _T_10366_24 : _T_12799; // @[Mux.scala 46:16:@11918.4]
  assign _T_12802 = 5'h18 == _T_11317_28; // @[Mux.scala 46:19:@11919.4]
  assign _T_12803 = _T_12802 ? _T_10366_23 : _T_12801; // @[Mux.scala 46:16:@11920.4]
  assign _T_12804 = 5'h17 == _T_11317_28; // @[Mux.scala 46:19:@11921.4]
  assign _T_12805 = _T_12804 ? _T_10366_22 : _T_12803; // @[Mux.scala 46:16:@11922.4]
  assign _T_12806 = 5'h16 == _T_11317_28; // @[Mux.scala 46:19:@11923.4]
  assign _T_12807 = _T_12806 ? _T_10366_21 : _T_12805; // @[Mux.scala 46:16:@11924.4]
  assign _T_12808 = 5'h15 == _T_11317_28; // @[Mux.scala 46:19:@11925.4]
  assign _T_12809 = _T_12808 ? _T_10366_20 : _T_12807; // @[Mux.scala 46:16:@11926.4]
  assign _T_12810 = 5'h14 == _T_11317_28; // @[Mux.scala 46:19:@11927.4]
  assign _T_12811 = _T_12810 ? _T_10366_19 : _T_12809; // @[Mux.scala 46:16:@11928.4]
  assign _T_12812 = 5'h13 == _T_11317_28; // @[Mux.scala 46:19:@11929.4]
  assign _T_12813 = _T_12812 ? _T_10366_18 : _T_12811; // @[Mux.scala 46:16:@11930.4]
  assign _T_12814 = 5'h12 == _T_11317_28; // @[Mux.scala 46:19:@11931.4]
  assign _T_12815 = _T_12814 ? _T_10366_17 : _T_12813; // @[Mux.scala 46:16:@11932.4]
  assign _T_12816 = 5'h11 == _T_11317_28; // @[Mux.scala 46:19:@11933.4]
  assign _T_12817 = _T_12816 ? _T_10366_16 : _T_12815; // @[Mux.scala 46:16:@11934.4]
  assign _T_12818 = 5'h10 == _T_11317_28; // @[Mux.scala 46:19:@11935.4]
  assign _T_12819 = _T_12818 ? _T_10366_15 : _T_12817; // @[Mux.scala 46:16:@11936.4]
  assign _T_12820 = 5'hf == _T_11317_28; // @[Mux.scala 46:19:@11937.4]
  assign _T_12821 = _T_12820 ? _T_10366_14 : _T_12819; // @[Mux.scala 46:16:@11938.4]
  assign _T_12822 = 5'he == _T_11317_28; // @[Mux.scala 46:19:@11939.4]
  assign _T_12823 = _T_12822 ? _T_10366_13 : _T_12821; // @[Mux.scala 46:16:@11940.4]
  assign _T_12824 = 5'hd == _T_11317_28; // @[Mux.scala 46:19:@11941.4]
  assign _T_12825 = _T_12824 ? _T_10366_12 : _T_12823; // @[Mux.scala 46:16:@11942.4]
  assign _T_12826 = 5'hc == _T_11317_28; // @[Mux.scala 46:19:@11943.4]
  assign _T_12827 = _T_12826 ? _T_10366_11 : _T_12825; // @[Mux.scala 46:16:@11944.4]
  assign _T_12828 = 5'hb == _T_11317_28; // @[Mux.scala 46:19:@11945.4]
  assign _T_12829 = _T_12828 ? _T_10366_10 : _T_12827; // @[Mux.scala 46:16:@11946.4]
  assign _T_12830 = 5'ha == _T_11317_28; // @[Mux.scala 46:19:@11947.4]
  assign _T_12831 = _T_12830 ? _T_10366_9 : _T_12829; // @[Mux.scala 46:16:@11948.4]
  assign _T_12832 = 5'h9 == _T_11317_28; // @[Mux.scala 46:19:@11949.4]
  assign _T_12833 = _T_12832 ? _T_10366_8 : _T_12831; // @[Mux.scala 46:16:@11950.4]
  assign _T_12834 = 5'h8 == _T_11317_28; // @[Mux.scala 46:19:@11951.4]
  assign _T_12835 = _T_12834 ? _T_10366_7 : _T_12833; // @[Mux.scala 46:16:@11952.4]
  assign _T_12836 = 5'h7 == _T_11317_28; // @[Mux.scala 46:19:@11953.4]
  assign _T_12837 = _T_12836 ? _T_10366_6 : _T_12835; // @[Mux.scala 46:16:@11954.4]
  assign _T_12838 = 5'h6 == _T_11317_28; // @[Mux.scala 46:19:@11955.4]
  assign _T_12839 = _T_12838 ? _T_10366_5 : _T_12837; // @[Mux.scala 46:16:@11956.4]
  assign _T_12840 = 5'h5 == _T_11317_28; // @[Mux.scala 46:19:@11957.4]
  assign _T_12841 = _T_12840 ? _T_10366_4 : _T_12839; // @[Mux.scala 46:16:@11958.4]
  assign _T_12842 = 5'h4 == _T_11317_28; // @[Mux.scala 46:19:@11959.4]
  assign _T_12843 = _T_12842 ? _T_10366_3 : _T_12841; // @[Mux.scala 46:16:@11960.4]
  assign _T_12844 = 5'h3 == _T_11317_28; // @[Mux.scala 46:19:@11961.4]
  assign _T_12845 = _T_12844 ? _T_10366_2 : _T_12843; // @[Mux.scala 46:16:@11962.4]
  assign _T_12846 = 5'h2 == _T_11317_28; // @[Mux.scala 46:19:@11963.4]
  assign _T_12847 = _T_12846 ? _T_10366_1 : _T_12845; // @[Mux.scala 46:16:@11964.4]
  assign _T_12848 = 5'h1 == _T_11317_28; // @[Mux.scala 46:19:@11965.4]
  assign _T_12849 = _T_12848 ? _T_10366_0 : _T_12847; // @[Mux.scala 46:16:@11966.4]
  assign _T_12881 = 5'h1e == _T_11317_29; // @[Mux.scala 46:19:@11968.4]
  assign _T_12882 = _T_12881 ? _T_10366_29 : 8'h0; // @[Mux.scala 46:16:@11969.4]
  assign _T_12883 = 5'h1d == _T_11317_29; // @[Mux.scala 46:19:@11970.4]
  assign _T_12884 = _T_12883 ? _T_10366_28 : _T_12882; // @[Mux.scala 46:16:@11971.4]
  assign _T_12885 = 5'h1c == _T_11317_29; // @[Mux.scala 46:19:@11972.4]
  assign _T_12886 = _T_12885 ? _T_10366_27 : _T_12884; // @[Mux.scala 46:16:@11973.4]
  assign _T_12887 = 5'h1b == _T_11317_29; // @[Mux.scala 46:19:@11974.4]
  assign _T_12888 = _T_12887 ? _T_10366_26 : _T_12886; // @[Mux.scala 46:16:@11975.4]
  assign _T_12889 = 5'h1a == _T_11317_29; // @[Mux.scala 46:19:@11976.4]
  assign _T_12890 = _T_12889 ? _T_10366_25 : _T_12888; // @[Mux.scala 46:16:@11977.4]
  assign _T_12891 = 5'h19 == _T_11317_29; // @[Mux.scala 46:19:@11978.4]
  assign _T_12892 = _T_12891 ? _T_10366_24 : _T_12890; // @[Mux.scala 46:16:@11979.4]
  assign _T_12893 = 5'h18 == _T_11317_29; // @[Mux.scala 46:19:@11980.4]
  assign _T_12894 = _T_12893 ? _T_10366_23 : _T_12892; // @[Mux.scala 46:16:@11981.4]
  assign _T_12895 = 5'h17 == _T_11317_29; // @[Mux.scala 46:19:@11982.4]
  assign _T_12896 = _T_12895 ? _T_10366_22 : _T_12894; // @[Mux.scala 46:16:@11983.4]
  assign _T_12897 = 5'h16 == _T_11317_29; // @[Mux.scala 46:19:@11984.4]
  assign _T_12898 = _T_12897 ? _T_10366_21 : _T_12896; // @[Mux.scala 46:16:@11985.4]
  assign _T_12899 = 5'h15 == _T_11317_29; // @[Mux.scala 46:19:@11986.4]
  assign _T_12900 = _T_12899 ? _T_10366_20 : _T_12898; // @[Mux.scala 46:16:@11987.4]
  assign _T_12901 = 5'h14 == _T_11317_29; // @[Mux.scala 46:19:@11988.4]
  assign _T_12902 = _T_12901 ? _T_10366_19 : _T_12900; // @[Mux.scala 46:16:@11989.4]
  assign _T_12903 = 5'h13 == _T_11317_29; // @[Mux.scala 46:19:@11990.4]
  assign _T_12904 = _T_12903 ? _T_10366_18 : _T_12902; // @[Mux.scala 46:16:@11991.4]
  assign _T_12905 = 5'h12 == _T_11317_29; // @[Mux.scala 46:19:@11992.4]
  assign _T_12906 = _T_12905 ? _T_10366_17 : _T_12904; // @[Mux.scala 46:16:@11993.4]
  assign _T_12907 = 5'h11 == _T_11317_29; // @[Mux.scala 46:19:@11994.4]
  assign _T_12908 = _T_12907 ? _T_10366_16 : _T_12906; // @[Mux.scala 46:16:@11995.4]
  assign _T_12909 = 5'h10 == _T_11317_29; // @[Mux.scala 46:19:@11996.4]
  assign _T_12910 = _T_12909 ? _T_10366_15 : _T_12908; // @[Mux.scala 46:16:@11997.4]
  assign _T_12911 = 5'hf == _T_11317_29; // @[Mux.scala 46:19:@11998.4]
  assign _T_12912 = _T_12911 ? _T_10366_14 : _T_12910; // @[Mux.scala 46:16:@11999.4]
  assign _T_12913 = 5'he == _T_11317_29; // @[Mux.scala 46:19:@12000.4]
  assign _T_12914 = _T_12913 ? _T_10366_13 : _T_12912; // @[Mux.scala 46:16:@12001.4]
  assign _T_12915 = 5'hd == _T_11317_29; // @[Mux.scala 46:19:@12002.4]
  assign _T_12916 = _T_12915 ? _T_10366_12 : _T_12914; // @[Mux.scala 46:16:@12003.4]
  assign _T_12917 = 5'hc == _T_11317_29; // @[Mux.scala 46:19:@12004.4]
  assign _T_12918 = _T_12917 ? _T_10366_11 : _T_12916; // @[Mux.scala 46:16:@12005.4]
  assign _T_12919 = 5'hb == _T_11317_29; // @[Mux.scala 46:19:@12006.4]
  assign _T_12920 = _T_12919 ? _T_10366_10 : _T_12918; // @[Mux.scala 46:16:@12007.4]
  assign _T_12921 = 5'ha == _T_11317_29; // @[Mux.scala 46:19:@12008.4]
  assign _T_12922 = _T_12921 ? _T_10366_9 : _T_12920; // @[Mux.scala 46:16:@12009.4]
  assign _T_12923 = 5'h9 == _T_11317_29; // @[Mux.scala 46:19:@12010.4]
  assign _T_12924 = _T_12923 ? _T_10366_8 : _T_12922; // @[Mux.scala 46:16:@12011.4]
  assign _T_12925 = 5'h8 == _T_11317_29; // @[Mux.scala 46:19:@12012.4]
  assign _T_12926 = _T_12925 ? _T_10366_7 : _T_12924; // @[Mux.scala 46:16:@12013.4]
  assign _T_12927 = 5'h7 == _T_11317_29; // @[Mux.scala 46:19:@12014.4]
  assign _T_12928 = _T_12927 ? _T_10366_6 : _T_12926; // @[Mux.scala 46:16:@12015.4]
  assign _T_12929 = 5'h6 == _T_11317_29; // @[Mux.scala 46:19:@12016.4]
  assign _T_12930 = _T_12929 ? _T_10366_5 : _T_12928; // @[Mux.scala 46:16:@12017.4]
  assign _T_12931 = 5'h5 == _T_11317_29; // @[Mux.scala 46:19:@12018.4]
  assign _T_12932 = _T_12931 ? _T_10366_4 : _T_12930; // @[Mux.scala 46:16:@12019.4]
  assign _T_12933 = 5'h4 == _T_11317_29; // @[Mux.scala 46:19:@12020.4]
  assign _T_12934 = _T_12933 ? _T_10366_3 : _T_12932; // @[Mux.scala 46:16:@12021.4]
  assign _T_12935 = 5'h3 == _T_11317_29; // @[Mux.scala 46:19:@12022.4]
  assign _T_12936 = _T_12935 ? _T_10366_2 : _T_12934; // @[Mux.scala 46:16:@12023.4]
  assign _T_12937 = 5'h2 == _T_11317_29; // @[Mux.scala 46:19:@12024.4]
  assign _T_12938 = _T_12937 ? _T_10366_1 : _T_12936; // @[Mux.scala 46:16:@12025.4]
  assign _T_12939 = 5'h1 == _T_11317_29; // @[Mux.scala 46:19:@12026.4]
  assign _T_12940 = _T_12939 ? _T_10366_0 : _T_12938; // @[Mux.scala 46:16:@12027.4]
  assign _T_12973 = 5'h1f == _T_11317_30; // @[Mux.scala 46:19:@12029.4]
  assign _T_12974 = _T_12973 ? _T_10366_30 : 8'h0; // @[Mux.scala 46:16:@12030.4]
  assign _T_12975 = 5'h1e == _T_11317_30; // @[Mux.scala 46:19:@12031.4]
  assign _T_12976 = _T_12975 ? _T_10366_29 : _T_12974; // @[Mux.scala 46:16:@12032.4]
  assign _T_12977 = 5'h1d == _T_11317_30; // @[Mux.scala 46:19:@12033.4]
  assign _T_12978 = _T_12977 ? _T_10366_28 : _T_12976; // @[Mux.scala 46:16:@12034.4]
  assign _T_12979 = 5'h1c == _T_11317_30; // @[Mux.scala 46:19:@12035.4]
  assign _T_12980 = _T_12979 ? _T_10366_27 : _T_12978; // @[Mux.scala 46:16:@12036.4]
  assign _T_12981 = 5'h1b == _T_11317_30; // @[Mux.scala 46:19:@12037.4]
  assign _T_12982 = _T_12981 ? _T_10366_26 : _T_12980; // @[Mux.scala 46:16:@12038.4]
  assign _T_12983 = 5'h1a == _T_11317_30; // @[Mux.scala 46:19:@12039.4]
  assign _T_12984 = _T_12983 ? _T_10366_25 : _T_12982; // @[Mux.scala 46:16:@12040.4]
  assign _T_12985 = 5'h19 == _T_11317_30; // @[Mux.scala 46:19:@12041.4]
  assign _T_12986 = _T_12985 ? _T_10366_24 : _T_12984; // @[Mux.scala 46:16:@12042.4]
  assign _T_12987 = 5'h18 == _T_11317_30; // @[Mux.scala 46:19:@12043.4]
  assign _T_12988 = _T_12987 ? _T_10366_23 : _T_12986; // @[Mux.scala 46:16:@12044.4]
  assign _T_12989 = 5'h17 == _T_11317_30; // @[Mux.scala 46:19:@12045.4]
  assign _T_12990 = _T_12989 ? _T_10366_22 : _T_12988; // @[Mux.scala 46:16:@12046.4]
  assign _T_12991 = 5'h16 == _T_11317_30; // @[Mux.scala 46:19:@12047.4]
  assign _T_12992 = _T_12991 ? _T_10366_21 : _T_12990; // @[Mux.scala 46:16:@12048.4]
  assign _T_12993 = 5'h15 == _T_11317_30; // @[Mux.scala 46:19:@12049.4]
  assign _T_12994 = _T_12993 ? _T_10366_20 : _T_12992; // @[Mux.scala 46:16:@12050.4]
  assign _T_12995 = 5'h14 == _T_11317_30; // @[Mux.scala 46:19:@12051.4]
  assign _T_12996 = _T_12995 ? _T_10366_19 : _T_12994; // @[Mux.scala 46:16:@12052.4]
  assign _T_12997 = 5'h13 == _T_11317_30; // @[Mux.scala 46:19:@12053.4]
  assign _T_12998 = _T_12997 ? _T_10366_18 : _T_12996; // @[Mux.scala 46:16:@12054.4]
  assign _T_12999 = 5'h12 == _T_11317_30; // @[Mux.scala 46:19:@12055.4]
  assign _T_13000 = _T_12999 ? _T_10366_17 : _T_12998; // @[Mux.scala 46:16:@12056.4]
  assign _T_13001 = 5'h11 == _T_11317_30; // @[Mux.scala 46:19:@12057.4]
  assign _T_13002 = _T_13001 ? _T_10366_16 : _T_13000; // @[Mux.scala 46:16:@12058.4]
  assign _T_13003 = 5'h10 == _T_11317_30; // @[Mux.scala 46:19:@12059.4]
  assign _T_13004 = _T_13003 ? _T_10366_15 : _T_13002; // @[Mux.scala 46:16:@12060.4]
  assign _T_13005 = 5'hf == _T_11317_30; // @[Mux.scala 46:19:@12061.4]
  assign _T_13006 = _T_13005 ? _T_10366_14 : _T_13004; // @[Mux.scala 46:16:@12062.4]
  assign _T_13007 = 5'he == _T_11317_30; // @[Mux.scala 46:19:@12063.4]
  assign _T_13008 = _T_13007 ? _T_10366_13 : _T_13006; // @[Mux.scala 46:16:@12064.4]
  assign _T_13009 = 5'hd == _T_11317_30; // @[Mux.scala 46:19:@12065.4]
  assign _T_13010 = _T_13009 ? _T_10366_12 : _T_13008; // @[Mux.scala 46:16:@12066.4]
  assign _T_13011 = 5'hc == _T_11317_30; // @[Mux.scala 46:19:@12067.4]
  assign _T_13012 = _T_13011 ? _T_10366_11 : _T_13010; // @[Mux.scala 46:16:@12068.4]
  assign _T_13013 = 5'hb == _T_11317_30; // @[Mux.scala 46:19:@12069.4]
  assign _T_13014 = _T_13013 ? _T_10366_10 : _T_13012; // @[Mux.scala 46:16:@12070.4]
  assign _T_13015 = 5'ha == _T_11317_30; // @[Mux.scala 46:19:@12071.4]
  assign _T_13016 = _T_13015 ? _T_10366_9 : _T_13014; // @[Mux.scala 46:16:@12072.4]
  assign _T_13017 = 5'h9 == _T_11317_30; // @[Mux.scala 46:19:@12073.4]
  assign _T_13018 = _T_13017 ? _T_10366_8 : _T_13016; // @[Mux.scala 46:16:@12074.4]
  assign _T_13019 = 5'h8 == _T_11317_30; // @[Mux.scala 46:19:@12075.4]
  assign _T_13020 = _T_13019 ? _T_10366_7 : _T_13018; // @[Mux.scala 46:16:@12076.4]
  assign _T_13021 = 5'h7 == _T_11317_30; // @[Mux.scala 46:19:@12077.4]
  assign _T_13022 = _T_13021 ? _T_10366_6 : _T_13020; // @[Mux.scala 46:16:@12078.4]
  assign _T_13023 = 5'h6 == _T_11317_30; // @[Mux.scala 46:19:@12079.4]
  assign _T_13024 = _T_13023 ? _T_10366_5 : _T_13022; // @[Mux.scala 46:16:@12080.4]
  assign _T_13025 = 5'h5 == _T_11317_30; // @[Mux.scala 46:19:@12081.4]
  assign _T_13026 = _T_13025 ? _T_10366_4 : _T_13024; // @[Mux.scala 46:16:@12082.4]
  assign _T_13027 = 5'h4 == _T_11317_30; // @[Mux.scala 46:19:@12083.4]
  assign _T_13028 = _T_13027 ? _T_10366_3 : _T_13026; // @[Mux.scala 46:16:@12084.4]
  assign _T_13029 = 5'h3 == _T_11317_30; // @[Mux.scala 46:19:@12085.4]
  assign _T_13030 = _T_13029 ? _T_10366_2 : _T_13028; // @[Mux.scala 46:16:@12086.4]
  assign _T_13031 = 5'h2 == _T_11317_30; // @[Mux.scala 46:19:@12087.4]
  assign _T_13032 = _T_13031 ? _T_10366_1 : _T_13030; // @[Mux.scala 46:16:@12088.4]
  assign _T_13033 = 5'h1 == _T_11317_30; // @[Mux.scala 46:19:@12089.4]
  assign _T_13034 = _T_13033 ? _T_10366_0 : _T_13032; // @[Mux.scala 46:16:@12090.4]
  assign _T_13068 = 6'h20 == _T_11317_31; // @[Mux.scala 46:19:@12092.4]
  assign _T_13069 = _T_13068 ? _T_10366_31 : 8'h0; // @[Mux.scala 46:16:@12093.4]
  assign _T_13070 = 6'h1f == _T_11317_31; // @[Mux.scala 46:19:@12094.4]
  assign _T_13071 = _T_13070 ? _T_10366_30 : _T_13069; // @[Mux.scala 46:16:@12095.4]
  assign _T_13072 = 6'h1e == _T_11317_31; // @[Mux.scala 46:19:@12096.4]
  assign _T_13073 = _T_13072 ? _T_10366_29 : _T_13071; // @[Mux.scala 46:16:@12097.4]
  assign _T_13074 = 6'h1d == _T_11317_31; // @[Mux.scala 46:19:@12098.4]
  assign _T_13075 = _T_13074 ? _T_10366_28 : _T_13073; // @[Mux.scala 46:16:@12099.4]
  assign _T_13076 = 6'h1c == _T_11317_31; // @[Mux.scala 46:19:@12100.4]
  assign _T_13077 = _T_13076 ? _T_10366_27 : _T_13075; // @[Mux.scala 46:16:@12101.4]
  assign _T_13078 = 6'h1b == _T_11317_31; // @[Mux.scala 46:19:@12102.4]
  assign _T_13079 = _T_13078 ? _T_10366_26 : _T_13077; // @[Mux.scala 46:16:@12103.4]
  assign _T_13080 = 6'h1a == _T_11317_31; // @[Mux.scala 46:19:@12104.4]
  assign _T_13081 = _T_13080 ? _T_10366_25 : _T_13079; // @[Mux.scala 46:16:@12105.4]
  assign _T_13082 = 6'h19 == _T_11317_31; // @[Mux.scala 46:19:@12106.4]
  assign _T_13083 = _T_13082 ? _T_10366_24 : _T_13081; // @[Mux.scala 46:16:@12107.4]
  assign _T_13084 = 6'h18 == _T_11317_31; // @[Mux.scala 46:19:@12108.4]
  assign _T_13085 = _T_13084 ? _T_10366_23 : _T_13083; // @[Mux.scala 46:16:@12109.4]
  assign _T_13086 = 6'h17 == _T_11317_31; // @[Mux.scala 46:19:@12110.4]
  assign _T_13087 = _T_13086 ? _T_10366_22 : _T_13085; // @[Mux.scala 46:16:@12111.4]
  assign _T_13088 = 6'h16 == _T_11317_31; // @[Mux.scala 46:19:@12112.4]
  assign _T_13089 = _T_13088 ? _T_10366_21 : _T_13087; // @[Mux.scala 46:16:@12113.4]
  assign _T_13090 = 6'h15 == _T_11317_31; // @[Mux.scala 46:19:@12114.4]
  assign _T_13091 = _T_13090 ? _T_10366_20 : _T_13089; // @[Mux.scala 46:16:@12115.4]
  assign _T_13092 = 6'h14 == _T_11317_31; // @[Mux.scala 46:19:@12116.4]
  assign _T_13093 = _T_13092 ? _T_10366_19 : _T_13091; // @[Mux.scala 46:16:@12117.4]
  assign _T_13094 = 6'h13 == _T_11317_31; // @[Mux.scala 46:19:@12118.4]
  assign _T_13095 = _T_13094 ? _T_10366_18 : _T_13093; // @[Mux.scala 46:16:@12119.4]
  assign _T_13096 = 6'h12 == _T_11317_31; // @[Mux.scala 46:19:@12120.4]
  assign _T_13097 = _T_13096 ? _T_10366_17 : _T_13095; // @[Mux.scala 46:16:@12121.4]
  assign _T_13098 = 6'h11 == _T_11317_31; // @[Mux.scala 46:19:@12122.4]
  assign _T_13099 = _T_13098 ? _T_10366_16 : _T_13097; // @[Mux.scala 46:16:@12123.4]
  assign _T_13100 = 6'h10 == _T_11317_31; // @[Mux.scala 46:19:@12124.4]
  assign _T_13101 = _T_13100 ? _T_10366_15 : _T_13099; // @[Mux.scala 46:16:@12125.4]
  assign _T_13102 = 6'hf == _T_11317_31; // @[Mux.scala 46:19:@12126.4]
  assign _T_13103 = _T_13102 ? _T_10366_14 : _T_13101; // @[Mux.scala 46:16:@12127.4]
  assign _T_13104 = 6'he == _T_11317_31; // @[Mux.scala 46:19:@12128.4]
  assign _T_13105 = _T_13104 ? _T_10366_13 : _T_13103; // @[Mux.scala 46:16:@12129.4]
  assign _T_13106 = 6'hd == _T_11317_31; // @[Mux.scala 46:19:@12130.4]
  assign _T_13107 = _T_13106 ? _T_10366_12 : _T_13105; // @[Mux.scala 46:16:@12131.4]
  assign _T_13108 = 6'hc == _T_11317_31; // @[Mux.scala 46:19:@12132.4]
  assign _T_13109 = _T_13108 ? _T_10366_11 : _T_13107; // @[Mux.scala 46:16:@12133.4]
  assign _T_13110 = 6'hb == _T_11317_31; // @[Mux.scala 46:19:@12134.4]
  assign _T_13111 = _T_13110 ? _T_10366_10 : _T_13109; // @[Mux.scala 46:16:@12135.4]
  assign _T_13112 = 6'ha == _T_11317_31; // @[Mux.scala 46:19:@12136.4]
  assign _T_13113 = _T_13112 ? _T_10366_9 : _T_13111; // @[Mux.scala 46:16:@12137.4]
  assign _T_13114 = 6'h9 == _T_11317_31; // @[Mux.scala 46:19:@12138.4]
  assign _T_13115 = _T_13114 ? _T_10366_8 : _T_13113; // @[Mux.scala 46:16:@12139.4]
  assign _T_13116 = 6'h8 == _T_11317_31; // @[Mux.scala 46:19:@12140.4]
  assign _T_13117 = _T_13116 ? _T_10366_7 : _T_13115; // @[Mux.scala 46:16:@12141.4]
  assign _T_13118 = 6'h7 == _T_11317_31; // @[Mux.scala 46:19:@12142.4]
  assign _T_13119 = _T_13118 ? _T_10366_6 : _T_13117; // @[Mux.scala 46:16:@12143.4]
  assign _T_13120 = 6'h6 == _T_11317_31; // @[Mux.scala 46:19:@12144.4]
  assign _T_13121 = _T_13120 ? _T_10366_5 : _T_13119; // @[Mux.scala 46:16:@12145.4]
  assign _T_13122 = 6'h5 == _T_11317_31; // @[Mux.scala 46:19:@12146.4]
  assign _T_13123 = _T_13122 ? _T_10366_4 : _T_13121; // @[Mux.scala 46:16:@12147.4]
  assign _T_13124 = 6'h4 == _T_11317_31; // @[Mux.scala 46:19:@12148.4]
  assign _T_13125 = _T_13124 ? _T_10366_3 : _T_13123; // @[Mux.scala 46:16:@12149.4]
  assign _T_13126 = 6'h3 == _T_11317_31; // @[Mux.scala 46:19:@12150.4]
  assign _T_13127 = _T_13126 ? _T_10366_2 : _T_13125; // @[Mux.scala 46:16:@12151.4]
  assign _T_13128 = 6'h2 == _T_11317_31; // @[Mux.scala 46:19:@12152.4]
  assign _T_13129 = _T_13128 ? _T_10366_1 : _T_13127; // @[Mux.scala 46:16:@12153.4]
  assign _T_13130 = 6'h1 == _T_11317_31; // @[Mux.scala 46:19:@12154.4]
  assign _T_13131 = _T_13130 ? _T_10366_0 : _T_13129; // @[Mux.scala 46:16:@12155.4]
  assign _T_13166 = 6'h21 == _T_11317_32; // @[Mux.scala 46:19:@12157.4]
  assign _T_13167 = _T_13166 ? _T_10366_32 : 8'h0; // @[Mux.scala 46:16:@12158.4]
  assign _T_13168 = 6'h20 == _T_11317_32; // @[Mux.scala 46:19:@12159.4]
  assign _T_13169 = _T_13168 ? _T_10366_31 : _T_13167; // @[Mux.scala 46:16:@12160.4]
  assign _T_13170 = 6'h1f == _T_11317_32; // @[Mux.scala 46:19:@12161.4]
  assign _T_13171 = _T_13170 ? _T_10366_30 : _T_13169; // @[Mux.scala 46:16:@12162.4]
  assign _T_13172 = 6'h1e == _T_11317_32; // @[Mux.scala 46:19:@12163.4]
  assign _T_13173 = _T_13172 ? _T_10366_29 : _T_13171; // @[Mux.scala 46:16:@12164.4]
  assign _T_13174 = 6'h1d == _T_11317_32; // @[Mux.scala 46:19:@12165.4]
  assign _T_13175 = _T_13174 ? _T_10366_28 : _T_13173; // @[Mux.scala 46:16:@12166.4]
  assign _T_13176 = 6'h1c == _T_11317_32; // @[Mux.scala 46:19:@12167.4]
  assign _T_13177 = _T_13176 ? _T_10366_27 : _T_13175; // @[Mux.scala 46:16:@12168.4]
  assign _T_13178 = 6'h1b == _T_11317_32; // @[Mux.scala 46:19:@12169.4]
  assign _T_13179 = _T_13178 ? _T_10366_26 : _T_13177; // @[Mux.scala 46:16:@12170.4]
  assign _T_13180 = 6'h1a == _T_11317_32; // @[Mux.scala 46:19:@12171.4]
  assign _T_13181 = _T_13180 ? _T_10366_25 : _T_13179; // @[Mux.scala 46:16:@12172.4]
  assign _T_13182 = 6'h19 == _T_11317_32; // @[Mux.scala 46:19:@12173.4]
  assign _T_13183 = _T_13182 ? _T_10366_24 : _T_13181; // @[Mux.scala 46:16:@12174.4]
  assign _T_13184 = 6'h18 == _T_11317_32; // @[Mux.scala 46:19:@12175.4]
  assign _T_13185 = _T_13184 ? _T_10366_23 : _T_13183; // @[Mux.scala 46:16:@12176.4]
  assign _T_13186 = 6'h17 == _T_11317_32; // @[Mux.scala 46:19:@12177.4]
  assign _T_13187 = _T_13186 ? _T_10366_22 : _T_13185; // @[Mux.scala 46:16:@12178.4]
  assign _T_13188 = 6'h16 == _T_11317_32; // @[Mux.scala 46:19:@12179.4]
  assign _T_13189 = _T_13188 ? _T_10366_21 : _T_13187; // @[Mux.scala 46:16:@12180.4]
  assign _T_13190 = 6'h15 == _T_11317_32; // @[Mux.scala 46:19:@12181.4]
  assign _T_13191 = _T_13190 ? _T_10366_20 : _T_13189; // @[Mux.scala 46:16:@12182.4]
  assign _T_13192 = 6'h14 == _T_11317_32; // @[Mux.scala 46:19:@12183.4]
  assign _T_13193 = _T_13192 ? _T_10366_19 : _T_13191; // @[Mux.scala 46:16:@12184.4]
  assign _T_13194 = 6'h13 == _T_11317_32; // @[Mux.scala 46:19:@12185.4]
  assign _T_13195 = _T_13194 ? _T_10366_18 : _T_13193; // @[Mux.scala 46:16:@12186.4]
  assign _T_13196 = 6'h12 == _T_11317_32; // @[Mux.scala 46:19:@12187.4]
  assign _T_13197 = _T_13196 ? _T_10366_17 : _T_13195; // @[Mux.scala 46:16:@12188.4]
  assign _T_13198 = 6'h11 == _T_11317_32; // @[Mux.scala 46:19:@12189.4]
  assign _T_13199 = _T_13198 ? _T_10366_16 : _T_13197; // @[Mux.scala 46:16:@12190.4]
  assign _T_13200 = 6'h10 == _T_11317_32; // @[Mux.scala 46:19:@12191.4]
  assign _T_13201 = _T_13200 ? _T_10366_15 : _T_13199; // @[Mux.scala 46:16:@12192.4]
  assign _T_13202 = 6'hf == _T_11317_32; // @[Mux.scala 46:19:@12193.4]
  assign _T_13203 = _T_13202 ? _T_10366_14 : _T_13201; // @[Mux.scala 46:16:@12194.4]
  assign _T_13204 = 6'he == _T_11317_32; // @[Mux.scala 46:19:@12195.4]
  assign _T_13205 = _T_13204 ? _T_10366_13 : _T_13203; // @[Mux.scala 46:16:@12196.4]
  assign _T_13206 = 6'hd == _T_11317_32; // @[Mux.scala 46:19:@12197.4]
  assign _T_13207 = _T_13206 ? _T_10366_12 : _T_13205; // @[Mux.scala 46:16:@12198.4]
  assign _T_13208 = 6'hc == _T_11317_32; // @[Mux.scala 46:19:@12199.4]
  assign _T_13209 = _T_13208 ? _T_10366_11 : _T_13207; // @[Mux.scala 46:16:@12200.4]
  assign _T_13210 = 6'hb == _T_11317_32; // @[Mux.scala 46:19:@12201.4]
  assign _T_13211 = _T_13210 ? _T_10366_10 : _T_13209; // @[Mux.scala 46:16:@12202.4]
  assign _T_13212 = 6'ha == _T_11317_32; // @[Mux.scala 46:19:@12203.4]
  assign _T_13213 = _T_13212 ? _T_10366_9 : _T_13211; // @[Mux.scala 46:16:@12204.4]
  assign _T_13214 = 6'h9 == _T_11317_32; // @[Mux.scala 46:19:@12205.4]
  assign _T_13215 = _T_13214 ? _T_10366_8 : _T_13213; // @[Mux.scala 46:16:@12206.4]
  assign _T_13216 = 6'h8 == _T_11317_32; // @[Mux.scala 46:19:@12207.4]
  assign _T_13217 = _T_13216 ? _T_10366_7 : _T_13215; // @[Mux.scala 46:16:@12208.4]
  assign _T_13218 = 6'h7 == _T_11317_32; // @[Mux.scala 46:19:@12209.4]
  assign _T_13219 = _T_13218 ? _T_10366_6 : _T_13217; // @[Mux.scala 46:16:@12210.4]
  assign _T_13220 = 6'h6 == _T_11317_32; // @[Mux.scala 46:19:@12211.4]
  assign _T_13221 = _T_13220 ? _T_10366_5 : _T_13219; // @[Mux.scala 46:16:@12212.4]
  assign _T_13222 = 6'h5 == _T_11317_32; // @[Mux.scala 46:19:@12213.4]
  assign _T_13223 = _T_13222 ? _T_10366_4 : _T_13221; // @[Mux.scala 46:16:@12214.4]
  assign _T_13224 = 6'h4 == _T_11317_32; // @[Mux.scala 46:19:@12215.4]
  assign _T_13225 = _T_13224 ? _T_10366_3 : _T_13223; // @[Mux.scala 46:16:@12216.4]
  assign _T_13226 = 6'h3 == _T_11317_32; // @[Mux.scala 46:19:@12217.4]
  assign _T_13227 = _T_13226 ? _T_10366_2 : _T_13225; // @[Mux.scala 46:16:@12218.4]
  assign _T_13228 = 6'h2 == _T_11317_32; // @[Mux.scala 46:19:@12219.4]
  assign _T_13229 = _T_13228 ? _T_10366_1 : _T_13227; // @[Mux.scala 46:16:@12220.4]
  assign _T_13230 = 6'h1 == _T_11317_32; // @[Mux.scala 46:19:@12221.4]
  assign _T_13231 = _T_13230 ? _T_10366_0 : _T_13229; // @[Mux.scala 46:16:@12222.4]
  assign _T_13267 = 6'h22 == _T_11317_33; // @[Mux.scala 46:19:@12224.4]
  assign _T_13268 = _T_13267 ? _T_10366_33 : 8'h0; // @[Mux.scala 46:16:@12225.4]
  assign _T_13269 = 6'h21 == _T_11317_33; // @[Mux.scala 46:19:@12226.4]
  assign _T_13270 = _T_13269 ? _T_10366_32 : _T_13268; // @[Mux.scala 46:16:@12227.4]
  assign _T_13271 = 6'h20 == _T_11317_33; // @[Mux.scala 46:19:@12228.4]
  assign _T_13272 = _T_13271 ? _T_10366_31 : _T_13270; // @[Mux.scala 46:16:@12229.4]
  assign _T_13273 = 6'h1f == _T_11317_33; // @[Mux.scala 46:19:@12230.4]
  assign _T_13274 = _T_13273 ? _T_10366_30 : _T_13272; // @[Mux.scala 46:16:@12231.4]
  assign _T_13275 = 6'h1e == _T_11317_33; // @[Mux.scala 46:19:@12232.4]
  assign _T_13276 = _T_13275 ? _T_10366_29 : _T_13274; // @[Mux.scala 46:16:@12233.4]
  assign _T_13277 = 6'h1d == _T_11317_33; // @[Mux.scala 46:19:@12234.4]
  assign _T_13278 = _T_13277 ? _T_10366_28 : _T_13276; // @[Mux.scala 46:16:@12235.4]
  assign _T_13279 = 6'h1c == _T_11317_33; // @[Mux.scala 46:19:@12236.4]
  assign _T_13280 = _T_13279 ? _T_10366_27 : _T_13278; // @[Mux.scala 46:16:@12237.4]
  assign _T_13281 = 6'h1b == _T_11317_33; // @[Mux.scala 46:19:@12238.4]
  assign _T_13282 = _T_13281 ? _T_10366_26 : _T_13280; // @[Mux.scala 46:16:@12239.4]
  assign _T_13283 = 6'h1a == _T_11317_33; // @[Mux.scala 46:19:@12240.4]
  assign _T_13284 = _T_13283 ? _T_10366_25 : _T_13282; // @[Mux.scala 46:16:@12241.4]
  assign _T_13285 = 6'h19 == _T_11317_33; // @[Mux.scala 46:19:@12242.4]
  assign _T_13286 = _T_13285 ? _T_10366_24 : _T_13284; // @[Mux.scala 46:16:@12243.4]
  assign _T_13287 = 6'h18 == _T_11317_33; // @[Mux.scala 46:19:@12244.4]
  assign _T_13288 = _T_13287 ? _T_10366_23 : _T_13286; // @[Mux.scala 46:16:@12245.4]
  assign _T_13289 = 6'h17 == _T_11317_33; // @[Mux.scala 46:19:@12246.4]
  assign _T_13290 = _T_13289 ? _T_10366_22 : _T_13288; // @[Mux.scala 46:16:@12247.4]
  assign _T_13291 = 6'h16 == _T_11317_33; // @[Mux.scala 46:19:@12248.4]
  assign _T_13292 = _T_13291 ? _T_10366_21 : _T_13290; // @[Mux.scala 46:16:@12249.4]
  assign _T_13293 = 6'h15 == _T_11317_33; // @[Mux.scala 46:19:@12250.4]
  assign _T_13294 = _T_13293 ? _T_10366_20 : _T_13292; // @[Mux.scala 46:16:@12251.4]
  assign _T_13295 = 6'h14 == _T_11317_33; // @[Mux.scala 46:19:@12252.4]
  assign _T_13296 = _T_13295 ? _T_10366_19 : _T_13294; // @[Mux.scala 46:16:@12253.4]
  assign _T_13297 = 6'h13 == _T_11317_33; // @[Mux.scala 46:19:@12254.4]
  assign _T_13298 = _T_13297 ? _T_10366_18 : _T_13296; // @[Mux.scala 46:16:@12255.4]
  assign _T_13299 = 6'h12 == _T_11317_33; // @[Mux.scala 46:19:@12256.4]
  assign _T_13300 = _T_13299 ? _T_10366_17 : _T_13298; // @[Mux.scala 46:16:@12257.4]
  assign _T_13301 = 6'h11 == _T_11317_33; // @[Mux.scala 46:19:@12258.4]
  assign _T_13302 = _T_13301 ? _T_10366_16 : _T_13300; // @[Mux.scala 46:16:@12259.4]
  assign _T_13303 = 6'h10 == _T_11317_33; // @[Mux.scala 46:19:@12260.4]
  assign _T_13304 = _T_13303 ? _T_10366_15 : _T_13302; // @[Mux.scala 46:16:@12261.4]
  assign _T_13305 = 6'hf == _T_11317_33; // @[Mux.scala 46:19:@12262.4]
  assign _T_13306 = _T_13305 ? _T_10366_14 : _T_13304; // @[Mux.scala 46:16:@12263.4]
  assign _T_13307 = 6'he == _T_11317_33; // @[Mux.scala 46:19:@12264.4]
  assign _T_13308 = _T_13307 ? _T_10366_13 : _T_13306; // @[Mux.scala 46:16:@12265.4]
  assign _T_13309 = 6'hd == _T_11317_33; // @[Mux.scala 46:19:@12266.4]
  assign _T_13310 = _T_13309 ? _T_10366_12 : _T_13308; // @[Mux.scala 46:16:@12267.4]
  assign _T_13311 = 6'hc == _T_11317_33; // @[Mux.scala 46:19:@12268.4]
  assign _T_13312 = _T_13311 ? _T_10366_11 : _T_13310; // @[Mux.scala 46:16:@12269.4]
  assign _T_13313 = 6'hb == _T_11317_33; // @[Mux.scala 46:19:@12270.4]
  assign _T_13314 = _T_13313 ? _T_10366_10 : _T_13312; // @[Mux.scala 46:16:@12271.4]
  assign _T_13315 = 6'ha == _T_11317_33; // @[Mux.scala 46:19:@12272.4]
  assign _T_13316 = _T_13315 ? _T_10366_9 : _T_13314; // @[Mux.scala 46:16:@12273.4]
  assign _T_13317 = 6'h9 == _T_11317_33; // @[Mux.scala 46:19:@12274.4]
  assign _T_13318 = _T_13317 ? _T_10366_8 : _T_13316; // @[Mux.scala 46:16:@12275.4]
  assign _T_13319 = 6'h8 == _T_11317_33; // @[Mux.scala 46:19:@12276.4]
  assign _T_13320 = _T_13319 ? _T_10366_7 : _T_13318; // @[Mux.scala 46:16:@12277.4]
  assign _T_13321 = 6'h7 == _T_11317_33; // @[Mux.scala 46:19:@12278.4]
  assign _T_13322 = _T_13321 ? _T_10366_6 : _T_13320; // @[Mux.scala 46:16:@12279.4]
  assign _T_13323 = 6'h6 == _T_11317_33; // @[Mux.scala 46:19:@12280.4]
  assign _T_13324 = _T_13323 ? _T_10366_5 : _T_13322; // @[Mux.scala 46:16:@12281.4]
  assign _T_13325 = 6'h5 == _T_11317_33; // @[Mux.scala 46:19:@12282.4]
  assign _T_13326 = _T_13325 ? _T_10366_4 : _T_13324; // @[Mux.scala 46:16:@12283.4]
  assign _T_13327 = 6'h4 == _T_11317_33; // @[Mux.scala 46:19:@12284.4]
  assign _T_13328 = _T_13327 ? _T_10366_3 : _T_13326; // @[Mux.scala 46:16:@12285.4]
  assign _T_13329 = 6'h3 == _T_11317_33; // @[Mux.scala 46:19:@12286.4]
  assign _T_13330 = _T_13329 ? _T_10366_2 : _T_13328; // @[Mux.scala 46:16:@12287.4]
  assign _T_13331 = 6'h2 == _T_11317_33; // @[Mux.scala 46:19:@12288.4]
  assign _T_13332 = _T_13331 ? _T_10366_1 : _T_13330; // @[Mux.scala 46:16:@12289.4]
  assign _T_13333 = 6'h1 == _T_11317_33; // @[Mux.scala 46:19:@12290.4]
  assign _T_13334 = _T_13333 ? _T_10366_0 : _T_13332; // @[Mux.scala 46:16:@12291.4]
  assign _T_13371 = 6'h23 == _T_11317_34; // @[Mux.scala 46:19:@12293.4]
  assign _T_13372 = _T_13371 ? _T_10366_34 : 8'h0; // @[Mux.scala 46:16:@12294.4]
  assign _T_13373 = 6'h22 == _T_11317_34; // @[Mux.scala 46:19:@12295.4]
  assign _T_13374 = _T_13373 ? _T_10366_33 : _T_13372; // @[Mux.scala 46:16:@12296.4]
  assign _T_13375 = 6'h21 == _T_11317_34; // @[Mux.scala 46:19:@12297.4]
  assign _T_13376 = _T_13375 ? _T_10366_32 : _T_13374; // @[Mux.scala 46:16:@12298.4]
  assign _T_13377 = 6'h20 == _T_11317_34; // @[Mux.scala 46:19:@12299.4]
  assign _T_13378 = _T_13377 ? _T_10366_31 : _T_13376; // @[Mux.scala 46:16:@12300.4]
  assign _T_13379 = 6'h1f == _T_11317_34; // @[Mux.scala 46:19:@12301.4]
  assign _T_13380 = _T_13379 ? _T_10366_30 : _T_13378; // @[Mux.scala 46:16:@12302.4]
  assign _T_13381 = 6'h1e == _T_11317_34; // @[Mux.scala 46:19:@12303.4]
  assign _T_13382 = _T_13381 ? _T_10366_29 : _T_13380; // @[Mux.scala 46:16:@12304.4]
  assign _T_13383 = 6'h1d == _T_11317_34; // @[Mux.scala 46:19:@12305.4]
  assign _T_13384 = _T_13383 ? _T_10366_28 : _T_13382; // @[Mux.scala 46:16:@12306.4]
  assign _T_13385 = 6'h1c == _T_11317_34; // @[Mux.scala 46:19:@12307.4]
  assign _T_13386 = _T_13385 ? _T_10366_27 : _T_13384; // @[Mux.scala 46:16:@12308.4]
  assign _T_13387 = 6'h1b == _T_11317_34; // @[Mux.scala 46:19:@12309.4]
  assign _T_13388 = _T_13387 ? _T_10366_26 : _T_13386; // @[Mux.scala 46:16:@12310.4]
  assign _T_13389 = 6'h1a == _T_11317_34; // @[Mux.scala 46:19:@12311.4]
  assign _T_13390 = _T_13389 ? _T_10366_25 : _T_13388; // @[Mux.scala 46:16:@12312.4]
  assign _T_13391 = 6'h19 == _T_11317_34; // @[Mux.scala 46:19:@12313.4]
  assign _T_13392 = _T_13391 ? _T_10366_24 : _T_13390; // @[Mux.scala 46:16:@12314.4]
  assign _T_13393 = 6'h18 == _T_11317_34; // @[Mux.scala 46:19:@12315.4]
  assign _T_13394 = _T_13393 ? _T_10366_23 : _T_13392; // @[Mux.scala 46:16:@12316.4]
  assign _T_13395 = 6'h17 == _T_11317_34; // @[Mux.scala 46:19:@12317.4]
  assign _T_13396 = _T_13395 ? _T_10366_22 : _T_13394; // @[Mux.scala 46:16:@12318.4]
  assign _T_13397 = 6'h16 == _T_11317_34; // @[Mux.scala 46:19:@12319.4]
  assign _T_13398 = _T_13397 ? _T_10366_21 : _T_13396; // @[Mux.scala 46:16:@12320.4]
  assign _T_13399 = 6'h15 == _T_11317_34; // @[Mux.scala 46:19:@12321.4]
  assign _T_13400 = _T_13399 ? _T_10366_20 : _T_13398; // @[Mux.scala 46:16:@12322.4]
  assign _T_13401 = 6'h14 == _T_11317_34; // @[Mux.scala 46:19:@12323.4]
  assign _T_13402 = _T_13401 ? _T_10366_19 : _T_13400; // @[Mux.scala 46:16:@12324.4]
  assign _T_13403 = 6'h13 == _T_11317_34; // @[Mux.scala 46:19:@12325.4]
  assign _T_13404 = _T_13403 ? _T_10366_18 : _T_13402; // @[Mux.scala 46:16:@12326.4]
  assign _T_13405 = 6'h12 == _T_11317_34; // @[Mux.scala 46:19:@12327.4]
  assign _T_13406 = _T_13405 ? _T_10366_17 : _T_13404; // @[Mux.scala 46:16:@12328.4]
  assign _T_13407 = 6'h11 == _T_11317_34; // @[Mux.scala 46:19:@12329.4]
  assign _T_13408 = _T_13407 ? _T_10366_16 : _T_13406; // @[Mux.scala 46:16:@12330.4]
  assign _T_13409 = 6'h10 == _T_11317_34; // @[Mux.scala 46:19:@12331.4]
  assign _T_13410 = _T_13409 ? _T_10366_15 : _T_13408; // @[Mux.scala 46:16:@12332.4]
  assign _T_13411 = 6'hf == _T_11317_34; // @[Mux.scala 46:19:@12333.4]
  assign _T_13412 = _T_13411 ? _T_10366_14 : _T_13410; // @[Mux.scala 46:16:@12334.4]
  assign _T_13413 = 6'he == _T_11317_34; // @[Mux.scala 46:19:@12335.4]
  assign _T_13414 = _T_13413 ? _T_10366_13 : _T_13412; // @[Mux.scala 46:16:@12336.4]
  assign _T_13415 = 6'hd == _T_11317_34; // @[Mux.scala 46:19:@12337.4]
  assign _T_13416 = _T_13415 ? _T_10366_12 : _T_13414; // @[Mux.scala 46:16:@12338.4]
  assign _T_13417 = 6'hc == _T_11317_34; // @[Mux.scala 46:19:@12339.4]
  assign _T_13418 = _T_13417 ? _T_10366_11 : _T_13416; // @[Mux.scala 46:16:@12340.4]
  assign _T_13419 = 6'hb == _T_11317_34; // @[Mux.scala 46:19:@12341.4]
  assign _T_13420 = _T_13419 ? _T_10366_10 : _T_13418; // @[Mux.scala 46:16:@12342.4]
  assign _T_13421 = 6'ha == _T_11317_34; // @[Mux.scala 46:19:@12343.4]
  assign _T_13422 = _T_13421 ? _T_10366_9 : _T_13420; // @[Mux.scala 46:16:@12344.4]
  assign _T_13423 = 6'h9 == _T_11317_34; // @[Mux.scala 46:19:@12345.4]
  assign _T_13424 = _T_13423 ? _T_10366_8 : _T_13422; // @[Mux.scala 46:16:@12346.4]
  assign _T_13425 = 6'h8 == _T_11317_34; // @[Mux.scala 46:19:@12347.4]
  assign _T_13426 = _T_13425 ? _T_10366_7 : _T_13424; // @[Mux.scala 46:16:@12348.4]
  assign _T_13427 = 6'h7 == _T_11317_34; // @[Mux.scala 46:19:@12349.4]
  assign _T_13428 = _T_13427 ? _T_10366_6 : _T_13426; // @[Mux.scala 46:16:@12350.4]
  assign _T_13429 = 6'h6 == _T_11317_34; // @[Mux.scala 46:19:@12351.4]
  assign _T_13430 = _T_13429 ? _T_10366_5 : _T_13428; // @[Mux.scala 46:16:@12352.4]
  assign _T_13431 = 6'h5 == _T_11317_34; // @[Mux.scala 46:19:@12353.4]
  assign _T_13432 = _T_13431 ? _T_10366_4 : _T_13430; // @[Mux.scala 46:16:@12354.4]
  assign _T_13433 = 6'h4 == _T_11317_34; // @[Mux.scala 46:19:@12355.4]
  assign _T_13434 = _T_13433 ? _T_10366_3 : _T_13432; // @[Mux.scala 46:16:@12356.4]
  assign _T_13435 = 6'h3 == _T_11317_34; // @[Mux.scala 46:19:@12357.4]
  assign _T_13436 = _T_13435 ? _T_10366_2 : _T_13434; // @[Mux.scala 46:16:@12358.4]
  assign _T_13437 = 6'h2 == _T_11317_34; // @[Mux.scala 46:19:@12359.4]
  assign _T_13438 = _T_13437 ? _T_10366_1 : _T_13436; // @[Mux.scala 46:16:@12360.4]
  assign _T_13439 = 6'h1 == _T_11317_34; // @[Mux.scala 46:19:@12361.4]
  assign _T_13440 = _T_13439 ? _T_10366_0 : _T_13438; // @[Mux.scala 46:16:@12362.4]
  assign _T_13478 = 6'h24 == _T_11317_35; // @[Mux.scala 46:19:@12364.4]
  assign _T_13479 = _T_13478 ? _T_10366_35 : 8'h0; // @[Mux.scala 46:16:@12365.4]
  assign _T_13480 = 6'h23 == _T_11317_35; // @[Mux.scala 46:19:@12366.4]
  assign _T_13481 = _T_13480 ? _T_10366_34 : _T_13479; // @[Mux.scala 46:16:@12367.4]
  assign _T_13482 = 6'h22 == _T_11317_35; // @[Mux.scala 46:19:@12368.4]
  assign _T_13483 = _T_13482 ? _T_10366_33 : _T_13481; // @[Mux.scala 46:16:@12369.4]
  assign _T_13484 = 6'h21 == _T_11317_35; // @[Mux.scala 46:19:@12370.4]
  assign _T_13485 = _T_13484 ? _T_10366_32 : _T_13483; // @[Mux.scala 46:16:@12371.4]
  assign _T_13486 = 6'h20 == _T_11317_35; // @[Mux.scala 46:19:@12372.4]
  assign _T_13487 = _T_13486 ? _T_10366_31 : _T_13485; // @[Mux.scala 46:16:@12373.4]
  assign _T_13488 = 6'h1f == _T_11317_35; // @[Mux.scala 46:19:@12374.4]
  assign _T_13489 = _T_13488 ? _T_10366_30 : _T_13487; // @[Mux.scala 46:16:@12375.4]
  assign _T_13490 = 6'h1e == _T_11317_35; // @[Mux.scala 46:19:@12376.4]
  assign _T_13491 = _T_13490 ? _T_10366_29 : _T_13489; // @[Mux.scala 46:16:@12377.4]
  assign _T_13492 = 6'h1d == _T_11317_35; // @[Mux.scala 46:19:@12378.4]
  assign _T_13493 = _T_13492 ? _T_10366_28 : _T_13491; // @[Mux.scala 46:16:@12379.4]
  assign _T_13494 = 6'h1c == _T_11317_35; // @[Mux.scala 46:19:@12380.4]
  assign _T_13495 = _T_13494 ? _T_10366_27 : _T_13493; // @[Mux.scala 46:16:@12381.4]
  assign _T_13496 = 6'h1b == _T_11317_35; // @[Mux.scala 46:19:@12382.4]
  assign _T_13497 = _T_13496 ? _T_10366_26 : _T_13495; // @[Mux.scala 46:16:@12383.4]
  assign _T_13498 = 6'h1a == _T_11317_35; // @[Mux.scala 46:19:@12384.4]
  assign _T_13499 = _T_13498 ? _T_10366_25 : _T_13497; // @[Mux.scala 46:16:@12385.4]
  assign _T_13500 = 6'h19 == _T_11317_35; // @[Mux.scala 46:19:@12386.4]
  assign _T_13501 = _T_13500 ? _T_10366_24 : _T_13499; // @[Mux.scala 46:16:@12387.4]
  assign _T_13502 = 6'h18 == _T_11317_35; // @[Mux.scala 46:19:@12388.4]
  assign _T_13503 = _T_13502 ? _T_10366_23 : _T_13501; // @[Mux.scala 46:16:@12389.4]
  assign _T_13504 = 6'h17 == _T_11317_35; // @[Mux.scala 46:19:@12390.4]
  assign _T_13505 = _T_13504 ? _T_10366_22 : _T_13503; // @[Mux.scala 46:16:@12391.4]
  assign _T_13506 = 6'h16 == _T_11317_35; // @[Mux.scala 46:19:@12392.4]
  assign _T_13507 = _T_13506 ? _T_10366_21 : _T_13505; // @[Mux.scala 46:16:@12393.4]
  assign _T_13508 = 6'h15 == _T_11317_35; // @[Mux.scala 46:19:@12394.4]
  assign _T_13509 = _T_13508 ? _T_10366_20 : _T_13507; // @[Mux.scala 46:16:@12395.4]
  assign _T_13510 = 6'h14 == _T_11317_35; // @[Mux.scala 46:19:@12396.4]
  assign _T_13511 = _T_13510 ? _T_10366_19 : _T_13509; // @[Mux.scala 46:16:@12397.4]
  assign _T_13512 = 6'h13 == _T_11317_35; // @[Mux.scala 46:19:@12398.4]
  assign _T_13513 = _T_13512 ? _T_10366_18 : _T_13511; // @[Mux.scala 46:16:@12399.4]
  assign _T_13514 = 6'h12 == _T_11317_35; // @[Mux.scala 46:19:@12400.4]
  assign _T_13515 = _T_13514 ? _T_10366_17 : _T_13513; // @[Mux.scala 46:16:@12401.4]
  assign _T_13516 = 6'h11 == _T_11317_35; // @[Mux.scala 46:19:@12402.4]
  assign _T_13517 = _T_13516 ? _T_10366_16 : _T_13515; // @[Mux.scala 46:16:@12403.4]
  assign _T_13518 = 6'h10 == _T_11317_35; // @[Mux.scala 46:19:@12404.4]
  assign _T_13519 = _T_13518 ? _T_10366_15 : _T_13517; // @[Mux.scala 46:16:@12405.4]
  assign _T_13520 = 6'hf == _T_11317_35; // @[Mux.scala 46:19:@12406.4]
  assign _T_13521 = _T_13520 ? _T_10366_14 : _T_13519; // @[Mux.scala 46:16:@12407.4]
  assign _T_13522 = 6'he == _T_11317_35; // @[Mux.scala 46:19:@12408.4]
  assign _T_13523 = _T_13522 ? _T_10366_13 : _T_13521; // @[Mux.scala 46:16:@12409.4]
  assign _T_13524 = 6'hd == _T_11317_35; // @[Mux.scala 46:19:@12410.4]
  assign _T_13525 = _T_13524 ? _T_10366_12 : _T_13523; // @[Mux.scala 46:16:@12411.4]
  assign _T_13526 = 6'hc == _T_11317_35; // @[Mux.scala 46:19:@12412.4]
  assign _T_13527 = _T_13526 ? _T_10366_11 : _T_13525; // @[Mux.scala 46:16:@12413.4]
  assign _T_13528 = 6'hb == _T_11317_35; // @[Mux.scala 46:19:@12414.4]
  assign _T_13529 = _T_13528 ? _T_10366_10 : _T_13527; // @[Mux.scala 46:16:@12415.4]
  assign _T_13530 = 6'ha == _T_11317_35; // @[Mux.scala 46:19:@12416.4]
  assign _T_13531 = _T_13530 ? _T_10366_9 : _T_13529; // @[Mux.scala 46:16:@12417.4]
  assign _T_13532 = 6'h9 == _T_11317_35; // @[Mux.scala 46:19:@12418.4]
  assign _T_13533 = _T_13532 ? _T_10366_8 : _T_13531; // @[Mux.scala 46:16:@12419.4]
  assign _T_13534 = 6'h8 == _T_11317_35; // @[Mux.scala 46:19:@12420.4]
  assign _T_13535 = _T_13534 ? _T_10366_7 : _T_13533; // @[Mux.scala 46:16:@12421.4]
  assign _T_13536 = 6'h7 == _T_11317_35; // @[Mux.scala 46:19:@12422.4]
  assign _T_13537 = _T_13536 ? _T_10366_6 : _T_13535; // @[Mux.scala 46:16:@12423.4]
  assign _T_13538 = 6'h6 == _T_11317_35; // @[Mux.scala 46:19:@12424.4]
  assign _T_13539 = _T_13538 ? _T_10366_5 : _T_13537; // @[Mux.scala 46:16:@12425.4]
  assign _T_13540 = 6'h5 == _T_11317_35; // @[Mux.scala 46:19:@12426.4]
  assign _T_13541 = _T_13540 ? _T_10366_4 : _T_13539; // @[Mux.scala 46:16:@12427.4]
  assign _T_13542 = 6'h4 == _T_11317_35; // @[Mux.scala 46:19:@12428.4]
  assign _T_13543 = _T_13542 ? _T_10366_3 : _T_13541; // @[Mux.scala 46:16:@12429.4]
  assign _T_13544 = 6'h3 == _T_11317_35; // @[Mux.scala 46:19:@12430.4]
  assign _T_13545 = _T_13544 ? _T_10366_2 : _T_13543; // @[Mux.scala 46:16:@12431.4]
  assign _T_13546 = 6'h2 == _T_11317_35; // @[Mux.scala 46:19:@12432.4]
  assign _T_13547 = _T_13546 ? _T_10366_1 : _T_13545; // @[Mux.scala 46:16:@12433.4]
  assign _T_13548 = 6'h1 == _T_11317_35; // @[Mux.scala 46:19:@12434.4]
  assign _T_13549 = _T_13548 ? _T_10366_0 : _T_13547; // @[Mux.scala 46:16:@12435.4]
  assign _T_13588 = 6'h25 == _T_11317_36; // @[Mux.scala 46:19:@12437.4]
  assign _T_13589 = _T_13588 ? _T_10366_36 : 8'h0; // @[Mux.scala 46:16:@12438.4]
  assign _T_13590 = 6'h24 == _T_11317_36; // @[Mux.scala 46:19:@12439.4]
  assign _T_13591 = _T_13590 ? _T_10366_35 : _T_13589; // @[Mux.scala 46:16:@12440.4]
  assign _T_13592 = 6'h23 == _T_11317_36; // @[Mux.scala 46:19:@12441.4]
  assign _T_13593 = _T_13592 ? _T_10366_34 : _T_13591; // @[Mux.scala 46:16:@12442.4]
  assign _T_13594 = 6'h22 == _T_11317_36; // @[Mux.scala 46:19:@12443.4]
  assign _T_13595 = _T_13594 ? _T_10366_33 : _T_13593; // @[Mux.scala 46:16:@12444.4]
  assign _T_13596 = 6'h21 == _T_11317_36; // @[Mux.scala 46:19:@12445.4]
  assign _T_13597 = _T_13596 ? _T_10366_32 : _T_13595; // @[Mux.scala 46:16:@12446.4]
  assign _T_13598 = 6'h20 == _T_11317_36; // @[Mux.scala 46:19:@12447.4]
  assign _T_13599 = _T_13598 ? _T_10366_31 : _T_13597; // @[Mux.scala 46:16:@12448.4]
  assign _T_13600 = 6'h1f == _T_11317_36; // @[Mux.scala 46:19:@12449.4]
  assign _T_13601 = _T_13600 ? _T_10366_30 : _T_13599; // @[Mux.scala 46:16:@12450.4]
  assign _T_13602 = 6'h1e == _T_11317_36; // @[Mux.scala 46:19:@12451.4]
  assign _T_13603 = _T_13602 ? _T_10366_29 : _T_13601; // @[Mux.scala 46:16:@12452.4]
  assign _T_13604 = 6'h1d == _T_11317_36; // @[Mux.scala 46:19:@12453.4]
  assign _T_13605 = _T_13604 ? _T_10366_28 : _T_13603; // @[Mux.scala 46:16:@12454.4]
  assign _T_13606 = 6'h1c == _T_11317_36; // @[Mux.scala 46:19:@12455.4]
  assign _T_13607 = _T_13606 ? _T_10366_27 : _T_13605; // @[Mux.scala 46:16:@12456.4]
  assign _T_13608 = 6'h1b == _T_11317_36; // @[Mux.scala 46:19:@12457.4]
  assign _T_13609 = _T_13608 ? _T_10366_26 : _T_13607; // @[Mux.scala 46:16:@12458.4]
  assign _T_13610 = 6'h1a == _T_11317_36; // @[Mux.scala 46:19:@12459.4]
  assign _T_13611 = _T_13610 ? _T_10366_25 : _T_13609; // @[Mux.scala 46:16:@12460.4]
  assign _T_13612 = 6'h19 == _T_11317_36; // @[Mux.scala 46:19:@12461.4]
  assign _T_13613 = _T_13612 ? _T_10366_24 : _T_13611; // @[Mux.scala 46:16:@12462.4]
  assign _T_13614 = 6'h18 == _T_11317_36; // @[Mux.scala 46:19:@12463.4]
  assign _T_13615 = _T_13614 ? _T_10366_23 : _T_13613; // @[Mux.scala 46:16:@12464.4]
  assign _T_13616 = 6'h17 == _T_11317_36; // @[Mux.scala 46:19:@12465.4]
  assign _T_13617 = _T_13616 ? _T_10366_22 : _T_13615; // @[Mux.scala 46:16:@12466.4]
  assign _T_13618 = 6'h16 == _T_11317_36; // @[Mux.scala 46:19:@12467.4]
  assign _T_13619 = _T_13618 ? _T_10366_21 : _T_13617; // @[Mux.scala 46:16:@12468.4]
  assign _T_13620 = 6'h15 == _T_11317_36; // @[Mux.scala 46:19:@12469.4]
  assign _T_13621 = _T_13620 ? _T_10366_20 : _T_13619; // @[Mux.scala 46:16:@12470.4]
  assign _T_13622 = 6'h14 == _T_11317_36; // @[Mux.scala 46:19:@12471.4]
  assign _T_13623 = _T_13622 ? _T_10366_19 : _T_13621; // @[Mux.scala 46:16:@12472.4]
  assign _T_13624 = 6'h13 == _T_11317_36; // @[Mux.scala 46:19:@12473.4]
  assign _T_13625 = _T_13624 ? _T_10366_18 : _T_13623; // @[Mux.scala 46:16:@12474.4]
  assign _T_13626 = 6'h12 == _T_11317_36; // @[Mux.scala 46:19:@12475.4]
  assign _T_13627 = _T_13626 ? _T_10366_17 : _T_13625; // @[Mux.scala 46:16:@12476.4]
  assign _T_13628 = 6'h11 == _T_11317_36; // @[Mux.scala 46:19:@12477.4]
  assign _T_13629 = _T_13628 ? _T_10366_16 : _T_13627; // @[Mux.scala 46:16:@12478.4]
  assign _T_13630 = 6'h10 == _T_11317_36; // @[Mux.scala 46:19:@12479.4]
  assign _T_13631 = _T_13630 ? _T_10366_15 : _T_13629; // @[Mux.scala 46:16:@12480.4]
  assign _T_13632 = 6'hf == _T_11317_36; // @[Mux.scala 46:19:@12481.4]
  assign _T_13633 = _T_13632 ? _T_10366_14 : _T_13631; // @[Mux.scala 46:16:@12482.4]
  assign _T_13634 = 6'he == _T_11317_36; // @[Mux.scala 46:19:@12483.4]
  assign _T_13635 = _T_13634 ? _T_10366_13 : _T_13633; // @[Mux.scala 46:16:@12484.4]
  assign _T_13636 = 6'hd == _T_11317_36; // @[Mux.scala 46:19:@12485.4]
  assign _T_13637 = _T_13636 ? _T_10366_12 : _T_13635; // @[Mux.scala 46:16:@12486.4]
  assign _T_13638 = 6'hc == _T_11317_36; // @[Mux.scala 46:19:@12487.4]
  assign _T_13639 = _T_13638 ? _T_10366_11 : _T_13637; // @[Mux.scala 46:16:@12488.4]
  assign _T_13640 = 6'hb == _T_11317_36; // @[Mux.scala 46:19:@12489.4]
  assign _T_13641 = _T_13640 ? _T_10366_10 : _T_13639; // @[Mux.scala 46:16:@12490.4]
  assign _T_13642 = 6'ha == _T_11317_36; // @[Mux.scala 46:19:@12491.4]
  assign _T_13643 = _T_13642 ? _T_10366_9 : _T_13641; // @[Mux.scala 46:16:@12492.4]
  assign _T_13644 = 6'h9 == _T_11317_36; // @[Mux.scala 46:19:@12493.4]
  assign _T_13645 = _T_13644 ? _T_10366_8 : _T_13643; // @[Mux.scala 46:16:@12494.4]
  assign _T_13646 = 6'h8 == _T_11317_36; // @[Mux.scala 46:19:@12495.4]
  assign _T_13647 = _T_13646 ? _T_10366_7 : _T_13645; // @[Mux.scala 46:16:@12496.4]
  assign _T_13648 = 6'h7 == _T_11317_36; // @[Mux.scala 46:19:@12497.4]
  assign _T_13649 = _T_13648 ? _T_10366_6 : _T_13647; // @[Mux.scala 46:16:@12498.4]
  assign _T_13650 = 6'h6 == _T_11317_36; // @[Mux.scala 46:19:@12499.4]
  assign _T_13651 = _T_13650 ? _T_10366_5 : _T_13649; // @[Mux.scala 46:16:@12500.4]
  assign _T_13652 = 6'h5 == _T_11317_36; // @[Mux.scala 46:19:@12501.4]
  assign _T_13653 = _T_13652 ? _T_10366_4 : _T_13651; // @[Mux.scala 46:16:@12502.4]
  assign _T_13654 = 6'h4 == _T_11317_36; // @[Mux.scala 46:19:@12503.4]
  assign _T_13655 = _T_13654 ? _T_10366_3 : _T_13653; // @[Mux.scala 46:16:@12504.4]
  assign _T_13656 = 6'h3 == _T_11317_36; // @[Mux.scala 46:19:@12505.4]
  assign _T_13657 = _T_13656 ? _T_10366_2 : _T_13655; // @[Mux.scala 46:16:@12506.4]
  assign _T_13658 = 6'h2 == _T_11317_36; // @[Mux.scala 46:19:@12507.4]
  assign _T_13659 = _T_13658 ? _T_10366_1 : _T_13657; // @[Mux.scala 46:16:@12508.4]
  assign _T_13660 = 6'h1 == _T_11317_36; // @[Mux.scala 46:19:@12509.4]
  assign _T_13661 = _T_13660 ? _T_10366_0 : _T_13659; // @[Mux.scala 46:16:@12510.4]
  assign _T_13701 = 6'h26 == _T_11317_37; // @[Mux.scala 46:19:@12512.4]
  assign _T_13702 = _T_13701 ? _T_10366_37 : 8'h0; // @[Mux.scala 46:16:@12513.4]
  assign _T_13703 = 6'h25 == _T_11317_37; // @[Mux.scala 46:19:@12514.4]
  assign _T_13704 = _T_13703 ? _T_10366_36 : _T_13702; // @[Mux.scala 46:16:@12515.4]
  assign _T_13705 = 6'h24 == _T_11317_37; // @[Mux.scala 46:19:@12516.4]
  assign _T_13706 = _T_13705 ? _T_10366_35 : _T_13704; // @[Mux.scala 46:16:@12517.4]
  assign _T_13707 = 6'h23 == _T_11317_37; // @[Mux.scala 46:19:@12518.4]
  assign _T_13708 = _T_13707 ? _T_10366_34 : _T_13706; // @[Mux.scala 46:16:@12519.4]
  assign _T_13709 = 6'h22 == _T_11317_37; // @[Mux.scala 46:19:@12520.4]
  assign _T_13710 = _T_13709 ? _T_10366_33 : _T_13708; // @[Mux.scala 46:16:@12521.4]
  assign _T_13711 = 6'h21 == _T_11317_37; // @[Mux.scala 46:19:@12522.4]
  assign _T_13712 = _T_13711 ? _T_10366_32 : _T_13710; // @[Mux.scala 46:16:@12523.4]
  assign _T_13713 = 6'h20 == _T_11317_37; // @[Mux.scala 46:19:@12524.4]
  assign _T_13714 = _T_13713 ? _T_10366_31 : _T_13712; // @[Mux.scala 46:16:@12525.4]
  assign _T_13715 = 6'h1f == _T_11317_37; // @[Mux.scala 46:19:@12526.4]
  assign _T_13716 = _T_13715 ? _T_10366_30 : _T_13714; // @[Mux.scala 46:16:@12527.4]
  assign _T_13717 = 6'h1e == _T_11317_37; // @[Mux.scala 46:19:@12528.4]
  assign _T_13718 = _T_13717 ? _T_10366_29 : _T_13716; // @[Mux.scala 46:16:@12529.4]
  assign _T_13719 = 6'h1d == _T_11317_37; // @[Mux.scala 46:19:@12530.4]
  assign _T_13720 = _T_13719 ? _T_10366_28 : _T_13718; // @[Mux.scala 46:16:@12531.4]
  assign _T_13721 = 6'h1c == _T_11317_37; // @[Mux.scala 46:19:@12532.4]
  assign _T_13722 = _T_13721 ? _T_10366_27 : _T_13720; // @[Mux.scala 46:16:@12533.4]
  assign _T_13723 = 6'h1b == _T_11317_37; // @[Mux.scala 46:19:@12534.4]
  assign _T_13724 = _T_13723 ? _T_10366_26 : _T_13722; // @[Mux.scala 46:16:@12535.4]
  assign _T_13725 = 6'h1a == _T_11317_37; // @[Mux.scala 46:19:@12536.4]
  assign _T_13726 = _T_13725 ? _T_10366_25 : _T_13724; // @[Mux.scala 46:16:@12537.4]
  assign _T_13727 = 6'h19 == _T_11317_37; // @[Mux.scala 46:19:@12538.4]
  assign _T_13728 = _T_13727 ? _T_10366_24 : _T_13726; // @[Mux.scala 46:16:@12539.4]
  assign _T_13729 = 6'h18 == _T_11317_37; // @[Mux.scala 46:19:@12540.4]
  assign _T_13730 = _T_13729 ? _T_10366_23 : _T_13728; // @[Mux.scala 46:16:@12541.4]
  assign _T_13731 = 6'h17 == _T_11317_37; // @[Mux.scala 46:19:@12542.4]
  assign _T_13732 = _T_13731 ? _T_10366_22 : _T_13730; // @[Mux.scala 46:16:@12543.4]
  assign _T_13733 = 6'h16 == _T_11317_37; // @[Mux.scala 46:19:@12544.4]
  assign _T_13734 = _T_13733 ? _T_10366_21 : _T_13732; // @[Mux.scala 46:16:@12545.4]
  assign _T_13735 = 6'h15 == _T_11317_37; // @[Mux.scala 46:19:@12546.4]
  assign _T_13736 = _T_13735 ? _T_10366_20 : _T_13734; // @[Mux.scala 46:16:@12547.4]
  assign _T_13737 = 6'h14 == _T_11317_37; // @[Mux.scala 46:19:@12548.4]
  assign _T_13738 = _T_13737 ? _T_10366_19 : _T_13736; // @[Mux.scala 46:16:@12549.4]
  assign _T_13739 = 6'h13 == _T_11317_37; // @[Mux.scala 46:19:@12550.4]
  assign _T_13740 = _T_13739 ? _T_10366_18 : _T_13738; // @[Mux.scala 46:16:@12551.4]
  assign _T_13741 = 6'h12 == _T_11317_37; // @[Mux.scala 46:19:@12552.4]
  assign _T_13742 = _T_13741 ? _T_10366_17 : _T_13740; // @[Mux.scala 46:16:@12553.4]
  assign _T_13743 = 6'h11 == _T_11317_37; // @[Mux.scala 46:19:@12554.4]
  assign _T_13744 = _T_13743 ? _T_10366_16 : _T_13742; // @[Mux.scala 46:16:@12555.4]
  assign _T_13745 = 6'h10 == _T_11317_37; // @[Mux.scala 46:19:@12556.4]
  assign _T_13746 = _T_13745 ? _T_10366_15 : _T_13744; // @[Mux.scala 46:16:@12557.4]
  assign _T_13747 = 6'hf == _T_11317_37; // @[Mux.scala 46:19:@12558.4]
  assign _T_13748 = _T_13747 ? _T_10366_14 : _T_13746; // @[Mux.scala 46:16:@12559.4]
  assign _T_13749 = 6'he == _T_11317_37; // @[Mux.scala 46:19:@12560.4]
  assign _T_13750 = _T_13749 ? _T_10366_13 : _T_13748; // @[Mux.scala 46:16:@12561.4]
  assign _T_13751 = 6'hd == _T_11317_37; // @[Mux.scala 46:19:@12562.4]
  assign _T_13752 = _T_13751 ? _T_10366_12 : _T_13750; // @[Mux.scala 46:16:@12563.4]
  assign _T_13753 = 6'hc == _T_11317_37; // @[Mux.scala 46:19:@12564.4]
  assign _T_13754 = _T_13753 ? _T_10366_11 : _T_13752; // @[Mux.scala 46:16:@12565.4]
  assign _T_13755 = 6'hb == _T_11317_37; // @[Mux.scala 46:19:@12566.4]
  assign _T_13756 = _T_13755 ? _T_10366_10 : _T_13754; // @[Mux.scala 46:16:@12567.4]
  assign _T_13757 = 6'ha == _T_11317_37; // @[Mux.scala 46:19:@12568.4]
  assign _T_13758 = _T_13757 ? _T_10366_9 : _T_13756; // @[Mux.scala 46:16:@12569.4]
  assign _T_13759 = 6'h9 == _T_11317_37; // @[Mux.scala 46:19:@12570.4]
  assign _T_13760 = _T_13759 ? _T_10366_8 : _T_13758; // @[Mux.scala 46:16:@12571.4]
  assign _T_13761 = 6'h8 == _T_11317_37; // @[Mux.scala 46:19:@12572.4]
  assign _T_13762 = _T_13761 ? _T_10366_7 : _T_13760; // @[Mux.scala 46:16:@12573.4]
  assign _T_13763 = 6'h7 == _T_11317_37; // @[Mux.scala 46:19:@12574.4]
  assign _T_13764 = _T_13763 ? _T_10366_6 : _T_13762; // @[Mux.scala 46:16:@12575.4]
  assign _T_13765 = 6'h6 == _T_11317_37; // @[Mux.scala 46:19:@12576.4]
  assign _T_13766 = _T_13765 ? _T_10366_5 : _T_13764; // @[Mux.scala 46:16:@12577.4]
  assign _T_13767 = 6'h5 == _T_11317_37; // @[Mux.scala 46:19:@12578.4]
  assign _T_13768 = _T_13767 ? _T_10366_4 : _T_13766; // @[Mux.scala 46:16:@12579.4]
  assign _T_13769 = 6'h4 == _T_11317_37; // @[Mux.scala 46:19:@12580.4]
  assign _T_13770 = _T_13769 ? _T_10366_3 : _T_13768; // @[Mux.scala 46:16:@12581.4]
  assign _T_13771 = 6'h3 == _T_11317_37; // @[Mux.scala 46:19:@12582.4]
  assign _T_13772 = _T_13771 ? _T_10366_2 : _T_13770; // @[Mux.scala 46:16:@12583.4]
  assign _T_13773 = 6'h2 == _T_11317_37; // @[Mux.scala 46:19:@12584.4]
  assign _T_13774 = _T_13773 ? _T_10366_1 : _T_13772; // @[Mux.scala 46:16:@12585.4]
  assign _T_13775 = 6'h1 == _T_11317_37; // @[Mux.scala 46:19:@12586.4]
  assign _T_13776 = _T_13775 ? _T_10366_0 : _T_13774; // @[Mux.scala 46:16:@12587.4]
  assign _T_13817 = 6'h27 == _T_11317_38; // @[Mux.scala 46:19:@12589.4]
  assign _T_13818 = _T_13817 ? _T_10366_38 : 8'h0; // @[Mux.scala 46:16:@12590.4]
  assign _T_13819 = 6'h26 == _T_11317_38; // @[Mux.scala 46:19:@12591.4]
  assign _T_13820 = _T_13819 ? _T_10366_37 : _T_13818; // @[Mux.scala 46:16:@12592.4]
  assign _T_13821 = 6'h25 == _T_11317_38; // @[Mux.scala 46:19:@12593.4]
  assign _T_13822 = _T_13821 ? _T_10366_36 : _T_13820; // @[Mux.scala 46:16:@12594.4]
  assign _T_13823 = 6'h24 == _T_11317_38; // @[Mux.scala 46:19:@12595.4]
  assign _T_13824 = _T_13823 ? _T_10366_35 : _T_13822; // @[Mux.scala 46:16:@12596.4]
  assign _T_13825 = 6'h23 == _T_11317_38; // @[Mux.scala 46:19:@12597.4]
  assign _T_13826 = _T_13825 ? _T_10366_34 : _T_13824; // @[Mux.scala 46:16:@12598.4]
  assign _T_13827 = 6'h22 == _T_11317_38; // @[Mux.scala 46:19:@12599.4]
  assign _T_13828 = _T_13827 ? _T_10366_33 : _T_13826; // @[Mux.scala 46:16:@12600.4]
  assign _T_13829 = 6'h21 == _T_11317_38; // @[Mux.scala 46:19:@12601.4]
  assign _T_13830 = _T_13829 ? _T_10366_32 : _T_13828; // @[Mux.scala 46:16:@12602.4]
  assign _T_13831 = 6'h20 == _T_11317_38; // @[Mux.scala 46:19:@12603.4]
  assign _T_13832 = _T_13831 ? _T_10366_31 : _T_13830; // @[Mux.scala 46:16:@12604.4]
  assign _T_13833 = 6'h1f == _T_11317_38; // @[Mux.scala 46:19:@12605.4]
  assign _T_13834 = _T_13833 ? _T_10366_30 : _T_13832; // @[Mux.scala 46:16:@12606.4]
  assign _T_13835 = 6'h1e == _T_11317_38; // @[Mux.scala 46:19:@12607.4]
  assign _T_13836 = _T_13835 ? _T_10366_29 : _T_13834; // @[Mux.scala 46:16:@12608.4]
  assign _T_13837 = 6'h1d == _T_11317_38; // @[Mux.scala 46:19:@12609.4]
  assign _T_13838 = _T_13837 ? _T_10366_28 : _T_13836; // @[Mux.scala 46:16:@12610.4]
  assign _T_13839 = 6'h1c == _T_11317_38; // @[Mux.scala 46:19:@12611.4]
  assign _T_13840 = _T_13839 ? _T_10366_27 : _T_13838; // @[Mux.scala 46:16:@12612.4]
  assign _T_13841 = 6'h1b == _T_11317_38; // @[Mux.scala 46:19:@12613.4]
  assign _T_13842 = _T_13841 ? _T_10366_26 : _T_13840; // @[Mux.scala 46:16:@12614.4]
  assign _T_13843 = 6'h1a == _T_11317_38; // @[Mux.scala 46:19:@12615.4]
  assign _T_13844 = _T_13843 ? _T_10366_25 : _T_13842; // @[Mux.scala 46:16:@12616.4]
  assign _T_13845 = 6'h19 == _T_11317_38; // @[Mux.scala 46:19:@12617.4]
  assign _T_13846 = _T_13845 ? _T_10366_24 : _T_13844; // @[Mux.scala 46:16:@12618.4]
  assign _T_13847 = 6'h18 == _T_11317_38; // @[Mux.scala 46:19:@12619.4]
  assign _T_13848 = _T_13847 ? _T_10366_23 : _T_13846; // @[Mux.scala 46:16:@12620.4]
  assign _T_13849 = 6'h17 == _T_11317_38; // @[Mux.scala 46:19:@12621.4]
  assign _T_13850 = _T_13849 ? _T_10366_22 : _T_13848; // @[Mux.scala 46:16:@12622.4]
  assign _T_13851 = 6'h16 == _T_11317_38; // @[Mux.scala 46:19:@12623.4]
  assign _T_13852 = _T_13851 ? _T_10366_21 : _T_13850; // @[Mux.scala 46:16:@12624.4]
  assign _T_13853 = 6'h15 == _T_11317_38; // @[Mux.scala 46:19:@12625.4]
  assign _T_13854 = _T_13853 ? _T_10366_20 : _T_13852; // @[Mux.scala 46:16:@12626.4]
  assign _T_13855 = 6'h14 == _T_11317_38; // @[Mux.scala 46:19:@12627.4]
  assign _T_13856 = _T_13855 ? _T_10366_19 : _T_13854; // @[Mux.scala 46:16:@12628.4]
  assign _T_13857 = 6'h13 == _T_11317_38; // @[Mux.scala 46:19:@12629.4]
  assign _T_13858 = _T_13857 ? _T_10366_18 : _T_13856; // @[Mux.scala 46:16:@12630.4]
  assign _T_13859 = 6'h12 == _T_11317_38; // @[Mux.scala 46:19:@12631.4]
  assign _T_13860 = _T_13859 ? _T_10366_17 : _T_13858; // @[Mux.scala 46:16:@12632.4]
  assign _T_13861 = 6'h11 == _T_11317_38; // @[Mux.scala 46:19:@12633.4]
  assign _T_13862 = _T_13861 ? _T_10366_16 : _T_13860; // @[Mux.scala 46:16:@12634.4]
  assign _T_13863 = 6'h10 == _T_11317_38; // @[Mux.scala 46:19:@12635.4]
  assign _T_13864 = _T_13863 ? _T_10366_15 : _T_13862; // @[Mux.scala 46:16:@12636.4]
  assign _T_13865 = 6'hf == _T_11317_38; // @[Mux.scala 46:19:@12637.4]
  assign _T_13866 = _T_13865 ? _T_10366_14 : _T_13864; // @[Mux.scala 46:16:@12638.4]
  assign _T_13867 = 6'he == _T_11317_38; // @[Mux.scala 46:19:@12639.4]
  assign _T_13868 = _T_13867 ? _T_10366_13 : _T_13866; // @[Mux.scala 46:16:@12640.4]
  assign _T_13869 = 6'hd == _T_11317_38; // @[Mux.scala 46:19:@12641.4]
  assign _T_13870 = _T_13869 ? _T_10366_12 : _T_13868; // @[Mux.scala 46:16:@12642.4]
  assign _T_13871 = 6'hc == _T_11317_38; // @[Mux.scala 46:19:@12643.4]
  assign _T_13872 = _T_13871 ? _T_10366_11 : _T_13870; // @[Mux.scala 46:16:@12644.4]
  assign _T_13873 = 6'hb == _T_11317_38; // @[Mux.scala 46:19:@12645.4]
  assign _T_13874 = _T_13873 ? _T_10366_10 : _T_13872; // @[Mux.scala 46:16:@12646.4]
  assign _T_13875 = 6'ha == _T_11317_38; // @[Mux.scala 46:19:@12647.4]
  assign _T_13876 = _T_13875 ? _T_10366_9 : _T_13874; // @[Mux.scala 46:16:@12648.4]
  assign _T_13877 = 6'h9 == _T_11317_38; // @[Mux.scala 46:19:@12649.4]
  assign _T_13878 = _T_13877 ? _T_10366_8 : _T_13876; // @[Mux.scala 46:16:@12650.4]
  assign _T_13879 = 6'h8 == _T_11317_38; // @[Mux.scala 46:19:@12651.4]
  assign _T_13880 = _T_13879 ? _T_10366_7 : _T_13878; // @[Mux.scala 46:16:@12652.4]
  assign _T_13881 = 6'h7 == _T_11317_38; // @[Mux.scala 46:19:@12653.4]
  assign _T_13882 = _T_13881 ? _T_10366_6 : _T_13880; // @[Mux.scala 46:16:@12654.4]
  assign _T_13883 = 6'h6 == _T_11317_38; // @[Mux.scala 46:19:@12655.4]
  assign _T_13884 = _T_13883 ? _T_10366_5 : _T_13882; // @[Mux.scala 46:16:@12656.4]
  assign _T_13885 = 6'h5 == _T_11317_38; // @[Mux.scala 46:19:@12657.4]
  assign _T_13886 = _T_13885 ? _T_10366_4 : _T_13884; // @[Mux.scala 46:16:@12658.4]
  assign _T_13887 = 6'h4 == _T_11317_38; // @[Mux.scala 46:19:@12659.4]
  assign _T_13888 = _T_13887 ? _T_10366_3 : _T_13886; // @[Mux.scala 46:16:@12660.4]
  assign _T_13889 = 6'h3 == _T_11317_38; // @[Mux.scala 46:19:@12661.4]
  assign _T_13890 = _T_13889 ? _T_10366_2 : _T_13888; // @[Mux.scala 46:16:@12662.4]
  assign _T_13891 = 6'h2 == _T_11317_38; // @[Mux.scala 46:19:@12663.4]
  assign _T_13892 = _T_13891 ? _T_10366_1 : _T_13890; // @[Mux.scala 46:16:@12664.4]
  assign _T_13893 = 6'h1 == _T_11317_38; // @[Mux.scala 46:19:@12665.4]
  assign _T_13894 = _T_13893 ? _T_10366_0 : _T_13892; // @[Mux.scala 46:16:@12666.4]
  assign _T_13936 = 6'h28 == _T_11317_39; // @[Mux.scala 46:19:@12668.4]
  assign _T_13937 = _T_13936 ? _T_10366_39 : 8'h0; // @[Mux.scala 46:16:@12669.4]
  assign _T_13938 = 6'h27 == _T_11317_39; // @[Mux.scala 46:19:@12670.4]
  assign _T_13939 = _T_13938 ? _T_10366_38 : _T_13937; // @[Mux.scala 46:16:@12671.4]
  assign _T_13940 = 6'h26 == _T_11317_39; // @[Mux.scala 46:19:@12672.4]
  assign _T_13941 = _T_13940 ? _T_10366_37 : _T_13939; // @[Mux.scala 46:16:@12673.4]
  assign _T_13942 = 6'h25 == _T_11317_39; // @[Mux.scala 46:19:@12674.4]
  assign _T_13943 = _T_13942 ? _T_10366_36 : _T_13941; // @[Mux.scala 46:16:@12675.4]
  assign _T_13944 = 6'h24 == _T_11317_39; // @[Mux.scala 46:19:@12676.4]
  assign _T_13945 = _T_13944 ? _T_10366_35 : _T_13943; // @[Mux.scala 46:16:@12677.4]
  assign _T_13946 = 6'h23 == _T_11317_39; // @[Mux.scala 46:19:@12678.4]
  assign _T_13947 = _T_13946 ? _T_10366_34 : _T_13945; // @[Mux.scala 46:16:@12679.4]
  assign _T_13948 = 6'h22 == _T_11317_39; // @[Mux.scala 46:19:@12680.4]
  assign _T_13949 = _T_13948 ? _T_10366_33 : _T_13947; // @[Mux.scala 46:16:@12681.4]
  assign _T_13950 = 6'h21 == _T_11317_39; // @[Mux.scala 46:19:@12682.4]
  assign _T_13951 = _T_13950 ? _T_10366_32 : _T_13949; // @[Mux.scala 46:16:@12683.4]
  assign _T_13952 = 6'h20 == _T_11317_39; // @[Mux.scala 46:19:@12684.4]
  assign _T_13953 = _T_13952 ? _T_10366_31 : _T_13951; // @[Mux.scala 46:16:@12685.4]
  assign _T_13954 = 6'h1f == _T_11317_39; // @[Mux.scala 46:19:@12686.4]
  assign _T_13955 = _T_13954 ? _T_10366_30 : _T_13953; // @[Mux.scala 46:16:@12687.4]
  assign _T_13956 = 6'h1e == _T_11317_39; // @[Mux.scala 46:19:@12688.4]
  assign _T_13957 = _T_13956 ? _T_10366_29 : _T_13955; // @[Mux.scala 46:16:@12689.4]
  assign _T_13958 = 6'h1d == _T_11317_39; // @[Mux.scala 46:19:@12690.4]
  assign _T_13959 = _T_13958 ? _T_10366_28 : _T_13957; // @[Mux.scala 46:16:@12691.4]
  assign _T_13960 = 6'h1c == _T_11317_39; // @[Mux.scala 46:19:@12692.4]
  assign _T_13961 = _T_13960 ? _T_10366_27 : _T_13959; // @[Mux.scala 46:16:@12693.4]
  assign _T_13962 = 6'h1b == _T_11317_39; // @[Mux.scala 46:19:@12694.4]
  assign _T_13963 = _T_13962 ? _T_10366_26 : _T_13961; // @[Mux.scala 46:16:@12695.4]
  assign _T_13964 = 6'h1a == _T_11317_39; // @[Mux.scala 46:19:@12696.4]
  assign _T_13965 = _T_13964 ? _T_10366_25 : _T_13963; // @[Mux.scala 46:16:@12697.4]
  assign _T_13966 = 6'h19 == _T_11317_39; // @[Mux.scala 46:19:@12698.4]
  assign _T_13967 = _T_13966 ? _T_10366_24 : _T_13965; // @[Mux.scala 46:16:@12699.4]
  assign _T_13968 = 6'h18 == _T_11317_39; // @[Mux.scala 46:19:@12700.4]
  assign _T_13969 = _T_13968 ? _T_10366_23 : _T_13967; // @[Mux.scala 46:16:@12701.4]
  assign _T_13970 = 6'h17 == _T_11317_39; // @[Mux.scala 46:19:@12702.4]
  assign _T_13971 = _T_13970 ? _T_10366_22 : _T_13969; // @[Mux.scala 46:16:@12703.4]
  assign _T_13972 = 6'h16 == _T_11317_39; // @[Mux.scala 46:19:@12704.4]
  assign _T_13973 = _T_13972 ? _T_10366_21 : _T_13971; // @[Mux.scala 46:16:@12705.4]
  assign _T_13974 = 6'h15 == _T_11317_39; // @[Mux.scala 46:19:@12706.4]
  assign _T_13975 = _T_13974 ? _T_10366_20 : _T_13973; // @[Mux.scala 46:16:@12707.4]
  assign _T_13976 = 6'h14 == _T_11317_39; // @[Mux.scala 46:19:@12708.4]
  assign _T_13977 = _T_13976 ? _T_10366_19 : _T_13975; // @[Mux.scala 46:16:@12709.4]
  assign _T_13978 = 6'h13 == _T_11317_39; // @[Mux.scala 46:19:@12710.4]
  assign _T_13979 = _T_13978 ? _T_10366_18 : _T_13977; // @[Mux.scala 46:16:@12711.4]
  assign _T_13980 = 6'h12 == _T_11317_39; // @[Mux.scala 46:19:@12712.4]
  assign _T_13981 = _T_13980 ? _T_10366_17 : _T_13979; // @[Mux.scala 46:16:@12713.4]
  assign _T_13982 = 6'h11 == _T_11317_39; // @[Mux.scala 46:19:@12714.4]
  assign _T_13983 = _T_13982 ? _T_10366_16 : _T_13981; // @[Mux.scala 46:16:@12715.4]
  assign _T_13984 = 6'h10 == _T_11317_39; // @[Mux.scala 46:19:@12716.4]
  assign _T_13985 = _T_13984 ? _T_10366_15 : _T_13983; // @[Mux.scala 46:16:@12717.4]
  assign _T_13986 = 6'hf == _T_11317_39; // @[Mux.scala 46:19:@12718.4]
  assign _T_13987 = _T_13986 ? _T_10366_14 : _T_13985; // @[Mux.scala 46:16:@12719.4]
  assign _T_13988 = 6'he == _T_11317_39; // @[Mux.scala 46:19:@12720.4]
  assign _T_13989 = _T_13988 ? _T_10366_13 : _T_13987; // @[Mux.scala 46:16:@12721.4]
  assign _T_13990 = 6'hd == _T_11317_39; // @[Mux.scala 46:19:@12722.4]
  assign _T_13991 = _T_13990 ? _T_10366_12 : _T_13989; // @[Mux.scala 46:16:@12723.4]
  assign _T_13992 = 6'hc == _T_11317_39; // @[Mux.scala 46:19:@12724.4]
  assign _T_13993 = _T_13992 ? _T_10366_11 : _T_13991; // @[Mux.scala 46:16:@12725.4]
  assign _T_13994 = 6'hb == _T_11317_39; // @[Mux.scala 46:19:@12726.4]
  assign _T_13995 = _T_13994 ? _T_10366_10 : _T_13993; // @[Mux.scala 46:16:@12727.4]
  assign _T_13996 = 6'ha == _T_11317_39; // @[Mux.scala 46:19:@12728.4]
  assign _T_13997 = _T_13996 ? _T_10366_9 : _T_13995; // @[Mux.scala 46:16:@12729.4]
  assign _T_13998 = 6'h9 == _T_11317_39; // @[Mux.scala 46:19:@12730.4]
  assign _T_13999 = _T_13998 ? _T_10366_8 : _T_13997; // @[Mux.scala 46:16:@12731.4]
  assign _T_14000 = 6'h8 == _T_11317_39; // @[Mux.scala 46:19:@12732.4]
  assign _T_14001 = _T_14000 ? _T_10366_7 : _T_13999; // @[Mux.scala 46:16:@12733.4]
  assign _T_14002 = 6'h7 == _T_11317_39; // @[Mux.scala 46:19:@12734.4]
  assign _T_14003 = _T_14002 ? _T_10366_6 : _T_14001; // @[Mux.scala 46:16:@12735.4]
  assign _T_14004 = 6'h6 == _T_11317_39; // @[Mux.scala 46:19:@12736.4]
  assign _T_14005 = _T_14004 ? _T_10366_5 : _T_14003; // @[Mux.scala 46:16:@12737.4]
  assign _T_14006 = 6'h5 == _T_11317_39; // @[Mux.scala 46:19:@12738.4]
  assign _T_14007 = _T_14006 ? _T_10366_4 : _T_14005; // @[Mux.scala 46:16:@12739.4]
  assign _T_14008 = 6'h4 == _T_11317_39; // @[Mux.scala 46:19:@12740.4]
  assign _T_14009 = _T_14008 ? _T_10366_3 : _T_14007; // @[Mux.scala 46:16:@12741.4]
  assign _T_14010 = 6'h3 == _T_11317_39; // @[Mux.scala 46:19:@12742.4]
  assign _T_14011 = _T_14010 ? _T_10366_2 : _T_14009; // @[Mux.scala 46:16:@12743.4]
  assign _T_14012 = 6'h2 == _T_11317_39; // @[Mux.scala 46:19:@12744.4]
  assign _T_14013 = _T_14012 ? _T_10366_1 : _T_14011; // @[Mux.scala 46:16:@12745.4]
  assign _T_14014 = 6'h1 == _T_11317_39; // @[Mux.scala 46:19:@12746.4]
  assign _T_14015 = _T_14014 ? _T_10366_0 : _T_14013; // @[Mux.scala 46:16:@12747.4]
  assign _T_14058 = 6'h29 == _T_11317_40; // @[Mux.scala 46:19:@12749.4]
  assign _T_14059 = _T_14058 ? _T_10366_40 : 8'h0; // @[Mux.scala 46:16:@12750.4]
  assign _T_14060 = 6'h28 == _T_11317_40; // @[Mux.scala 46:19:@12751.4]
  assign _T_14061 = _T_14060 ? _T_10366_39 : _T_14059; // @[Mux.scala 46:16:@12752.4]
  assign _T_14062 = 6'h27 == _T_11317_40; // @[Mux.scala 46:19:@12753.4]
  assign _T_14063 = _T_14062 ? _T_10366_38 : _T_14061; // @[Mux.scala 46:16:@12754.4]
  assign _T_14064 = 6'h26 == _T_11317_40; // @[Mux.scala 46:19:@12755.4]
  assign _T_14065 = _T_14064 ? _T_10366_37 : _T_14063; // @[Mux.scala 46:16:@12756.4]
  assign _T_14066 = 6'h25 == _T_11317_40; // @[Mux.scala 46:19:@12757.4]
  assign _T_14067 = _T_14066 ? _T_10366_36 : _T_14065; // @[Mux.scala 46:16:@12758.4]
  assign _T_14068 = 6'h24 == _T_11317_40; // @[Mux.scala 46:19:@12759.4]
  assign _T_14069 = _T_14068 ? _T_10366_35 : _T_14067; // @[Mux.scala 46:16:@12760.4]
  assign _T_14070 = 6'h23 == _T_11317_40; // @[Mux.scala 46:19:@12761.4]
  assign _T_14071 = _T_14070 ? _T_10366_34 : _T_14069; // @[Mux.scala 46:16:@12762.4]
  assign _T_14072 = 6'h22 == _T_11317_40; // @[Mux.scala 46:19:@12763.4]
  assign _T_14073 = _T_14072 ? _T_10366_33 : _T_14071; // @[Mux.scala 46:16:@12764.4]
  assign _T_14074 = 6'h21 == _T_11317_40; // @[Mux.scala 46:19:@12765.4]
  assign _T_14075 = _T_14074 ? _T_10366_32 : _T_14073; // @[Mux.scala 46:16:@12766.4]
  assign _T_14076 = 6'h20 == _T_11317_40; // @[Mux.scala 46:19:@12767.4]
  assign _T_14077 = _T_14076 ? _T_10366_31 : _T_14075; // @[Mux.scala 46:16:@12768.4]
  assign _T_14078 = 6'h1f == _T_11317_40; // @[Mux.scala 46:19:@12769.4]
  assign _T_14079 = _T_14078 ? _T_10366_30 : _T_14077; // @[Mux.scala 46:16:@12770.4]
  assign _T_14080 = 6'h1e == _T_11317_40; // @[Mux.scala 46:19:@12771.4]
  assign _T_14081 = _T_14080 ? _T_10366_29 : _T_14079; // @[Mux.scala 46:16:@12772.4]
  assign _T_14082 = 6'h1d == _T_11317_40; // @[Mux.scala 46:19:@12773.4]
  assign _T_14083 = _T_14082 ? _T_10366_28 : _T_14081; // @[Mux.scala 46:16:@12774.4]
  assign _T_14084 = 6'h1c == _T_11317_40; // @[Mux.scala 46:19:@12775.4]
  assign _T_14085 = _T_14084 ? _T_10366_27 : _T_14083; // @[Mux.scala 46:16:@12776.4]
  assign _T_14086 = 6'h1b == _T_11317_40; // @[Mux.scala 46:19:@12777.4]
  assign _T_14087 = _T_14086 ? _T_10366_26 : _T_14085; // @[Mux.scala 46:16:@12778.4]
  assign _T_14088 = 6'h1a == _T_11317_40; // @[Mux.scala 46:19:@12779.4]
  assign _T_14089 = _T_14088 ? _T_10366_25 : _T_14087; // @[Mux.scala 46:16:@12780.4]
  assign _T_14090 = 6'h19 == _T_11317_40; // @[Mux.scala 46:19:@12781.4]
  assign _T_14091 = _T_14090 ? _T_10366_24 : _T_14089; // @[Mux.scala 46:16:@12782.4]
  assign _T_14092 = 6'h18 == _T_11317_40; // @[Mux.scala 46:19:@12783.4]
  assign _T_14093 = _T_14092 ? _T_10366_23 : _T_14091; // @[Mux.scala 46:16:@12784.4]
  assign _T_14094 = 6'h17 == _T_11317_40; // @[Mux.scala 46:19:@12785.4]
  assign _T_14095 = _T_14094 ? _T_10366_22 : _T_14093; // @[Mux.scala 46:16:@12786.4]
  assign _T_14096 = 6'h16 == _T_11317_40; // @[Mux.scala 46:19:@12787.4]
  assign _T_14097 = _T_14096 ? _T_10366_21 : _T_14095; // @[Mux.scala 46:16:@12788.4]
  assign _T_14098 = 6'h15 == _T_11317_40; // @[Mux.scala 46:19:@12789.4]
  assign _T_14099 = _T_14098 ? _T_10366_20 : _T_14097; // @[Mux.scala 46:16:@12790.4]
  assign _T_14100 = 6'h14 == _T_11317_40; // @[Mux.scala 46:19:@12791.4]
  assign _T_14101 = _T_14100 ? _T_10366_19 : _T_14099; // @[Mux.scala 46:16:@12792.4]
  assign _T_14102 = 6'h13 == _T_11317_40; // @[Mux.scala 46:19:@12793.4]
  assign _T_14103 = _T_14102 ? _T_10366_18 : _T_14101; // @[Mux.scala 46:16:@12794.4]
  assign _T_14104 = 6'h12 == _T_11317_40; // @[Mux.scala 46:19:@12795.4]
  assign _T_14105 = _T_14104 ? _T_10366_17 : _T_14103; // @[Mux.scala 46:16:@12796.4]
  assign _T_14106 = 6'h11 == _T_11317_40; // @[Mux.scala 46:19:@12797.4]
  assign _T_14107 = _T_14106 ? _T_10366_16 : _T_14105; // @[Mux.scala 46:16:@12798.4]
  assign _T_14108 = 6'h10 == _T_11317_40; // @[Mux.scala 46:19:@12799.4]
  assign _T_14109 = _T_14108 ? _T_10366_15 : _T_14107; // @[Mux.scala 46:16:@12800.4]
  assign _T_14110 = 6'hf == _T_11317_40; // @[Mux.scala 46:19:@12801.4]
  assign _T_14111 = _T_14110 ? _T_10366_14 : _T_14109; // @[Mux.scala 46:16:@12802.4]
  assign _T_14112 = 6'he == _T_11317_40; // @[Mux.scala 46:19:@12803.4]
  assign _T_14113 = _T_14112 ? _T_10366_13 : _T_14111; // @[Mux.scala 46:16:@12804.4]
  assign _T_14114 = 6'hd == _T_11317_40; // @[Mux.scala 46:19:@12805.4]
  assign _T_14115 = _T_14114 ? _T_10366_12 : _T_14113; // @[Mux.scala 46:16:@12806.4]
  assign _T_14116 = 6'hc == _T_11317_40; // @[Mux.scala 46:19:@12807.4]
  assign _T_14117 = _T_14116 ? _T_10366_11 : _T_14115; // @[Mux.scala 46:16:@12808.4]
  assign _T_14118 = 6'hb == _T_11317_40; // @[Mux.scala 46:19:@12809.4]
  assign _T_14119 = _T_14118 ? _T_10366_10 : _T_14117; // @[Mux.scala 46:16:@12810.4]
  assign _T_14120 = 6'ha == _T_11317_40; // @[Mux.scala 46:19:@12811.4]
  assign _T_14121 = _T_14120 ? _T_10366_9 : _T_14119; // @[Mux.scala 46:16:@12812.4]
  assign _T_14122 = 6'h9 == _T_11317_40; // @[Mux.scala 46:19:@12813.4]
  assign _T_14123 = _T_14122 ? _T_10366_8 : _T_14121; // @[Mux.scala 46:16:@12814.4]
  assign _T_14124 = 6'h8 == _T_11317_40; // @[Mux.scala 46:19:@12815.4]
  assign _T_14125 = _T_14124 ? _T_10366_7 : _T_14123; // @[Mux.scala 46:16:@12816.4]
  assign _T_14126 = 6'h7 == _T_11317_40; // @[Mux.scala 46:19:@12817.4]
  assign _T_14127 = _T_14126 ? _T_10366_6 : _T_14125; // @[Mux.scala 46:16:@12818.4]
  assign _T_14128 = 6'h6 == _T_11317_40; // @[Mux.scala 46:19:@12819.4]
  assign _T_14129 = _T_14128 ? _T_10366_5 : _T_14127; // @[Mux.scala 46:16:@12820.4]
  assign _T_14130 = 6'h5 == _T_11317_40; // @[Mux.scala 46:19:@12821.4]
  assign _T_14131 = _T_14130 ? _T_10366_4 : _T_14129; // @[Mux.scala 46:16:@12822.4]
  assign _T_14132 = 6'h4 == _T_11317_40; // @[Mux.scala 46:19:@12823.4]
  assign _T_14133 = _T_14132 ? _T_10366_3 : _T_14131; // @[Mux.scala 46:16:@12824.4]
  assign _T_14134 = 6'h3 == _T_11317_40; // @[Mux.scala 46:19:@12825.4]
  assign _T_14135 = _T_14134 ? _T_10366_2 : _T_14133; // @[Mux.scala 46:16:@12826.4]
  assign _T_14136 = 6'h2 == _T_11317_40; // @[Mux.scala 46:19:@12827.4]
  assign _T_14137 = _T_14136 ? _T_10366_1 : _T_14135; // @[Mux.scala 46:16:@12828.4]
  assign _T_14138 = 6'h1 == _T_11317_40; // @[Mux.scala 46:19:@12829.4]
  assign _T_14139 = _T_14138 ? _T_10366_0 : _T_14137; // @[Mux.scala 46:16:@12830.4]
  assign _T_14183 = 6'h2a == _T_11317_41; // @[Mux.scala 46:19:@12832.4]
  assign _T_14184 = _T_14183 ? _T_10366_41 : 8'h0; // @[Mux.scala 46:16:@12833.4]
  assign _T_14185 = 6'h29 == _T_11317_41; // @[Mux.scala 46:19:@12834.4]
  assign _T_14186 = _T_14185 ? _T_10366_40 : _T_14184; // @[Mux.scala 46:16:@12835.4]
  assign _T_14187 = 6'h28 == _T_11317_41; // @[Mux.scala 46:19:@12836.4]
  assign _T_14188 = _T_14187 ? _T_10366_39 : _T_14186; // @[Mux.scala 46:16:@12837.4]
  assign _T_14189 = 6'h27 == _T_11317_41; // @[Mux.scala 46:19:@12838.4]
  assign _T_14190 = _T_14189 ? _T_10366_38 : _T_14188; // @[Mux.scala 46:16:@12839.4]
  assign _T_14191 = 6'h26 == _T_11317_41; // @[Mux.scala 46:19:@12840.4]
  assign _T_14192 = _T_14191 ? _T_10366_37 : _T_14190; // @[Mux.scala 46:16:@12841.4]
  assign _T_14193 = 6'h25 == _T_11317_41; // @[Mux.scala 46:19:@12842.4]
  assign _T_14194 = _T_14193 ? _T_10366_36 : _T_14192; // @[Mux.scala 46:16:@12843.4]
  assign _T_14195 = 6'h24 == _T_11317_41; // @[Mux.scala 46:19:@12844.4]
  assign _T_14196 = _T_14195 ? _T_10366_35 : _T_14194; // @[Mux.scala 46:16:@12845.4]
  assign _T_14197 = 6'h23 == _T_11317_41; // @[Mux.scala 46:19:@12846.4]
  assign _T_14198 = _T_14197 ? _T_10366_34 : _T_14196; // @[Mux.scala 46:16:@12847.4]
  assign _T_14199 = 6'h22 == _T_11317_41; // @[Mux.scala 46:19:@12848.4]
  assign _T_14200 = _T_14199 ? _T_10366_33 : _T_14198; // @[Mux.scala 46:16:@12849.4]
  assign _T_14201 = 6'h21 == _T_11317_41; // @[Mux.scala 46:19:@12850.4]
  assign _T_14202 = _T_14201 ? _T_10366_32 : _T_14200; // @[Mux.scala 46:16:@12851.4]
  assign _T_14203 = 6'h20 == _T_11317_41; // @[Mux.scala 46:19:@12852.4]
  assign _T_14204 = _T_14203 ? _T_10366_31 : _T_14202; // @[Mux.scala 46:16:@12853.4]
  assign _T_14205 = 6'h1f == _T_11317_41; // @[Mux.scala 46:19:@12854.4]
  assign _T_14206 = _T_14205 ? _T_10366_30 : _T_14204; // @[Mux.scala 46:16:@12855.4]
  assign _T_14207 = 6'h1e == _T_11317_41; // @[Mux.scala 46:19:@12856.4]
  assign _T_14208 = _T_14207 ? _T_10366_29 : _T_14206; // @[Mux.scala 46:16:@12857.4]
  assign _T_14209 = 6'h1d == _T_11317_41; // @[Mux.scala 46:19:@12858.4]
  assign _T_14210 = _T_14209 ? _T_10366_28 : _T_14208; // @[Mux.scala 46:16:@12859.4]
  assign _T_14211 = 6'h1c == _T_11317_41; // @[Mux.scala 46:19:@12860.4]
  assign _T_14212 = _T_14211 ? _T_10366_27 : _T_14210; // @[Mux.scala 46:16:@12861.4]
  assign _T_14213 = 6'h1b == _T_11317_41; // @[Mux.scala 46:19:@12862.4]
  assign _T_14214 = _T_14213 ? _T_10366_26 : _T_14212; // @[Mux.scala 46:16:@12863.4]
  assign _T_14215 = 6'h1a == _T_11317_41; // @[Mux.scala 46:19:@12864.4]
  assign _T_14216 = _T_14215 ? _T_10366_25 : _T_14214; // @[Mux.scala 46:16:@12865.4]
  assign _T_14217 = 6'h19 == _T_11317_41; // @[Mux.scala 46:19:@12866.4]
  assign _T_14218 = _T_14217 ? _T_10366_24 : _T_14216; // @[Mux.scala 46:16:@12867.4]
  assign _T_14219 = 6'h18 == _T_11317_41; // @[Mux.scala 46:19:@12868.4]
  assign _T_14220 = _T_14219 ? _T_10366_23 : _T_14218; // @[Mux.scala 46:16:@12869.4]
  assign _T_14221 = 6'h17 == _T_11317_41; // @[Mux.scala 46:19:@12870.4]
  assign _T_14222 = _T_14221 ? _T_10366_22 : _T_14220; // @[Mux.scala 46:16:@12871.4]
  assign _T_14223 = 6'h16 == _T_11317_41; // @[Mux.scala 46:19:@12872.4]
  assign _T_14224 = _T_14223 ? _T_10366_21 : _T_14222; // @[Mux.scala 46:16:@12873.4]
  assign _T_14225 = 6'h15 == _T_11317_41; // @[Mux.scala 46:19:@12874.4]
  assign _T_14226 = _T_14225 ? _T_10366_20 : _T_14224; // @[Mux.scala 46:16:@12875.4]
  assign _T_14227 = 6'h14 == _T_11317_41; // @[Mux.scala 46:19:@12876.4]
  assign _T_14228 = _T_14227 ? _T_10366_19 : _T_14226; // @[Mux.scala 46:16:@12877.4]
  assign _T_14229 = 6'h13 == _T_11317_41; // @[Mux.scala 46:19:@12878.4]
  assign _T_14230 = _T_14229 ? _T_10366_18 : _T_14228; // @[Mux.scala 46:16:@12879.4]
  assign _T_14231 = 6'h12 == _T_11317_41; // @[Mux.scala 46:19:@12880.4]
  assign _T_14232 = _T_14231 ? _T_10366_17 : _T_14230; // @[Mux.scala 46:16:@12881.4]
  assign _T_14233 = 6'h11 == _T_11317_41; // @[Mux.scala 46:19:@12882.4]
  assign _T_14234 = _T_14233 ? _T_10366_16 : _T_14232; // @[Mux.scala 46:16:@12883.4]
  assign _T_14235 = 6'h10 == _T_11317_41; // @[Mux.scala 46:19:@12884.4]
  assign _T_14236 = _T_14235 ? _T_10366_15 : _T_14234; // @[Mux.scala 46:16:@12885.4]
  assign _T_14237 = 6'hf == _T_11317_41; // @[Mux.scala 46:19:@12886.4]
  assign _T_14238 = _T_14237 ? _T_10366_14 : _T_14236; // @[Mux.scala 46:16:@12887.4]
  assign _T_14239 = 6'he == _T_11317_41; // @[Mux.scala 46:19:@12888.4]
  assign _T_14240 = _T_14239 ? _T_10366_13 : _T_14238; // @[Mux.scala 46:16:@12889.4]
  assign _T_14241 = 6'hd == _T_11317_41; // @[Mux.scala 46:19:@12890.4]
  assign _T_14242 = _T_14241 ? _T_10366_12 : _T_14240; // @[Mux.scala 46:16:@12891.4]
  assign _T_14243 = 6'hc == _T_11317_41; // @[Mux.scala 46:19:@12892.4]
  assign _T_14244 = _T_14243 ? _T_10366_11 : _T_14242; // @[Mux.scala 46:16:@12893.4]
  assign _T_14245 = 6'hb == _T_11317_41; // @[Mux.scala 46:19:@12894.4]
  assign _T_14246 = _T_14245 ? _T_10366_10 : _T_14244; // @[Mux.scala 46:16:@12895.4]
  assign _T_14247 = 6'ha == _T_11317_41; // @[Mux.scala 46:19:@12896.4]
  assign _T_14248 = _T_14247 ? _T_10366_9 : _T_14246; // @[Mux.scala 46:16:@12897.4]
  assign _T_14249 = 6'h9 == _T_11317_41; // @[Mux.scala 46:19:@12898.4]
  assign _T_14250 = _T_14249 ? _T_10366_8 : _T_14248; // @[Mux.scala 46:16:@12899.4]
  assign _T_14251 = 6'h8 == _T_11317_41; // @[Mux.scala 46:19:@12900.4]
  assign _T_14252 = _T_14251 ? _T_10366_7 : _T_14250; // @[Mux.scala 46:16:@12901.4]
  assign _T_14253 = 6'h7 == _T_11317_41; // @[Mux.scala 46:19:@12902.4]
  assign _T_14254 = _T_14253 ? _T_10366_6 : _T_14252; // @[Mux.scala 46:16:@12903.4]
  assign _T_14255 = 6'h6 == _T_11317_41; // @[Mux.scala 46:19:@12904.4]
  assign _T_14256 = _T_14255 ? _T_10366_5 : _T_14254; // @[Mux.scala 46:16:@12905.4]
  assign _T_14257 = 6'h5 == _T_11317_41; // @[Mux.scala 46:19:@12906.4]
  assign _T_14258 = _T_14257 ? _T_10366_4 : _T_14256; // @[Mux.scala 46:16:@12907.4]
  assign _T_14259 = 6'h4 == _T_11317_41; // @[Mux.scala 46:19:@12908.4]
  assign _T_14260 = _T_14259 ? _T_10366_3 : _T_14258; // @[Mux.scala 46:16:@12909.4]
  assign _T_14261 = 6'h3 == _T_11317_41; // @[Mux.scala 46:19:@12910.4]
  assign _T_14262 = _T_14261 ? _T_10366_2 : _T_14260; // @[Mux.scala 46:16:@12911.4]
  assign _T_14263 = 6'h2 == _T_11317_41; // @[Mux.scala 46:19:@12912.4]
  assign _T_14264 = _T_14263 ? _T_10366_1 : _T_14262; // @[Mux.scala 46:16:@12913.4]
  assign _T_14265 = 6'h1 == _T_11317_41; // @[Mux.scala 46:19:@12914.4]
  assign _T_14266 = _T_14265 ? _T_10366_0 : _T_14264; // @[Mux.scala 46:16:@12915.4]
  assign _T_14311 = 6'h2b == _T_11317_42; // @[Mux.scala 46:19:@12917.4]
  assign _T_14312 = _T_14311 ? _T_10366_42 : 8'h0; // @[Mux.scala 46:16:@12918.4]
  assign _T_14313 = 6'h2a == _T_11317_42; // @[Mux.scala 46:19:@12919.4]
  assign _T_14314 = _T_14313 ? _T_10366_41 : _T_14312; // @[Mux.scala 46:16:@12920.4]
  assign _T_14315 = 6'h29 == _T_11317_42; // @[Mux.scala 46:19:@12921.4]
  assign _T_14316 = _T_14315 ? _T_10366_40 : _T_14314; // @[Mux.scala 46:16:@12922.4]
  assign _T_14317 = 6'h28 == _T_11317_42; // @[Mux.scala 46:19:@12923.4]
  assign _T_14318 = _T_14317 ? _T_10366_39 : _T_14316; // @[Mux.scala 46:16:@12924.4]
  assign _T_14319 = 6'h27 == _T_11317_42; // @[Mux.scala 46:19:@12925.4]
  assign _T_14320 = _T_14319 ? _T_10366_38 : _T_14318; // @[Mux.scala 46:16:@12926.4]
  assign _T_14321 = 6'h26 == _T_11317_42; // @[Mux.scala 46:19:@12927.4]
  assign _T_14322 = _T_14321 ? _T_10366_37 : _T_14320; // @[Mux.scala 46:16:@12928.4]
  assign _T_14323 = 6'h25 == _T_11317_42; // @[Mux.scala 46:19:@12929.4]
  assign _T_14324 = _T_14323 ? _T_10366_36 : _T_14322; // @[Mux.scala 46:16:@12930.4]
  assign _T_14325 = 6'h24 == _T_11317_42; // @[Mux.scala 46:19:@12931.4]
  assign _T_14326 = _T_14325 ? _T_10366_35 : _T_14324; // @[Mux.scala 46:16:@12932.4]
  assign _T_14327 = 6'h23 == _T_11317_42; // @[Mux.scala 46:19:@12933.4]
  assign _T_14328 = _T_14327 ? _T_10366_34 : _T_14326; // @[Mux.scala 46:16:@12934.4]
  assign _T_14329 = 6'h22 == _T_11317_42; // @[Mux.scala 46:19:@12935.4]
  assign _T_14330 = _T_14329 ? _T_10366_33 : _T_14328; // @[Mux.scala 46:16:@12936.4]
  assign _T_14331 = 6'h21 == _T_11317_42; // @[Mux.scala 46:19:@12937.4]
  assign _T_14332 = _T_14331 ? _T_10366_32 : _T_14330; // @[Mux.scala 46:16:@12938.4]
  assign _T_14333 = 6'h20 == _T_11317_42; // @[Mux.scala 46:19:@12939.4]
  assign _T_14334 = _T_14333 ? _T_10366_31 : _T_14332; // @[Mux.scala 46:16:@12940.4]
  assign _T_14335 = 6'h1f == _T_11317_42; // @[Mux.scala 46:19:@12941.4]
  assign _T_14336 = _T_14335 ? _T_10366_30 : _T_14334; // @[Mux.scala 46:16:@12942.4]
  assign _T_14337 = 6'h1e == _T_11317_42; // @[Mux.scala 46:19:@12943.4]
  assign _T_14338 = _T_14337 ? _T_10366_29 : _T_14336; // @[Mux.scala 46:16:@12944.4]
  assign _T_14339 = 6'h1d == _T_11317_42; // @[Mux.scala 46:19:@12945.4]
  assign _T_14340 = _T_14339 ? _T_10366_28 : _T_14338; // @[Mux.scala 46:16:@12946.4]
  assign _T_14341 = 6'h1c == _T_11317_42; // @[Mux.scala 46:19:@12947.4]
  assign _T_14342 = _T_14341 ? _T_10366_27 : _T_14340; // @[Mux.scala 46:16:@12948.4]
  assign _T_14343 = 6'h1b == _T_11317_42; // @[Mux.scala 46:19:@12949.4]
  assign _T_14344 = _T_14343 ? _T_10366_26 : _T_14342; // @[Mux.scala 46:16:@12950.4]
  assign _T_14345 = 6'h1a == _T_11317_42; // @[Mux.scala 46:19:@12951.4]
  assign _T_14346 = _T_14345 ? _T_10366_25 : _T_14344; // @[Mux.scala 46:16:@12952.4]
  assign _T_14347 = 6'h19 == _T_11317_42; // @[Mux.scala 46:19:@12953.4]
  assign _T_14348 = _T_14347 ? _T_10366_24 : _T_14346; // @[Mux.scala 46:16:@12954.4]
  assign _T_14349 = 6'h18 == _T_11317_42; // @[Mux.scala 46:19:@12955.4]
  assign _T_14350 = _T_14349 ? _T_10366_23 : _T_14348; // @[Mux.scala 46:16:@12956.4]
  assign _T_14351 = 6'h17 == _T_11317_42; // @[Mux.scala 46:19:@12957.4]
  assign _T_14352 = _T_14351 ? _T_10366_22 : _T_14350; // @[Mux.scala 46:16:@12958.4]
  assign _T_14353 = 6'h16 == _T_11317_42; // @[Mux.scala 46:19:@12959.4]
  assign _T_14354 = _T_14353 ? _T_10366_21 : _T_14352; // @[Mux.scala 46:16:@12960.4]
  assign _T_14355 = 6'h15 == _T_11317_42; // @[Mux.scala 46:19:@12961.4]
  assign _T_14356 = _T_14355 ? _T_10366_20 : _T_14354; // @[Mux.scala 46:16:@12962.4]
  assign _T_14357 = 6'h14 == _T_11317_42; // @[Mux.scala 46:19:@12963.4]
  assign _T_14358 = _T_14357 ? _T_10366_19 : _T_14356; // @[Mux.scala 46:16:@12964.4]
  assign _T_14359 = 6'h13 == _T_11317_42; // @[Mux.scala 46:19:@12965.4]
  assign _T_14360 = _T_14359 ? _T_10366_18 : _T_14358; // @[Mux.scala 46:16:@12966.4]
  assign _T_14361 = 6'h12 == _T_11317_42; // @[Mux.scala 46:19:@12967.4]
  assign _T_14362 = _T_14361 ? _T_10366_17 : _T_14360; // @[Mux.scala 46:16:@12968.4]
  assign _T_14363 = 6'h11 == _T_11317_42; // @[Mux.scala 46:19:@12969.4]
  assign _T_14364 = _T_14363 ? _T_10366_16 : _T_14362; // @[Mux.scala 46:16:@12970.4]
  assign _T_14365 = 6'h10 == _T_11317_42; // @[Mux.scala 46:19:@12971.4]
  assign _T_14366 = _T_14365 ? _T_10366_15 : _T_14364; // @[Mux.scala 46:16:@12972.4]
  assign _T_14367 = 6'hf == _T_11317_42; // @[Mux.scala 46:19:@12973.4]
  assign _T_14368 = _T_14367 ? _T_10366_14 : _T_14366; // @[Mux.scala 46:16:@12974.4]
  assign _T_14369 = 6'he == _T_11317_42; // @[Mux.scala 46:19:@12975.4]
  assign _T_14370 = _T_14369 ? _T_10366_13 : _T_14368; // @[Mux.scala 46:16:@12976.4]
  assign _T_14371 = 6'hd == _T_11317_42; // @[Mux.scala 46:19:@12977.4]
  assign _T_14372 = _T_14371 ? _T_10366_12 : _T_14370; // @[Mux.scala 46:16:@12978.4]
  assign _T_14373 = 6'hc == _T_11317_42; // @[Mux.scala 46:19:@12979.4]
  assign _T_14374 = _T_14373 ? _T_10366_11 : _T_14372; // @[Mux.scala 46:16:@12980.4]
  assign _T_14375 = 6'hb == _T_11317_42; // @[Mux.scala 46:19:@12981.4]
  assign _T_14376 = _T_14375 ? _T_10366_10 : _T_14374; // @[Mux.scala 46:16:@12982.4]
  assign _T_14377 = 6'ha == _T_11317_42; // @[Mux.scala 46:19:@12983.4]
  assign _T_14378 = _T_14377 ? _T_10366_9 : _T_14376; // @[Mux.scala 46:16:@12984.4]
  assign _T_14379 = 6'h9 == _T_11317_42; // @[Mux.scala 46:19:@12985.4]
  assign _T_14380 = _T_14379 ? _T_10366_8 : _T_14378; // @[Mux.scala 46:16:@12986.4]
  assign _T_14381 = 6'h8 == _T_11317_42; // @[Mux.scala 46:19:@12987.4]
  assign _T_14382 = _T_14381 ? _T_10366_7 : _T_14380; // @[Mux.scala 46:16:@12988.4]
  assign _T_14383 = 6'h7 == _T_11317_42; // @[Mux.scala 46:19:@12989.4]
  assign _T_14384 = _T_14383 ? _T_10366_6 : _T_14382; // @[Mux.scala 46:16:@12990.4]
  assign _T_14385 = 6'h6 == _T_11317_42; // @[Mux.scala 46:19:@12991.4]
  assign _T_14386 = _T_14385 ? _T_10366_5 : _T_14384; // @[Mux.scala 46:16:@12992.4]
  assign _T_14387 = 6'h5 == _T_11317_42; // @[Mux.scala 46:19:@12993.4]
  assign _T_14388 = _T_14387 ? _T_10366_4 : _T_14386; // @[Mux.scala 46:16:@12994.4]
  assign _T_14389 = 6'h4 == _T_11317_42; // @[Mux.scala 46:19:@12995.4]
  assign _T_14390 = _T_14389 ? _T_10366_3 : _T_14388; // @[Mux.scala 46:16:@12996.4]
  assign _T_14391 = 6'h3 == _T_11317_42; // @[Mux.scala 46:19:@12997.4]
  assign _T_14392 = _T_14391 ? _T_10366_2 : _T_14390; // @[Mux.scala 46:16:@12998.4]
  assign _T_14393 = 6'h2 == _T_11317_42; // @[Mux.scala 46:19:@12999.4]
  assign _T_14394 = _T_14393 ? _T_10366_1 : _T_14392; // @[Mux.scala 46:16:@13000.4]
  assign _T_14395 = 6'h1 == _T_11317_42; // @[Mux.scala 46:19:@13001.4]
  assign _T_14396 = _T_14395 ? _T_10366_0 : _T_14394; // @[Mux.scala 46:16:@13002.4]
  assign _T_14442 = 6'h2c == _T_11317_43; // @[Mux.scala 46:19:@13004.4]
  assign _T_14443 = _T_14442 ? _T_10366_43 : 8'h0; // @[Mux.scala 46:16:@13005.4]
  assign _T_14444 = 6'h2b == _T_11317_43; // @[Mux.scala 46:19:@13006.4]
  assign _T_14445 = _T_14444 ? _T_10366_42 : _T_14443; // @[Mux.scala 46:16:@13007.4]
  assign _T_14446 = 6'h2a == _T_11317_43; // @[Mux.scala 46:19:@13008.4]
  assign _T_14447 = _T_14446 ? _T_10366_41 : _T_14445; // @[Mux.scala 46:16:@13009.4]
  assign _T_14448 = 6'h29 == _T_11317_43; // @[Mux.scala 46:19:@13010.4]
  assign _T_14449 = _T_14448 ? _T_10366_40 : _T_14447; // @[Mux.scala 46:16:@13011.4]
  assign _T_14450 = 6'h28 == _T_11317_43; // @[Mux.scala 46:19:@13012.4]
  assign _T_14451 = _T_14450 ? _T_10366_39 : _T_14449; // @[Mux.scala 46:16:@13013.4]
  assign _T_14452 = 6'h27 == _T_11317_43; // @[Mux.scala 46:19:@13014.4]
  assign _T_14453 = _T_14452 ? _T_10366_38 : _T_14451; // @[Mux.scala 46:16:@13015.4]
  assign _T_14454 = 6'h26 == _T_11317_43; // @[Mux.scala 46:19:@13016.4]
  assign _T_14455 = _T_14454 ? _T_10366_37 : _T_14453; // @[Mux.scala 46:16:@13017.4]
  assign _T_14456 = 6'h25 == _T_11317_43; // @[Mux.scala 46:19:@13018.4]
  assign _T_14457 = _T_14456 ? _T_10366_36 : _T_14455; // @[Mux.scala 46:16:@13019.4]
  assign _T_14458 = 6'h24 == _T_11317_43; // @[Mux.scala 46:19:@13020.4]
  assign _T_14459 = _T_14458 ? _T_10366_35 : _T_14457; // @[Mux.scala 46:16:@13021.4]
  assign _T_14460 = 6'h23 == _T_11317_43; // @[Mux.scala 46:19:@13022.4]
  assign _T_14461 = _T_14460 ? _T_10366_34 : _T_14459; // @[Mux.scala 46:16:@13023.4]
  assign _T_14462 = 6'h22 == _T_11317_43; // @[Mux.scala 46:19:@13024.4]
  assign _T_14463 = _T_14462 ? _T_10366_33 : _T_14461; // @[Mux.scala 46:16:@13025.4]
  assign _T_14464 = 6'h21 == _T_11317_43; // @[Mux.scala 46:19:@13026.4]
  assign _T_14465 = _T_14464 ? _T_10366_32 : _T_14463; // @[Mux.scala 46:16:@13027.4]
  assign _T_14466 = 6'h20 == _T_11317_43; // @[Mux.scala 46:19:@13028.4]
  assign _T_14467 = _T_14466 ? _T_10366_31 : _T_14465; // @[Mux.scala 46:16:@13029.4]
  assign _T_14468 = 6'h1f == _T_11317_43; // @[Mux.scala 46:19:@13030.4]
  assign _T_14469 = _T_14468 ? _T_10366_30 : _T_14467; // @[Mux.scala 46:16:@13031.4]
  assign _T_14470 = 6'h1e == _T_11317_43; // @[Mux.scala 46:19:@13032.4]
  assign _T_14471 = _T_14470 ? _T_10366_29 : _T_14469; // @[Mux.scala 46:16:@13033.4]
  assign _T_14472 = 6'h1d == _T_11317_43; // @[Mux.scala 46:19:@13034.4]
  assign _T_14473 = _T_14472 ? _T_10366_28 : _T_14471; // @[Mux.scala 46:16:@13035.4]
  assign _T_14474 = 6'h1c == _T_11317_43; // @[Mux.scala 46:19:@13036.4]
  assign _T_14475 = _T_14474 ? _T_10366_27 : _T_14473; // @[Mux.scala 46:16:@13037.4]
  assign _T_14476 = 6'h1b == _T_11317_43; // @[Mux.scala 46:19:@13038.4]
  assign _T_14477 = _T_14476 ? _T_10366_26 : _T_14475; // @[Mux.scala 46:16:@13039.4]
  assign _T_14478 = 6'h1a == _T_11317_43; // @[Mux.scala 46:19:@13040.4]
  assign _T_14479 = _T_14478 ? _T_10366_25 : _T_14477; // @[Mux.scala 46:16:@13041.4]
  assign _T_14480 = 6'h19 == _T_11317_43; // @[Mux.scala 46:19:@13042.4]
  assign _T_14481 = _T_14480 ? _T_10366_24 : _T_14479; // @[Mux.scala 46:16:@13043.4]
  assign _T_14482 = 6'h18 == _T_11317_43; // @[Mux.scala 46:19:@13044.4]
  assign _T_14483 = _T_14482 ? _T_10366_23 : _T_14481; // @[Mux.scala 46:16:@13045.4]
  assign _T_14484 = 6'h17 == _T_11317_43; // @[Mux.scala 46:19:@13046.4]
  assign _T_14485 = _T_14484 ? _T_10366_22 : _T_14483; // @[Mux.scala 46:16:@13047.4]
  assign _T_14486 = 6'h16 == _T_11317_43; // @[Mux.scala 46:19:@13048.4]
  assign _T_14487 = _T_14486 ? _T_10366_21 : _T_14485; // @[Mux.scala 46:16:@13049.4]
  assign _T_14488 = 6'h15 == _T_11317_43; // @[Mux.scala 46:19:@13050.4]
  assign _T_14489 = _T_14488 ? _T_10366_20 : _T_14487; // @[Mux.scala 46:16:@13051.4]
  assign _T_14490 = 6'h14 == _T_11317_43; // @[Mux.scala 46:19:@13052.4]
  assign _T_14491 = _T_14490 ? _T_10366_19 : _T_14489; // @[Mux.scala 46:16:@13053.4]
  assign _T_14492 = 6'h13 == _T_11317_43; // @[Mux.scala 46:19:@13054.4]
  assign _T_14493 = _T_14492 ? _T_10366_18 : _T_14491; // @[Mux.scala 46:16:@13055.4]
  assign _T_14494 = 6'h12 == _T_11317_43; // @[Mux.scala 46:19:@13056.4]
  assign _T_14495 = _T_14494 ? _T_10366_17 : _T_14493; // @[Mux.scala 46:16:@13057.4]
  assign _T_14496 = 6'h11 == _T_11317_43; // @[Mux.scala 46:19:@13058.4]
  assign _T_14497 = _T_14496 ? _T_10366_16 : _T_14495; // @[Mux.scala 46:16:@13059.4]
  assign _T_14498 = 6'h10 == _T_11317_43; // @[Mux.scala 46:19:@13060.4]
  assign _T_14499 = _T_14498 ? _T_10366_15 : _T_14497; // @[Mux.scala 46:16:@13061.4]
  assign _T_14500 = 6'hf == _T_11317_43; // @[Mux.scala 46:19:@13062.4]
  assign _T_14501 = _T_14500 ? _T_10366_14 : _T_14499; // @[Mux.scala 46:16:@13063.4]
  assign _T_14502 = 6'he == _T_11317_43; // @[Mux.scala 46:19:@13064.4]
  assign _T_14503 = _T_14502 ? _T_10366_13 : _T_14501; // @[Mux.scala 46:16:@13065.4]
  assign _T_14504 = 6'hd == _T_11317_43; // @[Mux.scala 46:19:@13066.4]
  assign _T_14505 = _T_14504 ? _T_10366_12 : _T_14503; // @[Mux.scala 46:16:@13067.4]
  assign _T_14506 = 6'hc == _T_11317_43; // @[Mux.scala 46:19:@13068.4]
  assign _T_14507 = _T_14506 ? _T_10366_11 : _T_14505; // @[Mux.scala 46:16:@13069.4]
  assign _T_14508 = 6'hb == _T_11317_43; // @[Mux.scala 46:19:@13070.4]
  assign _T_14509 = _T_14508 ? _T_10366_10 : _T_14507; // @[Mux.scala 46:16:@13071.4]
  assign _T_14510 = 6'ha == _T_11317_43; // @[Mux.scala 46:19:@13072.4]
  assign _T_14511 = _T_14510 ? _T_10366_9 : _T_14509; // @[Mux.scala 46:16:@13073.4]
  assign _T_14512 = 6'h9 == _T_11317_43; // @[Mux.scala 46:19:@13074.4]
  assign _T_14513 = _T_14512 ? _T_10366_8 : _T_14511; // @[Mux.scala 46:16:@13075.4]
  assign _T_14514 = 6'h8 == _T_11317_43; // @[Mux.scala 46:19:@13076.4]
  assign _T_14515 = _T_14514 ? _T_10366_7 : _T_14513; // @[Mux.scala 46:16:@13077.4]
  assign _T_14516 = 6'h7 == _T_11317_43; // @[Mux.scala 46:19:@13078.4]
  assign _T_14517 = _T_14516 ? _T_10366_6 : _T_14515; // @[Mux.scala 46:16:@13079.4]
  assign _T_14518 = 6'h6 == _T_11317_43; // @[Mux.scala 46:19:@13080.4]
  assign _T_14519 = _T_14518 ? _T_10366_5 : _T_14517; // @[Mux.scala 46:16:@13081.4]
  assign _T_14520 = 6'h5 == _T_11317_43; // @[Mux.scala 46:19:@13082.4]
  assign _T_14521 = _T_14520 ? _T_10366_4 : _T_14519; // @[Mux.scala 46:16:@13083.4]
  assign _T_14522 = 6'h4 == _T_11317_43; // @[Mux.scala 46:19:@13084.4]
  assign _T_14523 = _T_14522 ? _T_10366_3 : _T_14521; // @[Mux.scala 46:16:@13085.4]
  assign _T_14524 = 6'h3 == _T_11317_43; // @[Mux.scala 46:19:@13086.4]
  assign _T_14525 = _T_14524 ? _T_10366_2 : _T_14523; // @[Mux.scala 46:16:@13087.4]
  assign _T_14526 = 6'h2 == _T_11317_43; // @[Mux.scala 46:19:@13088.4]
  assign _T_14527 = _T_14526 ? _T_10366_1 : _T_14525; // @[Mux.scala 46:16:@13089.4]
  assign _T_14528 = 6'h1 == _T_11317_43; // @[Mux.scala 46:19:@13090.4]
  assign _T_14529 = _T_14528 ? _T_10366_0 : _T_14527; // @[Mux.scala 46:16:@13091.4]
  assign _T_14576 = 6'h2d == _T_11317_44; // @[Mux.scala 46:19:@13093.4]
  assign _T_14577 = _T_14576 ? _T_10366_44 : 8'h0; // @[Mux.scala 46:16:@13094.4]
  assign _T_14578 = 6'h2c == _T_11317_44; // @[Mux.scala 46:19:@13095.4]
  assign _T_14579 = _T_14578 ? _T_10366_43 : _T_14577; // @[Mux.scala 46:16:@13096.4]
  assign _T_14580 = 6'h2b == _T_11317_44; // @[Mux.scala 46:19:@13097.4]
  assign _T_14581 = _T_14580 ? _T_10366_42 : _T_14579; // @[Mux.scala 46:16:@13098.4]
  assign _T_14582 = 6'h2a == _T_11317_44; // @[Mux.scala 46:19:@13099.4]
  assign _T_14583 = _T_14582 ? _T_10366_41 : _T_14581; // @[Mux.scala 46:16:@13100.4]
  assign _T_14584 = 6'h29 == _T_11317_44; // @[Mux.scala 46:19:@13101.4]
  assign _T_14585 = _T_14584 ? _T_10366_40 : _T_14583; // @[Mux.scala 46:16:@13102.4]
  assign _T_14586 = 6'h28 == _T_11317_44; // @[Mux.scala 46:19:@13103.4]
  assign _T_14587 = _T_14586 ? _T_10366_39 : _T_14585; // @[Mux.scala 46:16:@13104.4]
  assign _T_14588 = 6'h27 == _T_11317_44; // @[Mux.scala 46:19:@13105.4]
  assign _T_14589 = _T_14588 ? _T_10366_38 : _T_14587; // @[Mux.scala 46:16:@13106.4]
  assign _T_14590 = 6'h26 == _T_11317_44; // @[Mux.scala 46:19:@13107.4]
  assign _T_14591 = _T_14590 ? _T_10366_37 : _T_14589; // @[Mux.scala 46:16:@13108.4]
  assign _T_14592 = 6'h25 == _T_11317_44; // @[Mux.scala 46:19:@13109.4]
  assign _T_14593 = _T_14592 ? _T_10366_36 : _T_14591; // @[Mux.scala 46:16:@13110.4]
  assign _T_14594 = 6'h24 == _T_11317_44; // @[Mux.scala 46:19:@13111.4]
  assign _T_14595 = _T_14594 ? _T_10366_35 : _T_14593; // @[Mux.scala 46:16:@13112.4]
  assign _T_14596 = 6'h23 == _T_11317_44; // @[Mux.scala 46:19:@13113.4]
  assign _T_14597 = _T_14596 ? _T_10366_34 : _T_14595; // @[Mux.scala 46:16:@13114.4]
  assign _T_14598 = 6'h22 == _T_11317_44; // @[Mux.scala 46:19:@13115.4]
  assign _T_14599 = _T_14598 ? _T_10366_33 : _T_14597; // @[Mux.scala 46:16:@13116.4]
  assign _T_14600 = 6'h21 == _T_11317_44; // @[Mux.scala 46:19:@13117.4]
  assign _T_14601 = _T_14600 ? _T_10366_32 : _T_14599; // @[Mux.scala 46:16:@13118.4]
  assign _T_14602 = 6'h20 == _T_11317_44; // @[Mux.scala 46:19:@13119.4]
  assign _T_14603 = _T_14602 ? _T_10366_31 : _T_14601; // @[Mux.scala 46:16:@13120.4]
  assign _T_14604 = 6'h1f == _T_11317_44; // @[Mux.scala 46:19:@13121.4]
  assign _T_14605 = _T_14604 ? _T_10366_30 : _T_14603; // @[Mux.scala 46:16:@13122.4]
  assign _T_14606 = 6'h1e == _T_11317_44; // @[Mux.scala 46:19:@13123.4]
  assign _T_14607 = _T_14606 ? _T_10366_29 : _T_14605; // @[Mux.scala 46:16:@13124.4]
  assign _T_14608 = 6'h1d == _T_11317_44; // @[Mux.scala 46:19:@13125.4]
  assign _T_14609 = _T_14608 ? _T_10366_28 : _T_14607; // @[Mux.scala 46:16:@13126.4]
  assign _T_14610 = 6'h1c == _T_11317_44; // @[Mux.scala 46:19:@13127.4]
  assign _T_14611 = _T_14610 ? _T_10366_27 : _T_14609; // @[Mux.scala 46:16:@13128.4]
  assign _T_14612 = 6'h1b == _T_11317_44; // @[Mux.scala 46:19:@13129.4]
  assign _T_14613 = _T_14612 ? _T_10366_26 : _T_14611; // @[Mux.scala 46:16:@13130.4]
  assign _T_14614 = 6'h1a == _T_11317_44; // @[Mux.scala 46:19:@13131.4]
  assign _T_14615 = _T_14614 ? _T_10366_25 : _T_14613; // @[Mux.scala 46:16:@13132.4]
  assign _T_14616 = 6'h19 == _T_11317_44; // @[Mux.scala 46:19:@13133.4]
  assign _T_14617 = _T_14616 ? _T_10366_24 : _T_14615; // @[Mux.scala 46:16:@13134.4]
  assign _T_14618 = 6'h18 == _T_11317_44; // @[Mux.scala 46:19:@13135.4]
  assign _T_14619 = _T_14618 ? _T_10366_23 : _T_14617; // @[Mux.scala 46:16:@13136.4]
  assign _T_14620 = 6'h17 == _T_11317_44; // @[Mux.scala 46:19:@13137.4]
  assign _T_14621 = _T_14620 ? _T_10366_22 : _T_14619; // @[Mux.scala 46:16:@13138.4]
  assign _T_14622 = 6'h16 == _T_11317_44; // @[Mux.scala 46:19:@13139.4]
  assign _T_14623 = _T_14622 ? _T_10366_21 : _T_14621; // @[Mux.scala 46:16:@13140.4]
  assign _T_14624 = 6'h15 == _T_11317_44; // @[Mux.scala 46:19:@13141.4]
  assign _T_14625 = _T_14624 ? _T_10366_20 : _T_14623; // @[Mux.scala 46:16:@13142.4]
  assign _T_14626 = 6'h14 == _T_11317_44; // @[Mux.scala 46:19:@13143.4]
  assign _T_14627 = _T_14626 ? _T_10366_19 : _T_14625; // @[Mux.scala 46:16:@13144.4]
  assign _T_14628 = 6'h13 == _T_11317_44; // @[Mux.scala 46:19:@13145.4]
  assign _T_14629 = _T_14628 ? _T_10366_18 : _T_14627; // @[Mux.scala 46:16:@13146.4]
  assign _T_14630 = 6'h12 == _T_11317_44; // @[Mux.scala 46:19:@13147.4]
  assign _T_14631 = _T_14630 ? _T_10366_17 : _T_14629; // @[Mux.scala 46:16:@13148.4]
  assign _T_14632 = 6'h11 == _T_11317_44; // @[Mux.scala 46:19:@13149.4]
  assign _T_14633 = _T_14632 ? _T_10366_16 : _T_14631; // @[Mux.scala 46:16:@13150.4]
  assign _T_14634 = 6'h10 == _T_11317_44; // @[Mux.scala 46:19:@13151.4]
  assign _T_14635 = _T_14634 ? _T_10366_15 : _T_14633; // @[Mux.scala 46:16:@13152.4]
  assign _T_14636 = 6'hf == _T_11317_44; // @[Mux.scala 46:19:@13153.4]
  assign _T_14637 = _T_14636 ? _T_10366_14 : _T_14635; // @[Mux.scala 46:16:@13154.4]
  assign _T_14638 = 6'he == _T_11317_44; // @[Mux.scala 46:19:@13155.4]
  assign _T_14639 = _T_14638 ? _T_10366_13 : _T_14637; // @[Mux.scala 46:16:@13156.4]
  assign _T_14640 = 6'hd == _T_11317_44; // @[Mux.scala 46:19:@13157.4]
  assign _T_14641 = _T_14640 ? _T_10366_12 : _T_14639; // @[Mux.scala 46:16:@13158.4]
  assign _T_14642 = 6'hc == _T_11317_44; // @[Mux.scala 46:19:@13159.4]
  assign _T_14643 = _T_14642 ? _T_10366_11 : _T_14641; // @[Mux.scala 46:16:@13160.4]
  assign _T_14644 = 6'hb == _T_11317_44; // @[Mux.scala 46:19:@13161.4]
  assign _T_14645 = _T_14644 ? _T_10366_10 : _T_14643; // @[Mux.scala 46:16:@13162.4]
  assign _T_14646 = 6'ha == _T_11317_44; // @[Mux.scala 46:19:@13163.4]
  assign _T_14647 = _T_14646 ? _T_10366_9 : _T_14645; // @[Mux.scala 46:16:@13164.4]
  assign _T_14648 = 6'h9 == _T_11317_44; // @[Mux.scala 46:19:@13165.4]
  assign _T_14649 = _T_14648 ? _T_10366_8 : _T_14647; // @[Mux.scala 46:16:@13166.4]
  assign _T_14650 = 6'h8 == _T_11317_44; // @[Mux.scala 46:19:@13167.4]
  assign _T_14651 = _T_14650 ? _T_10366_7 : _T_14649; // @[Mux.scala 46:16:@13168.4]
  assign _T_14652 = 6'h7 == _T_11317_44; // @[Mux.scala 46:19:@13169.4]
  assign _T_14653 = _T_14652 ? _T_10366_6 : _T_14651; // @[Mux.scala 46:16:@13170.4]
  assign _T_14654 = 6'h6 == _T_11317_44; // @[Mux.scala 46:19:@13171.4]
  assign _T_14655 = _T_14654 ? _T_10366_5 : _T_14653; // @[Mux.scala 46:16:@13172.4]
  assign _T_14656 = 6'h5 == _T_11317_44; // @[Mux.scala 46:19:@13173.4]
  assign _T_14657 = _T_14656 ? _T_10366_4 : _T_14655; // @[Mux.scala 46:16:@13174.4]
  assign _T_14658 = 6'h4 == _T_11317_44; // @[Mux.scala 46:19:@13175.4]
  assign _T_14659 = _T_14658 ? _T_10366_3 : _T_14657; // @[Mux.scala 46:16:@13176.4]
  assign _T_14660 = 6'h3 == _T_11317_44; // @[Mux.scala 46:19:@13177.4]
  assign _T_14661 = _T_14660 ? _T_10366_2 : _T_14659; // @[Mux.scala 46:16:@13178.4]
  assign _T_14662 = 6'h2 == _T_11317_44; // @[Mux.scala 46:19:@13179.4]
  assign _T_14663 = _T_14662 ? _T_10366_1 : _T_14661; // @[Mux.scala 46:16:@13180.4]
  assign _T_14664 = 6'h1 == _T_11317_44; // @[Mux.scala 46:19:@13181.4]
  assign _T_14665 = _T_14664 ? _T_10366_0 : _T_14663; // @[Mux.scala 46:16:@13182.4]
  assign _T_14713 = 6'h2e == _T_11317_45; // @[Mux.scala 46:19:@13184.4]
  assign _T_14714 = _T_14713 ? _T_10366_45 : 8'h0; // @[Mux.scala 46:16:@13185.4]
  assign _T_14715 = 6'h2d == _T_11317_45; // @[Mux.scala 46:19:@13186.4]
  assign _T_14716 = _T_14715 ? _T_10366_44 : _T_14714; // @[Mux.scala 46:16:@13187.4]
  assign _T_14717 = 6'h2c == _T_11317_45; // @[Mux.scala 46:19:@13188.4]
  assign _T_14718 = _T_14717 ? _T_10366_43 : _T_14716; // @[Mux.scala 46:16:@13189.4]
  assign _T_14719 = 6'h2b == _T_11317_45; // @[Mux.scala 46:19:@13190.4]
  assign _T_14720 = _T_14719 ? _T_10366_42 : _T_14718; // @[Mux.scala 46:16:@13191.4]
  assign _T_14721 = 6'h2a == _T_11317_45; // @[Mux.scala 46:19:@13192.4]
  assign _T_14722 = _T_14721 ? _T_10366_41 : _T_14720; // @[Mux.scala 46:16:@13193.4]
  assign _T_14723 = 6'h29 == _T_11317_45; // @[Mux.scala 46:19:@13194.4]
  assign _T_14724 = _T_14723 ? _T_10366_40 : _T_14722; // @[Mux.scala 46:16:@13195.4]
  assign _T_14725 = 6'h28 == _T_11317_45; // @[Mux.scala 46:19:@13196.4]
  assign _T_14726 = _T_14725 ? _T_10366_39 : _T_14724; // @[Mux.scala 46:16:@13197.4]
  assign _T_14727 = 6'h27 == _T_11317_45; // @[Mux.scala 46:19:@13198.4]
  assign _T_14728 = _T_14727 ? _T_10366_38 : _T_14726; // @[Mux.scala 46:16:@13199.4]
  assign _T_14729 = 6'h26 == _T_11317_45; // @[Mux.scala 46:19:@13200.4]
  assign _T_14730 = _T_14729 ? _T_10366_37 : _T_14728; // @[Mux.scala 46:16:@13201.4]
  assign _T_14731 = 6'h25 == _T_11317_45; // @[Mux.scala 46:19:@13202.4]
  assign _T_14732 = _T_14731 ? _T_10366_36 : _T_14730; // @[Mux.scala 46:16:@13203.4]
  assign _T_14733 = 6'h24 == _T_11317_45; // @[Mux.scala 46:19:@13204.4]
  assign _T_14734 = _T_14733 ? _T_10366_35 : _T_14732; // @[Mux.scala 46:16:@13205.4]
  assign _T_14735 = 6'h23 == _T_11317_45; // @[Mux.scala 46:19:@13206.4]
  assign _T_14736 = _T_14735 ? _T_10366_34 : _T_14734; // @[Mux.scala 46:16:@13207.4]
  assign _T_14737 = 6'h22 == _T_11317_45; // @[Mux.scala 46:19:@13208.4]
  assign _T_14738 = _T_14737 ? _T_10366_33 : _T_14736; // @[Mux.scala 46:16:@13209.4]
  assign _T_14739 = 6'h21 == _T_11317_45; // @[Mux.scala 46:19:@13210.4]
  assign _T_14740 = _T_14739 ? _T_10366_32 : _T_14738; // @[Mux.scala 46:16:@13211.4]
  assign _T_14741 = 6'h20 == _T_11317_45; // @[Mux.scala 46:19:@13212.4]
  assign _T_14742 = _T_14741 ? _T_10366_31 : _T_14740; // @[Mux.scala 46:16:@13213.4]
  assign _T_14743 = 6'h1f == _T_11317_45; // @[Mux.scala 46:19:@13214.4]
  assign _T_14744 = _T_14743 ? _T_10366_30 : _T_14742; // @[Mux.scala 46:16:@13215.4]
  assign _T_14745 = 6'h1e == _T_11317_45; // @[Mux.scala 46:19:@13216.4]
  assign _T_14746 = _T_14745 ? _T_10366_29 : _T_14744; // @[Mux.scala 46:16:@13217.4]
  assign _T_14747 = 6'h1d == _T_11317_45; // @[Mux.scala 46:19:@13218.4]
  assign _T_14748 = _T_14747 ? _T_10366_28 : _T_14746; // @[Mux.scala 46:16:@13219.4]
  assign _T_14749 = 6'h1c == _T_11317_45; // @[Mux.scala 46:19:@13220.4]
  assign _T_14750 = _T_14749 ? _T_10366_27 : _T_14748; // @[Mux.scala 46:16:@13221.4]
  assign _T_14751 = 6'h1b == _T_11317_45; // @[Mux.scala 46:19:@13222.4]
  assign _T_14752 = _T_14751 ? _T_10366_26 : _T_14750; // @[Mux.scala 46:16:@13223.4]
  assign _T_14753 = 6'h1a == _T_11317_45; // @[Mux.scala 46:19:@13224.4]
  assign _T_14754 = _T_14753 ? _T_10366_25 : _T_14752; // @[Mux.scala 46:16:@13225.4]
  assign _T_14755 = 6'h19 == _T_11317_45; // @[Mux.scala 46:19:@13226.4]
  assign _T_14756 = _T_14755 ? _T_10366_24 : _T_14754; // @[Mux.scala 46:16:@13227.4]
  assign _T_14757 = 6'h18 == _T_11317_45; // @[Mux.scala 46:19:@13228.4]
  assign _T_14758 = _T_14757 ? _T_10366_23 : _T_14756; // @[Mux.scala 46:16:@13229.4]
  assign _T_14759 = 6'h17 == _T_11317_45; // @[Mux.scala 46:19:@13230.4]
  assign _T_14760 = _T_14759 ? _T_10366_22 : _T_14758; // @[Mux.scala 46:16:@13231.4]
  assign _T_14761 = 6'h16 == _T_11317_45; // @[Mux.scala 46:19:@13232.4]
  assign _T_14762 = _T_14761 ? _T_10366_21 : _T_14760; // @[Mux.scala 46:16:@13233.4]
  assign _T_14763 = 6'h15 == _T_11317_45; // @[Mux.scala 46:19:@13234.4]
  assign _T_14764 = _T_14763 ? _T_10366_20 : _T_14762; // @[Mux.scala 46:16:@13235.4]
  assign _T_14765 = 6'h14 == _T_11317_45; // @[Mux.scala 46:19:@13236.4]
  assign _T_14766 = _T_14765 ? _T_10366_19 : _T_14764; // @[Mux.scala 46:16:@13237.4]
  assign _T_14767 = 6'h13 == _T_11317_45; // @[Mux.scala 46:19:@13238.4]
  assign _T_14768 = _T_14767 ? _T_10366_18 : _T_14766; // @[Mux.scala 46:16:@13239.4]
  assign _T_14769 = 6'h12 == _T_11317_45; // @[Mux.scala 46:19:@13240.4]
  assign _T_14770 = _T_14769 ? _T_10366_17 : _T_14768; // @[Mux.scala 46:16:@13241.4]
  assign _T_14771 = 6'h11 == _T_11317_45; // @[Mux.scala 46:19:@13242.4]
  assign _T_14772 = _T_14771 ? _T_10366_16 : _T_14770; // @[Mux.scala 46:16:@13243.4]
  assign _T_14773 = 6'h10 == _T_11317_45; // @[Mux.scala 46:19:@13244.4]
  assign _T_14774 = _T_14773 ? _T_10366_15 : _T_14772; // @[Mux.scala 46:16:@13245.4]
  assign _T_14775 = 6'hf == _T_11317_45; // @[Mux.scala 46:19:@13246.4]
  assign _T_14776 = _T_14775 ? _T_10366_14 : _T_14774; // @[Mux.scala 46:16:@13247.4]
  assign _T_14777 = 6'he == _T_11317_45; // @[Mux.scala 46:19:@13248.4]
  assign _T_14778 = _T_14777 ? _T_10366_13 : _T_14776; // @[Mux.scala 46:16:@13249.4]
  assign _T_14779 = 6'hd == _T_11317_45; // @[Mux.scala 46:19:@13250.4]
  assign _T_14780 = _T_14779 ? _T_10366_12 : _T_14778; // @[Mux.scala 46:16:@13251.4]
  assign _T_14781 = 6'hc == _T_11317_45; // @[Mux.scala 46:19:@13252.4]
  assign _T_14782 = _T_14781 ? _T_10366_11 : _T_14780; // @[Mux.scala 46:16:@13253.4]
  assign _T_14783 = 6'hb == _T_11317_45; // @[Mux.scala 46:19:@13254.4]
  assign _T_14784 = _T_14783 ? _T_10366_10 : _T_14782; // @[Mux.scala 46:16:@13255.4]
  assign _T_14785 = 6'ha == _T_11317_45; // @[Mux.scala 46:19:@13256.4]
  assign _T_14786 = _T_14785 ? _T_10366_9 : _T_14784; // @[Mux.scala 46:16:@13257.4]
  assign _T_14787 = 6'h9 == _T_11317_45; // @[Mux.scala 46:19:@13258.4]
  assign _T_14788 = _T_14787 ? _T_10366_8 : _T_14786; // @[Mux.scala 46:16:@13259.4]
  assign _T_14789 = 6'h8 == _T_11317_45; // @[Mux.scala 46:19:@13260.4]
  assign _T_14790 = _T_14789 ? _T_10366_7 : _T_14788; // @[Mux.scala 46:16:@13261.4]
  assign _T_14791 = 6'h7 == _T_11317_45; // @[Mux.scala 46:19:@13262.4]
  assign _T_14792 = _T_14791 ? _T_10366_6 : _T_14790; // @[Mux.scala 46:16:@13263.4]
  assign _T_14793 = 6'h6 == _T_11317_45; // @[Mux.scala 46:19:@13264.4]
  assign _T_14794 = _T_14793 ? _T_10366_5 : _T_14792; // @[Mux.scala 46:16:@13265.4]
  assign _T_14795 = 6'h5 == _T_11317_45; // @[Mux.scala 46:19:@13266.4]
  assign _T_14796 = _T_14795 ? _T_10366_4 : _T_14794; // @[Mux.scala 46:16:@13267.4]
  assign _T_14797 = 6'h4 == _T_11317_45; // @[Mux.scala 46:19:@13268.4]
  assign _T_14798 = _T_14797 ? _T_10366_3 : _T_14796; // @[Mux.scala 46:16:@13269.4]
  assign _T_14799 = 6'h3 == _T_11317_45; // @[Mux.scala 46:19:@13270.4]
  assign _T_14800 = _T_14799 ? _T_10366_2 : _T_14798; // @[Mux.scala 46:16:@13271.4]
  assign _T_14801 = 6'h2 == _T_11317_45; // @[Mux.scala 46:19:@13272.4]
  assign _T_14802 = _T_14801 ? _T_10366_1 : _T_14800; // @[Mux.scala 46:16:@13273.4]
  assign _T_14803 = 6'h1 == _T_11317_45; // @[Mux.scala 46:19:@13274.4]
  assign _T_14804 = _T_14803 ? _T_10366_0 : _T_14802; // @[Mux.scala 46:16:@13275.4]
  assign _T_14853 = 6'h2f == _T_11317_46; // @[Mux.scala 46:19:@13277.4]
  assign _T_14854 = _T_14853 ? _T_10366_46 : 8'h0; // @[Mux.scala 46:16:@13278.4]
  assign _T_14855 = 6'h2e == _T_11317_46; // @[Mux.scala 46:19:@13279.4]
  assign _T_14856 = _T_14855 ? _T_10366_45 : _T_14854; // @[Mux.scala 46:16:@13280.4]
  assign _T_14857 = 6'h2d == _T_11317_46; // @[Mux.scala 46:19:@13281.4]
  assign _T_14858 = _T_14857 ? _T_10366_44 : _T_14856; // @[Mux.scala 46:16:@13282.4]
  assign _T_14859 = 6'h2c == _T_11317_46; // @[Mux.scala 46:19:@13283.4]
  assign _T_14860 = _T_14859 ? _T_10366_43 : _T_14858; // @[Mux.scala 46:16:@13284.4]
  assign _T_14861 = 6'h2b == _T_11317_46; // @[Mux.scala 46:19:@13285.4]
  assign _T_14862 = _T_14861 ? _T_10366_42 : _T_14860; // @[Mux.scala 46:16:@13286.4]
  assign _T_14863 = 6'h2a == _T_11317_46; // @[Mux.scala 46:19:@13287.4]
  assign _T_14864 = _T_14863 ? _T_10366_41 : _T_14862; // @[Mux.scala 46:16:@13288.4]
  assign _T_14865 = 6'h29 == _T_11317_46; // @[Mux.scala 46:19:@13289.4]
  assign _T_14866 = _T_14865 ? _T_10366_40 : _T_14864; // @[Mux.scala 46:16:@13290.4]
  assign _T_14867 = 6'h28 == _T_11317_46; // @[Mux.scala 46:19:@13291.4]
  assign _T_14868 = _T_14867 ? _T_10366_39 : _T_14866; // @[Mux.scala 46:16:@13292.4]
  assign _T_14869 = 6'h27 == _T_11317_46; // @[Mux.scala 46:19:@13293.4]
  assign _T_14870 = _T_14869 ? _T_10366_38 : _T_14868; // @[Mux.scala 46:16:@13294.4]
  assign _T_14871 = 6'h26 == _T_11317_46; // @[Mux.scala 46:19:@13295.4]
  assign _T_14872 = _T_14871 ? _T_10366_37 : _T_14870; // @[Mux.scala 46:16:@13296.4]
  assign _T_14873 = 6'h25 == _T_11317_46; // @[Mux.scala 46:19:@13297.4]
  assign _T_14874 = _T_14873 ? _T_10366_36 : _T_14872; // @[Mux.scala 46:16:@13298.4]
  assign _T_14875 = 6'h24 == _T_11317_46; // @[Mux.scala 46:19:@13299.4]
  assign _T_14876 = _T_14875 ? _T_10366_35 : _T_14874; // @[Mux.scala 46:16:@13300.4]
  assign _T_14877 = 6'h23 == _T_11317_46; // @[Mux.scala 46:19:@13301.4]
  assign _T_14878 = _T_14877 ? _T_10366_34 : _T_14876; // @[Mux.scala 46:16:@13302.4]
  assign _T_14879 = 6'h22 == _T_11317_46; // @[Mux.scala 46:19:@13303.4]
  assign _T_14880 = _T_14879 ? _T_10366_33 : _T_14878; // @[Mux.scala 46:16:@13304.4]
  assign _T_14881 = 6'h21 == _T_11317_46; // @[Mux.scala 46:19:@13305.4]
  assign _T_14882 = _T_14881 ? _T_10366_32 : _T_14880; // @[Mux.scala 46:16:@13306.4]
  assign _T_14883 = 6'h20 == _T_11317_46; // @[Mux.scala 46:19:@13307.4]
  assign _T_14884 = _T_14883 ? _T_10366_31 : _T_14882; // @[Mux.scala 46:16:@13308.4]
  assign _T_14885 = 6'h1f == _T_11317_46; // @[Mux.scala 46:19:@13309.4]
  assign _T_14886 = _T_14885 ? _T_10366_30 : _T_14884; // @[Mux.scala 46:16:@13310.4]
  assign _T_14887 = 6'h1e == _T_11317_46; // @[Mux.scala 46:19:@13311.4]
  assign _T_14888 = _T_14887 ? _T_10366_29 : _T_14886; // @[Mux.scala 46:16:@13312.4]
  assign _T_14889 = 6'h1d == _T_11317_46; // @[Mux.scala 46:19:@13313.4]
  assign _T_14890 = _T_14889 ? _T_10366_28 : _T_14888; // @[Mux.scala 46:16:@13314.4]
  assign _T_14891 = 6'h1c == _T_11317_46; // @[Mux.scala 46:19:@13315.4]
  assign _T_14892 = _T_14891 ? _T_10366_27 : _T_14890; // @[Mux.scala 46:16:@13316.4]
  assign _T_14893 = 6'h1b == _T_11317_46; // @[Mux.scala 46:19:@13317.4]
  assign _T_14894 = _T_14893 ? _T_10366_26 : _T_14892; // @[Mux.scala 46:16:@13318.4]
  assign _T_14895 = 6'h1a == _T_11317_46; // @[Mux.scala 46:19:@13319.4]
  assign _T_14896 = _T_14895 ? _T_10366_25 : _T_14894; // @[Mux.scala 46:16:@13320.4]
  assign _T_14897 = 6'h19 == _T_11317_46; // @[Mux.scala 46:19:@13321.4]
  assign _T_14898 = _T_14897 ? _T_10366_24 : _T_14896; // @[Mux.scala 46:16:@13322.4]
  assign _T_14899 = 6'h18 == _T_11317_46; // @[Mux.scala 46:19:@13323.4]
  assign _T_14900 = _T_14899 ? _T_10366_23 : _T_14898; // @[Mux.scala 46:16:@13324.4]
  assign _T_14901 = 6'h17 == _T_11317_46; // @[Mux.scala 46:19:@13325.4]
  assign _T_14902 = _T_14901 ? _T_10366_22 : _T_14900; // @[Mux.scala 46:16:@13326.4]
  assign _T_14903 = 6'h16 == _T_11317_46; // @[Mux.scala 46:19:@13327.4]
  assign _T_14904 = _T_14903 ? _T_10366_21 : _T_14902; // @[Mux.scala 46:16:@13328.4]
  assign _T_14905 = 6'h15 == _T_11317_46; // @[Mux.scala 46:19:@13329.4]
  assign _T_14906 = _T_14905 ? _T_10366_20 : _T_14904; // @[Mux.scala 46:16:@13330.4]
  assign _T_14907 = 6'h14 == _T_11317_46; // @[Mux.scala 46:19:@13331.4]
  assign _T_14908 = _T_14907 ? _T_10366_19 : _T_14906; // @[Mux.scala 46:16:@13332.4]
  assign _T_14909 = 6'h13 == _T_11317_46; // @[Mux.scala 46:19:@13333.4]
  assign _T_14910 = _T_14909 ? _T_10366_18 : _T_14908; // @[Mux.scala 46:16:@13334.4]
  assign _T_14911 = 6'h12 == _T_11317_46; // @[Mux.scala 46:19:@13335.4]
  assign _T_14912 = _T_14911 ? _T_10366_17 : _T_14910; // @[Mux.scala 46:16:@13336.4]
  assign _T_14913 = 6'h11 == _T_11317_46; // @[Mux.scala 46:19:@13337.4]
  assign _T_14914 = _T_14913 ? _T_10366_16 : _T_14912; // @[Mux.scala 46:16:@13338.4]
  assign _T_14915 = 6'h10 == _T_11317_46; // @[Mux.scala 46:19:@13339.4]
  assign _T_14916 = _T_14915 ? _T_10366_15 : _T_14914; // @[Mux.scala 46:16:@13340.4]
  assign _T_14917 = 6'hf == _T_11317_46; // @[Mux.scala 46:19:@13341.4]
  assign _T_14918 = _T_14917 ? _T_10366_14 : _T_14916; // @[Mux.scala 46:16:@13342.4]
  assign _T_14919 = 6'he == _T_11317_46; // @[Mux.scala 46:19:@13343.4]
  assign _T_14920 = _T_14919 ? _T_10366_13 : _T_14918; // @[Mux.scala 46:16:@13344.4]
  assign _T_14921 = 6'hd == _T_11317_46; // @[Mux.scala 46:19:@13345.4]
  assign _T_14922 = _T_14921 ? _T_10366_12 : _T_14920; // @[Mux.scala 46:16:@13346.4]
  assign _T_14923 = 6'hc == _T_11317_46; // @[Mux.scala 46:19:@13347.4]
  assign _T_14924 = _T_14923 ? _T_10366_11 : _T_14922; // @[Mux.scala 46:16:@13348.4]
  assign _T_14925 = 6'hb == _T_11317_46; // @[Mux.scala 46:19:@13349.4]
  assign _T_14926 = _T_14925 ? _T_10366_10 : _T_14924; // @[Mux.scala 46:16:@13350.4]
  assign _T_14927 = 6'ha == _T_11317_46; // @[Mux.scala 46:19:@13351.4]
  assign _T_14928 = _T_14927 ? _T_10366_9 : _T_14926; // @[Mux.scala 46:16:@13352.4]
  assign _T_14929 = 6'h9 == _T_11317_46; // @[Mux.scala 46:19:@13353.4]
  assign _T_14930 = _T_14929 ? _T_10366_8 : _T_14928; // @[Mux.scala 46:16:@13354.4]
  assign _T_14931 = 6'h8 == _T_11317_46; // @[Mux.scala 46:19:@13355.4]
  assign _T_14932 = _T_14931 ? _T_10366_7 : _T_14930; // @[Mux.scala 46:16:@13356.4]
  assign _T_14933 = 6'h7 == _T_11317_46; // @[Mux.scala 46:19:@13357.4]
  assign _T_14934 = _T_14933 ? _T_10366_6 : _T_14932; // @[Mux.scala 46:16:@13358.4]
  assign _T_14935 = 6'h6 == _T_11317_46; // @[Mux.scala 46:19:@13359.4]
  assign _T_14936 = _T_14935 ? _T_10366_5 : _T_14934; // @[Mux.scala 46:16:@13360.4]
  assign _T_14937 = 6'h5 == _T_11317_46; // @[Mux.scala 46:19:@13361.4]
  assign _T_14938 = _T_14937 ? _T_10366_4 : _T_14936; // @[Mux.scala 46:16:@13362.4]
  assign _T_14939 = 6'h4 == _T_11317_46; // @[Mux.scala 46:19:@13363.4]
  assign _T_14940 = _T_14939 ? _T_10366_3 : _T_14938; // @[Mux.scala 46:16:@13364.4]
  assign _T_14941 = 6'h3 == _T_11317_46; // @[Mux.scala 46:19:@13365.4]
  assign _T_14942 = _T_14941 ? _T_10366_2 : _T_14940; // @[Mux.scala 46:16:@13366.4]
  assign _T_14943 = 6'h2 == _T_11317_46; // @[Mux.scala 46:19:@13367.4]
  assign _T_14944 = _T_14943 ? _T_10366_1 : _T_14942; // @[Mux.scala 46:16:@13368.4]
  assign _T_14945 = 6'h1 == _T_11317_46; // @[Mux.scala 46:19:@13369.4]
  assign _T_14946 = _T_14945 ? _T_10366_0 : _T_14944; // @[Mux.scala 46:16:@13370.4]
  assign _T_14996 = 6'h30 == _T_11317_47; // @[Mux.scala 46:19:@13372.4]
  assign _T_14997 = _T_14996 ? _T_10366_47 : 8'h0; // @[Mux.scala 46:16:@13373.4]
  assign _T_14998 = 6'h2f == _T_11317_47; // @[Mux.scala 46:19:@13374.4]
  assign _T_14999 = _T_14998 ? _T_10366_46 : _T_14997; // @[Mux.scala 46:16:@13375.4]
  assign _T_15000 = 6'h2e == _T_11317_47; // @[Mux.scala 46:19:@13376.4]
  assign _T_15001 = _T_15000 ? _T_10366_45 : _T_14999; // @[Mux.scala 46:16:@13377.4]
  assign _T_15002 = 6'h2d == _T_11317_47; // @[Mux.scala 46:19:@13378.4]
  assign _T_15003 = _T_15002 ? _T_10366_44 : _T_15001; // @[Mux.scala 46:16:@13379.4]
  assign _T_15004 = 6'h2c == _T_11317_47; // @[Mux.scala 46:19:@13380.4]
  assign _T_15005 = _T_15004 ? _T_10366_43 : _T_15003; // @[Mux.scala 46:16:@13381.4]
  assign _T_15006 = 6'h2b == _T_11317_47; // @[Mux.scala 46:19:@13382.4]
  assign _T_15007 = _T_15006 ? _T_10366_42 : _T_15005; // @[Mux.scala 46:16:@13383.4]
  assign _T_15008 = 6'h2a == _T_11317_47; // @[Mux.scala 46:19:@13384.4]
  assign _T_15009 = _T_15008 ? _T_10366_41 : _T_15007; // @[Mux.scala 46:16:@13385.4]
  assign _T_15010 = 6'h29 == _T_11317_47; // @[Mux.scala 46:19:@13386.4]
  assign _T_15011 = _T_15010 ? _T_10366_40 : _T_15009; // @[Mux.scala 46:16:@13387.4]
  assign _T_15012 = 6'h28 == _T_11317_47; // @[Mux.scala 46:19:@13388.4]
  assign _T_15013 = _T_15012 ? _T_10366_39 : _T_15011; // @[Mux.scala 46:16:@13389.4]
  assign _T_15014 = 6'h27 == _T_11317_47; // @[Mux.scala 46:19:@13390.4]
  assign _T_15015 = _T_15014 ? _T_10366_38 : _T_15013; // @[Mux.scala 46:16:@13391.4]
  assign _T_15016 = 6'h26 == _T_11317_47; // @[Mux.scala 46:19:@13392.4]
  assign _T_15017 = _T_15016 ? _T_10366_37 : _T_15015; // @[Mux.scala 46:16:@13393.4]
  assign _T_15018 = 6'h25 == _T_11317_47; // @[Mux.scala 46:19:@13394.4]
  assign _T_15019 = _T_15018 ? _T_10366_36 : _T_15017; // @[Mux.scala 46:16:@13395.4]
  assign _T_15020 = 6'h24 == _T_11317_47; // @[Mux.scala 46:19:@13396.4]
  assign _T_15021 = _T_15020 ? _T_10366_35 : _T_15019; // @[Mux.scala 46:16:@13397.4]
  assign _T_15022 = 6'h23 == _T_11317_47; // @[Mux.scala 46:19:@13398.4]
  assign _T_15023 = _T_15022 ? _T_10366_34 : _T_15021; // @[Mux.scala 46:16:@13399.4]
  assign _T_15024 = 6'h22 == _T_11317_47; // @[Mux.scala 46:19:@13400.4]
  assign _T_15025 = _T_15024 ? _T_10366_33 : _T_15023; // @[Mux.scala 46:16:@13401.4]
  assign _T_15026 = 6'h21 == _T_11317_47; // @[Mux.scala 46:19:@13402.4]
  assign _T_15027 = _T_15026 ? _T_10366_32 : _T_15025; // @[Mux.scala 46:16:@13403.4]
  assign _T_15028 = 6'h20 == _T_11317_47; // @[Mux.scala 46:19:@13404.4]
  assign _T_15029 = _T_15028 ? _T_10366_31 : _T_15027; // @[Mux.scala 46:16:@13405.4]
  assign _T_15030 = 6'h1f == _T_11317_47; // @[Mux.scala 46:19:@13406.4]
  assign _T_15031 = _T_15030 ? _T_10366_30 : _T_15029; // @[Mux.scala 46:16:@13407.4]
  assign _T_15032 = 6'h1e == _T_11317_47; // @[Mux.scala 46:19:@13408.4]
  assign _T_15033 = _T_15032 ? _T_10366_29 : _T_15031; // @[Mux.scala 46:16:@13409.4]
  assign _T_15034 = 6'h1d == _T_11317_47; // @[Mux.scala 46:19:@13410.4]
  assign _T_15035 = _T_15034 ? _T_10366_28 : _T_15033; // @[Mux.scala 46:16:@13411.4]
  assign _T_15036 = 6'h1c == _T_11317_47; // @[Mux.scala 46:19:@13412.4]
  assign _T_15037 = _T_15036 ? _T_10366_27 : _T_15035; // @[Mux.scala 46:16:@13413.4]
  assign _T_15038 = 6'h1b == _T_11317_47; // @[Mux.scala 46:19:@13414.4]
  assign _T_15039 = _T_15038 ? _T_10366_26 : _T_15037; // @[Mux.scala 46:16:@13415.4]
  assign _T_15040 = 6'h1a == _T_11317_47; // @[Mux.scala 46:19:@13416.4]
  assign _T_15041 = _T_15040 ? _T_10366_25 : _T_15039; // @[Mux.scala 46:16:@13417.4]
  assign _T_15042 = 6'h19 == _T_11317_47; // @[Mux.scala 46:19:@13418.4]
  assign _T_15043 = _T_15042 ? _T_10366_24 : _T_15041; // @[Mux.scala 46:16:@13419.4]
  assign _T_15044 = 6'h18 == _T_11317_47; // @[Mux.scala 46:19:@13420.4]
  assign _T_15045 = _T_15044 ? _T_10366_23 : _T_15043; // @[Mux.scala 46:16:@13421.4]
  assign _T_15046 = 6'h17 == _T_11317_47; // @[Mux.scala 46:19:@13422.4]
  assign _T_15047 = _T_15046 ? _T_10366_22 : _T_15045; // @[Mux.scala 46:16:@13423.4]
  assign _T_15048 = 6'h16 == _T_11317_47; // @[Mux.scala 46:19:@13424.4]
  assign _T_15049 = _T_15048 ? _T_10366_21 : _T_15047; // @[Mux.scala 46:16:@13425.4]
  assign _T_15050 = 6'h15 == _T_11317_47; // @[Mux.scala 46:19:@13426.4]
  assign _T_15051 = _T_15050 ? _T_10366_20 : _T_15049; // @[Mux.scala 46:16:@13427.4]
  assign _T_15052 = 6'h14 == _T_11317_47; // @[Mux.scala 46:19:@13428.4]
  assign _T_15053 = _T_15052 ? _T_10366_19 : _T_15051; // @[Mux.scala 46:16:@13429.4]
  assign _T_15054 = 6'h13 == _T_11317_47; // @[Mux.scala 46:19:@13430.4]
  assign _T_15055 = _T_15054 ? _T_10366_18 : _T_15053; // @[Mux.scala 46:16:@13431.4]
  assign _T_15056 = 6'h12 == _T_11317_47; // @[Mux.scala 46:19:@13432.4]
  assign _T_15057 = _T_15056 ? _T_10366_17 : _T_15055; // @[Mux.scala 46:16:@13433.4]
  assign _T_15058 = 6'h11 == _T_11317_47; // @[Mux.scala 46:19:@13434.4]
  assign _T_15059 = _T_15058 ? _T_10366_16 : _T_15057; // @[Mux.scala 46:16:@13435.4]
  assign _T_15060 = 6'h10 == _T_11317_47; // @[Mux.scala 46:19:@13436.4]
  assign _T_15061 = _T_15060 ? _T_10366_15 : _T_15059; // @[Mux.scala 46:16:@13437.4]
  assign _T_15062 = 6'hf == _T_11317_47; // @[Mux.scala 46:19:@13438.4]
  assign _T_15063 = _T_15062 ? _T_10366_14 : _T_15061; // @[Mux.scala 46:16:@13439.4]
  assign _T_15064 = 6'he == _T_11317_47; // @[Mux.scala 46:19:@13440.4]
  assign _T_15065 = _T_15064 ? _T_10366_13 : _T_15063; // @[Mux.scala 46:16:@13441.4]
  assign _T_15066 = 6'hd == _T_11317_47; // @[Mux.scala 46:19:@13442.4]
  assign _T_15067 = _T_15066 ? _T_10366_12 : _T_15065; // @[Mux.scala 46:16:@13443.4]
  assign _T_15068 = 6'hc == _T_11317_47; // @[Mux.scala 46:19:@13444.4]
  assign _T_15069 = _T_15068 ? _T_10366_11 : _T_15067; // @[Mux.scala 46:16:@13445.4]
  assign _T_15070 = 6'hb == _T_11317_47; // @[Mux.scala 46:19:@13446.4]
  assign _T_15071 = _T_15070 ? _T_10366_10 : _T_15069; // @[Mux.scala 46:16:@13447.4]
  assign _T_15072 = 6'ha == _T_11317_47; // @[Mux.scala 46:19:@13448.4]
  assign _T_15073 = _T_15072 ? _T_10366_9 : _T_15071; // @[Mux.scala 46:16:@13449.4]
  assign _T_15074 = 6'h9 == _T_11317_47; // @[Mux.scala 46:19:@13450.4]
  assign _T_15075 = _T_15074 ? _T_10366_8 : _T_15073; // @[Mux.scala 46:16:@13451.4]
  assign _T_15076 = 6'h8 == _T_11317_47; // @[Mux.scala 46:19:@13452.4]
  assign _T_15077 = _T_15076 ? _T_10366_7 : _T_15075; // @[Mux.scala 46:16:@13453.4]
  assign _T_15078 = 6'h7 == _T_11317_47; // @[Mux.scala 46:19:@13454.4]
  assign _T_15079 = _T_15078 ? _T_10366_6 : _T_15077; // @[Mux.scala 46:16:@13455.4]
  assign _T_15080 = 6'h6 == _T_11317_47; // @[Mux.scala 46:19:@13456.4]
  assign _T_15081 = _T_15080 ? _T_10366_5 : _T_15079; // @[Mux.scala 46:16:@13457.4]
  assign _T_15082 = 6'h5 == _T_11317_47; // @[Mux.scala 46:19:@13458.4]
  assign _T_15083 = _T_15082 ? _T_10366_4 : _T_15081; // @[Mux.scala 46:16:@13459.4]
  assign _T_15084 = 6'h4 == _T_11317_47; // @[Mux.scala 46:19:@13460.4]
  assign _T_15085 = _T_15084 ? _T_10366_3 : _T_15083; // @[Mux.scala 46:16:@13461.4]
  assign _T_15086 = 6'h3 == _T_11317_47; // @[Mux.scala 46:19:@13462.4]
  assign _T_15087 = _T_15086 ? _T_10366_2 : _T_15085; // @[Mux.scala 46:16:@13463.4]
  assign _T_15088 = 6'h2 == _T_11317_47; // @[Mux.scala 46:19:@13464.4]
  assign _T_15089 = _T_15088 ? _T_10366_1 : _T_15087; // @[Mux.scala 46:16:@13465.4]
  assign _T_15090 = 6'h1 == _T_11317_47; // @[Mux.scala 46:19:@13466.4]
  assign _T_15091 = _T_15090 ? _T_10366_0 : _T_15089; // @[Mux.scala 46:16:@13467.4]
  assign _T_15142 = 6'h31 == _T_11317_48; // @[Mux.scala 46:19:@13469.4]
  assign _T_15143 = _T_15142 ? _T_10366_48 : 8'h0; // @[Mux.scala 46:16:@13470.4]
  assign _T_15144 = 6'h30 == _T_11317_48; // @[Mux.scala 46:19:@13471.4]
  assign _T_15145 = _T_15144 ? _T_10366_47 : _T_15143; // @[Mux.scala 46:16:@13472.4]
  assign _T_15146 = 6'h2f == _T_11317_48; // @[Mux.scala 46:19:@13473.4]
  assign _T_15147 = _T_15146 ? _T_10366_46 : _T_15145; // @[Mux.scala 46:16:@13474.4]
  assign _T_15148 = 6'h2e == _T_11317_48; // @[Mux.scala 46:19:@13475.4]
  assign _T_15149 = _T_15148 ? _T_10366_45 : _T_15147; // @[Mux.scala 46:16:@13476.4]
  assign _T_15150 = 6'h2d == _T_11317_48; // @[Mux.scala 46:19:@13477.4]
  assign _T_15151 = _T_15150 ? _T_10366_44 : _T_15149; // @[Mux.scala 46:16:@13478.4]
  assign _T_15152 = 6'h2c == _T_11317_48; // @[Mux.scala 46:19:@13479.4]
  assign _T_15153 = _T_15152 ? _T_10366_43 : _T_15151; // @[Mux.scala 46:16:@13480.4]
  assign _T_15154 = 6'h2b == _T_11317_48; // @[Mux.scala 46:19:@13481.4]
  assign _T_15155 = _T_15154 ? _T_10366_42 : _T_15153; // @[Mux.scala 46:16:@13482.4]
  assign _T_15156 = 6'h2a == _T_11317_48; // @[Mux.scala 46:19:@13483.4]
  assign _T_15157 = _T_15156 ? _T_10366_41 : _T_15155; // @[Mux.scala 46:16:@13484.4]
  assign _T_15158 = 6'h29 == _T_11317_48; // @[Mux.scala 46:19:@13485.4]
  assign _T_15159 = _T_15158 ? _T_10366_40 : _T_15157; // @[Mux.scala 46:16:@13486.4]
  assign _T_15160 = 6'h28 == _T_11317_48; // @[Mux.scala 46:19:@13487.4]
  assign _T_15161 = _T_15160 ? _T_10366_39 : _T_15159; // @[Mux.scala 46:16:@13488.4]
  assign _T_15162 = 6'h27 == _T_11317_48; // @[Mux.scala 46:19:@13489.4]
  assign _T_15163 = _T_15162 ? _T_10366_38 : _T_15161; // @[Mux.scala 46:16:@13490.4]
  assign _T_15164 = 6'h26 == _T_11317_48; // @[Mux.scala 46:19:@13491.4]
  assign _T_15165 = _T_15164 ? _T_10366_37 : _T_15163; // @[Mux.scala 46:16:@13492.4]
  assign _T_15166 = 6'h25 == _T_11317_48; // @[Mux.scala 46:19:@13493.4]
  assign _T_15167 = _T_15166 ? _T_10366_36 : _T_15165; // @[Mux.scala 46:16:@13494.4]
  assign _T_15168 = 6'h24 == _T_11317_48; // @[Mux.scala 46:19:@13495.4]
  assign _T_15169 = _T_15168 ? _T_10366_35 : _T_15167; // @[Mux.scala 46:16:@13496.4]
  assign _T_15170 = 6'h23 == _T_11317_48; // @[Mux.scala 46:19:@13497.4]
  assign _T_15171 = _T_15170 ? _T_10366_34 : _T_15169; // @[Mux.scala 46:16:@13498.4]
  assign _T_15172 = 6'h22 == _T_11317_48; // @[Mux.scala 46:19:@13499.4]
  assign _T_15173 = _T_15172 ? _T_10366_33 : _T_15171; // @[Mux.scala 46:16:@13500.4]
  assign _T_15174 = 6'h21 == _T_11317_48; // @[Mux.scala 46:19:@13501.4]
  assign _T_15175 = _T_15174 ? _T_10366_32 : _T_15173; // @[Mux.scala 46:16:@13502.4]
  assign _T_15176 = 6'h20 == _T_11317_48; // @[Mux.scala 46:19:@13503.4]
  assign _T_15177 = _T_15176 ? _T_10366_31 : _T_15175; // @[Mux.scala 46:16:@13504.4]
  assign _T_15178 = 6'h1f == _T_11317_48; // @[Mux.scala 46:19:@13505.4]
  assign _T_15179 = _T_15178 ? _T_10366_30 : _T_15177; // @[Mux.scala 46:16:@13506.4]
  assign _T_15180 = 6'h1e == _T_11317_48; // @[Mux.scala 46:19:@13507.4]
  assign _T_15181 = _T_15180 ? _T_10366_29 : _T_15179; // @[Mux.scala 46:16:@13508.4]
  assign _T_15182 = 6'h1d == _T_11317_48; // @[Mux.scala 46:19:@13509.4]
  assign _T_15183 = _T_15182 ? _T_10366_28 : _T_15181; // @[Mux.scala 46:16:@13510.4]
  assign _T_15184 = 6'h1c == _T_11317_48; // @[Mux.scala 46:19:@13511.4]
  assign _T_15185 = _T_15184 ? _T_10366_27 : _T_15183; // @[Mux.scala 46:16:@13512.4]
  assign _T_15186 = 6'h1b == _T_11317_48; // @[Mux.scala 46:19:@13513.4]
  assign _T_15187 = _T_15186 ? _T_10366_26 : _T_15185; // @[Mux.scala 46:16:@13514.4]
  assign _T_15188 = 6'h1a == _T_11317_48; // @[Mux.scala 46:19:@13515.4]
  assign _T_15189 = _T_15188 ? _T_10366_25 : _T_15187; // @[Mux.scala 46:16:@13516.4]
  assign _T_15190 = 6'h19 == _T_11317_48; // @[Mux.scala 46:19:@13517.4]
  assign _T_15191 = _T_15190 ? _T_10366_24 : _T_15189; // @[Mux.scala 46:16:@13518.4]
  assign _T_15192 = 6'h18 == _T_11317_48; // @[Mux.scala 46:19:@13519.4]
  assign _T_15193 = _T_15192 ? _T_10366_23 : _T_15191; // @[Mux.scala 46:16:@13520.4]
  assign _T_15194 = 6'h17 == _T_11317_48; // @[Mux.scala 46:19:@13521.4]
  assign _T_15195 = _T_15194 ? _T_10366_22 : _T_15193; // @[Mux.scala 46:16:@13522.4]
  assign _T_15196 = 6'h16 == _T_11317_48; // @[Mux.scala 46:19:@13523.4]
  assign _T_15197 = _T_15196 ? _T_10366_21 : _T_15195; // @[Mux.scala 46:16:@13524.4]
  assign _T_15198 = 6'h15 == _T_11317_48; // @[Mux.scala 46:19:@13525.4]
  assign _T_15199 = _T_15198 ? _T_10366_20 : _T_15197; // @[Mux.scala 46:16:@13526.4]
  assign _T_15200 = 6'h14 == _T_11317_48; // @[Mux.scala 46:19:@13527.4]
  assign _T_15201 = _T_15200 ? _T_10366_19 : _T_15199; // @[Mux.scala 46:16:@13528.4]
  assign _T_15202 = 6'h13 == _T_11317_48; // @[Mux.scala 46:19:@13529.4]
  assign _T_15203 = _T_15202 ? _T_10366_18 : _T_15201; // @[Mux.scala 46:16:@13530.4]
  assign _T_15204 = 6'h12 == _T_11317_48; // @[Mux.scala 46:19:@13531.4]
  assign _T_15205 = _T_15204 ? _T_10366_17 : _T_15203; // @[Mux.scala 46:16:@13532.4]
  assign _T_15206 = 6'h11 == _T_11317_48; // @[Mux.scala 46:19:@13533.4]
  assign _T_15207 = _T_15206 ? _T_10366_16 : _T_15205; // @[Mux.scala 46:16:@13534.4]
  assign _T_15208 = 6'h10 == _T_11317_48; // @[Mux.scala 46:19:@13535.4]
  assign _T_15209 = _T_15208 ? _T_10366_15 : _T_15207; // @[Mux.scala 46:16:@13536.4]
  assign _T_15210 = 6'hf == _T_11317_48; // @[Mux.scala 46:19:@13537.4]
  assign _T_15211 = _T_15210 ? _T_10366_14 : _T_15209; // @[Mux.scala 46:16:@13538.4]
  assign _T_15212 = 6'he == _T_11317_48; // @[Mux.scala 46:19:@13539.4]
  assign _T_15213 = _T_15212 ? _T_10366_13 : _T_15211; // @[Mux.scala 46:16:@13540.4]
  assign _T_15214 = 6'hd == _T_11317_48; // @[Mux.scala 46:19:@13541.4]
  assign _T_15215 = _T_15214 ? _T_10366_12 : _T_15213; // @[Mux.scala 46:16:@13542.4]
  assign _T_15216 = 6'hc == _T_11317_48; // @[Mux.scala 46:19:@13543.4]
  assign _T_15217 = _T_15216 ? _T_10366_11 : _T_15215; // @[Mux.scala 46:16:@13544.4]
  assign _T_15218 = 6'hb == _T_11317_48; // @[Mux.scala 46:19:@13545.4]
  assign _T_15219 = _T_15218 ? _T_10366_10 : _T_15217; // @[Mux.scala 46:16:@13546.4]
  assign _T_15220 = 6'ha == _T_11317_48; // @[Mux.scala 46:19:@13547.4]
  assign _T_15221 = _T_15220 ? _T_10366_9 : _T_15219; // @[Mux.scala 46:16:@13548.4]
  assign _T_15222 = 6'h9 == _T_11317_48; // @[Mux.scala 46:19:@13549.4]
  assign _T_15223 = _T_15222 ? _T_10366_8 : _T_15221; // @[Mux.scala 46:16:@13550.4]
  assign _T_15224 = 6'h8 == _T_11317_48; // @[Mux.scala 46:19:@13551.4]
  assign _T_15225 = _T_15224 ? _T_10366_7 : _T_15223; // @[Mux.scala 46:16:@13552.4]
  assign _T_15226 = 6'h7 == _T_11317_48; // @[Mux.scala 46:19:@13553.4]
  assign _T_15227 = _T_15226 ? _T_10366_6 : _T_15225; // @[Mux.scala 46:16:@13554.4]
  assign _T_15228 = 6'h6 == _T_11317_48; // @[Mux.scala 46:19:@13555.4]
  assign _T_15229 = _T_15228 ? _T_10366_5 : _T_15227; // @[Mux.scala 46:16:@13556.4]
  assign _T_15230 = 6'h5 == _T_11317_48; // @[Mux.scala 46:19:@13557.4]
  assign _T_15231 = _T_15230 ? _T_10366_4 : _T_15229; // @[Mux.scala 46:16:@13558.4]
  assign _T_15232 = 6'h4 == _T_11317_48; // @[Mux.scala 46:19:@13559.4]
  assign _T_15233 = _T_15232 ? _T_10366_3 : _T_15231; // @[Mux.scala 46:16:@13560.4]
  assign _T_15234 = 6'h3 == _T_11317_48; // @[Mux.scala 46:19:@13561.4]
  assign _T_15235 = _T_15234 ? _T_10366_2 : _T_15233; // @[Mux.scala 46:16:@13562.4]
  assign _T_15236 = 6'h2 == _T_11317_48; // @[Mux.scala 46:19:@13563.4]
  assign _T_15237 = _T_15236 ? _T_10366_1 : _T_15235; // @[Mux.scala 46:16:@13564.4]
  assign _T_15238 = 6'h1 == _T_11317_48; // @[Mux.scala 46:19:@13565.4]
  assign _T_15239 = _T_15238 ? _T_10366_0 : _T_15237; // @[Mux.scala 46:16:@13566.4]
  assign _T_15291 = 6'h32 == _T_11317_49; // @[Mux.scala 46:19:@13568.4]
  assign _T_15292 = _T_15291 ? _T_10366_49 : 8'h0; // @[Mux.scala 46:16:@13569.4]
  assign _T_15293 = 6'h31 == _T_11317_49; // @[Mux.scala 46:19:@13570.4]
  assign _T_15294 = _T_15293 ? _T_10366_48 : _T_15292; // @[Mux.scala 46:16:@13571.4]
  assign _T_15295 = 6'h30 == _T_11317_49; // @[Mux.scala 46:19:@13572.4]
  assign _T_15296 = _T_15295 ? _T_10366_47 : _T_15294; // @[Mux.scala 46:16:@13573.4]
  assign _T_15297 = 6'h2f == _T_11317_49; // @[Mux.scala 46:19:@13574.4]
  assign _T_15298 = _T_15297 ? _T_10366_46 : _T_15296; // @[Mux.scala 46:16:@13575.4]
  assign _T_15299 = 6'h2e == _T_11317_49; // @[Mux.scala 46:19:@13576.4]
  assign _T_15300 = _T_15299 ? _T_10366_45 : _T_15298; // @[Mux.scala 46:16:@13577.4]
  assign _T_15301 = 6'h2d == _T_11317_49; // @[Mux.scala 46:19:@13578.4]
  assign _T_15302 = _T_15301 ? _T_10366_44 : _T_15300; // @[Mux.scala 46:16:@13579.4]
  assign _T_15303 = 6'h2c == _T_11317_49; // @[Mux.scala 46:19:@13580.4]
  assign _T_15304 = _T_15303 ? _T_10366_43 : _T_15302; // @[Mux.scala 46:16:@13581.4]
  assign _T_15305 = 6'h2b == _T_11317_49; // @[Mux.scala 46:19:@13582.4]
  assign _T_15306 = _T_15305 ? _T_10366_42 : _T_15304; // @[Mux.scala 46:16:@13583.4]
  assign _T_15307 = 6'h2a == _T_11317_49; // @[Mux.scala 46:19:@13584.4]
  assign _T_15308 = _T_15307 ? _T_10366_41 : _T_15306; // @[Mux.scala 46:16:@13585.4]
  assign _T_15309 = 6'h29 == _T_11317_49; // @[Mux.scala 46:19:@13586.4]
  assign _T_15310 = _T_15309 ? _T_10366_40 : _T_15308; // @[Mux.scala 46:16:@13587.4]
  assign _T_15311 = 6'h28 == _T_11317_49; // @[Mux.scala 46:19:@13588.4]
  assign _T_15312 = _T_15311 ? _T_10366_39 : _T_15310; // @[Mux.scala 46:16:@13589.4]
  assign _T_15313 = 6'h27 == _T_11317_49; // @[Mux.scala 46:19:@13590.4]
  assign _T_15314 = _T_15313 ? _T_10366_38 : _T_15312; // @[Mux.scala 46:16:@13591.4]
  assign _T_15315 = 6'h26 == _T_11317_49; // @[Mux.scala 46:19:@13592.4]
  assign _T_15316 = _T_15315 ? _T_10366_37 : _T_15314; // @[Mux.scala 46:16:@13593.4]
  assign _T_15317 = 6'h25 == _T_11317_49; // @[Mux.scala 46:19:@13594.4]
  assign _T_15318 = _T_15317 ? _T_10366_36 : _T_15316; // @[Mux.scala 46:16:@13595.4]
  assign _T_15319 = 6'h24 == _T_11317_49; // @[Mux.scala 46:19:@13596.4]
  assign _T_15320 = _T_15319 ? _T_10366_35 : _T_15318; // @[Mux.scala 46:16:@13597.4]
  assign _T_15321 = 6'h23 == _T_11317_49; // @[Mux.scala 46:19:@13598.4]
  assign _T_15322 = _T_15321 ? _T_10366_34 : _T_15320; // @[Mux.scala 46:16:@13599.4]
  assign _T_15323 = 6'h22 == _T_11317_49; // @[Mux.scala 46:19:@13600.4]
  assign _T_15324 = _T_15323 ? _T_10366_33 : _T_15322; // @[Mux.scala 46:16:@13601.4]
  assign _T_15325 = 6'h21 == _T_11317_49; // @[Mux.scala 46:19:@13602.4]
  assign _T_15326 = _T_15325 ? _T_10366_32 : _T_15324; // @[Mux.scala 46:16:@13603.4]
  assign _T_15327 = 6'h20 == _T_11317_49; // @[Mux.scala 46:19:@13604.4]
  assign _T_15328 = _T_15327 ? _T_10366_31 : _T_15326; // @[Mux.scala 46:16:@13605.4]
  assign _T_15329 = 6'h1f == _T_11317_49; // @[Mux.scala 46:19:@13606.4]
  assign _T_15330 = _T_15329 ? _T_10366_30 : _T_15328; // @[Mux.scala 46:16:@13607.4]
  assign _T_15331 = 6'h1e == _T_11317_49; // @[Mux.scala 46:19:@13608.4]
  assign _T_15332 = _T_15331 ? _T_10366_29 : _T_15330; // @[Mux.scala 46:16:@13609.4]
  assign _T_15333 = 6'h1d == _T_11317_49; // @[Mux.scala 46:19:@13610.4]
  assign _T_15334 = _T_15333 ? _T_10366_28 : _T_15332; // @[Mux.scala 46:16:@13611.4]
  assign _T_15335 = 6'h1c == _T_11317_49; // @[Mux.scala 46:19:@13612.4]
  assign _T_15336 = _T_15335 ? _T_10366_27 : _T_15334; // @[Mux.scala 46:16:@13613.4]
  assign _T_15337 = 6'h1b == _T_11317_49; // @[Mux.scala 46:19:@13614.4]
  assign _T_15338 = _T_15337 ? _T_10366_26 : _T_15336; // @[Mux.scala 46:16:@13615.4]
  assign _T_15339 = 6'h1a == _T_11317_49; // @[Mux.scala 46:19:@13616.4]
  assign _T_15340 = _T_15339 ? _T_10366_25 : _T_15338; // @[Mux.scala 46:16:@13617.4]
  assign _T_15341 = 6'h19 == _T_11317_49; // @[Mux.scala 46:19:@13618.4]
  assign _T_15342 = _T_15341 ? _T_10366_24 : _T_15340; // @[Mux.scala 46:16:@13619.4]
  assign _T_15343 = 6'h18 == _T_11317_49; // @[Mux.scala 46:19:@13620.4]
  assign _T_15344 = _T_15343 ? _T_10366_23 : _T_15342; // @[Mux.scala 46:16:@13621.4]
  assign _T_15345 = 6'h17 == _T_11317_49; // @[Mux.scala 46:19:@13622.4]
  assign _T_15346 = _T_15345 ? _T_10366_22 : _T_15344; // @[Mux.scala 46:16:@13623.4]
  assign _T_15347 = 6'h16 == _T_11317_49; // @[Mux.scala 46:19:@13624.4]
  assign _T_15348 = _T_15347 ? _T_10366_21 : _T_15346; // @[Mux.scala 46:16:@13625.4]
  assign _T_15349 = 6'h15 == _T_11317_49; // @[Mux.scala 46:19:@13626.4]
  assign _T_15350 = _T_15349 ? _T_10366_20 : _T_15348; // @[Mux.scala 46:16:@13627.4]
  assign _T_15351 = 6'h14 == _T_11317_49; // @[Mux.scala 46:19:@13628.4]
  assign _T_15352 = _T_15351 ? _T_10366_19 : _T_15350; // @[Mux.scala 46:16:@13629.4]
  assign _T_15353 = 6'h13 == _T_11317_49; // @[Mux.scala 46:19:@13630.4]
  assign _T_15354 = _T_15353 ? _T_10366_18 : _T_15352; // @[Mux.scala 46:16:@13631.4]
  assign _T_15355 = 6'h12 == _T_11317_49; // @[Mux.scala 46:19:@13632.4]
  assign _T_15356 = _T_15355 ? _T_10366_17 : _T_15354; // @[Mux.scala 46:16:@13633.4]
  assign _T_15357 = 6'h11 == _T_11317_49; // @[Mux.scala 46:19:@13634.4]
  assign _T_15358 = _T_15357 ? _T_10366_16 : _T_15356; // @[Mux.scala 46:16:@13635.4]
  assign _T_15359 = 6'h10 == _T_11317_49; // @[Mux.scala 46:19:@13636.4]
  assign _T_15360 = _T_15359 ? _T_10366_15 : _T_15358; // @[Mux.scala 46:16:@13637.4]
  assign _T_15361 = 6'hf == _T_11317_49; // @[Mux.scala 46:19:@13638.4]
  assign _T_15362 = _T_15361 ? _T_10366_14 : _T_15360; // @[Mux.scala 46:16:@13639.4]
  assign _T_15363 = 6'he == _T_11317_49; // @[Mux.scala 46:19:@13640.4]
  assign _T_15364 = _T_15363 ? _T_10366_13 : _T_15362; // @[Mux.scala 46:16:@13641.4]
  assign _T_15365 = 6'hd == _T_11317_49; // @[Mux.scala 46:19:@13642.4]
  assign _T_15366 = _T_15365 ? _T_10366_12 : _T_15364; // @[Mux.scala 46:16:@13643.4]
  assign _T_15367 = 6'hc == _T_11317_49; // @[Mux.scala 46:19:@13644.4]
  assign _T_15368 = _T_15367 ? _T_10366_11 : _T_15366; // @[Mux.scala 46:16:@13645.4]
  assign _T_15369 = 6'hb == _T_11317_49; // @[Mux.scala 46:19:@13646.4]
  assign _T_15370 = _T_15369 ? _T_10366_10 : _T_15368; // @[Mux.scala 46:16:@13647.4]
  assign _T_15371 = 6'ha == _T_11317_49; // @[Mux.scala 46:19:@13648.4]
  assign _T_15372 = _T_15371 ? _T_10366_9 : _T_15370; // @[Mux.scala 46:16:@13649.4]
  assign _T_15373 = 6'h9 == _T_11317_49; // @[Mux.scala 46:19:@13650.4]
  assign _T_15374 = _T_15373 ? _T_10366_8 : _T_15372; // @[Mux.scala 46:16:@13651.4]
  assign _T_15375 = 6'h8 == _T_11317_49; // @[Mux.scala 46:19:@13652.4]
  assign _T_15376 = _T_15375 ? _T_10366_7 : _T_15374; // @[Mux.scala 46:16:@13653.4]
  assign _T_15377 = 6'h7 == _T_11317_49; // @[Mux.scala 46:19:@13654.4]
  assign _T_15378 = _T_15377 ? _T_10366_6 : _T_15376; // @[Mux.scala 46:16:@13655.4]
  assign _T_15379 = 6'h6 == _T_11317_49; // @[Mux.scala 46:19:@13656.4]
  assign _T_15380 = _T_15379 ? _T_10366_5 : _T_15378; // @[Mux.scala 46:16:@13657.4]
  assign _T_15381 = 6'h5 == _T_11317_49; // @[Mux.scala 46:19:@13658.4]
  assign _T_15382 = _T_15381 ? _T_10366_4 : _T_15380; // @[Mux.scala 46:16:@13659.4]
  assign _T_15383 = 6'h4 == _T_11317_49; // @[Mux.scala 46:19:@13660.4]
  assign _T_15384 = _T_15383 ? _T_10366_3 : _T_15382; // @[Mux.scala 46:16:@13661.4]
  assign _T_15385 = 6'h3 == _T_11317_49; // @[Mux.scala 46:19:@13662.4]
  assign _T_15386 = _T_15385 ? _T_10366_2 : _T_15384; // @[Mux.scala 46:16:@13663.4]
  assign _T_15387 = 6'h2 == _T_11317_49; // @[Mux.scala 46:19:@13664.4]
  assign _T_15388 = _T_15387 ? _T_10366_1 : _T_15386; // @[Mux.scala 46:16:@13665.4]
  assign _T_15389 = 6'h1 == _T_11317_49; // @[Mux.scala 46:19:@13666.4]
  assign _T_15390 = _T_15389 ? _T_10366_0 : _T_15388; // @[Mux.scala 46:16:@13667.4]
  assign _T_15443 = 6'h33 == _T_11317_50; // @[Mux.scala 46:19:@13669.4]
  assign _T_15444 = _T_15443 ? _T_10366_50 : 8'h0; // @[Mux.scala 46:16:@13670.4]
  assign _T_15445 = 6'h32 == _T_11317_50; // @[Mux.scala 46:19:@13671.4]
  assign _T_15446 = _T_15445 ? _T_10366_49 : _T_15444; // @[Mux.scala 46:16:@13672.4]
  assign _T_15447 = 6'h31 == _T_11317_50; // @[Mux.scala 46:19:@13673.4]
  assign _T_15448 = _T_15447 ? _T_10366_48 : _T_15446; // @[Mux.scala 46:16:@13674.4]
  assign _T_15449 = 6'h30 == _T_11317_50; // @[Mux.scala 46:19:@13675.4]
  assign _T_15450 = _T_15449 ? _T_10366_47 : _T_15448; // @[Mux.scala 46:16:@13676.4]
  assign _T_15451 = 6'h2f == _T_11317_50; // @[Mux.scala 46:19:@13677.4]
  assign _T_15452 = _T_15451 ? _T_10366_46 : _T_15450; // @[Mux.scala 46:16:@13678.4]
  assign _T_15453 = 6'h2e == _T_11317_50; // @[Mux.scala 46:19:@13679.4]
  assign _T_15454 = _T_15453 ? _T_10366_45 : _T_15452; // @[Mux.scala 46:16:@13680.4]
  assign _T_15455 = 6'h2d == _T_11317_50; // @[Mux.scala 46:19:@13681.4]
  assign _T_15456 = _T_15455 ? _T_10366_44 : _T_15454; // @[Mux.scala 46:16:@13682.4]
  assign _T_15457 = 6'h2c == _T_11317_50; // @[Mux.scala 46:19:@13683.4]
  assign _T_15458 = _T_15457 ? _T_10366_43 : _T_15456; // @[Mux.scala 46:16:@13684.4]
  assign _T_15459 = 6'h2b == _T_11317_50; // @[Mux.scala 46:19:@13685.4]
  assign _T_15460 = _T_15459 ? _T_10366_42 : _T_15458; // @[Mux.scala 46:16:@13686.4]
  assign _T_15461 = 6'h2a == _T_11317_50; // @[Mux.scala 46:19:@13687.4]
  assign _T_15462 = _T_15461 ? _T_10366_41 : _T_15460; // @[Mux.scala 46:16:@13688.4]
  assign _T_15463 = 6'h29 == _T_11317_50; // @[Mux.scala 46:19:@13689.4]
  assign _T_15464 = _T_15463 ? _T_10366_40 : _T_15462; // @[Mux.scala 46:16:@13690.4]
  assign _T_15465 = 6'h28 == _T_11317_50; // @[Mux.scala 46:19:@13691.4]
  assign _T_15466 = _T_15465 ? _T_10366_39 : _T_15464; // @[Mux.scala 46:16:@13692.4]
  assign _T_15467 = 6'h27 == _T_11317_50; // @[Mux.scala 46:19:@13693.4]
  assign _T_15468 = _T_15467 ? _T_10366_38 : _T_15466; // @[Mux.scala 46:16:@13694.4]
  assign _T_15469 = 6'h26 == _T_11317_50; // @[Mux.scala 46:19:@13695.4]
  assign _T_15470 = _T_15469 ? _T_10366_37 : _T_15468; // @[Mux.scala 46:16:@13696.4]
  assign _T_15471 = 6'h25 == _T_11317_50; // @[Mux.scala 46:19:@13697.4]
  assign _T_15472 = _T_15471 ? _T_10366_36 : _T_15470; // @[Mux.scala 46:16:@13698.4]
  assign _T_15473 = 6'h24 == _T_11317_50; // @[Mux.scala 46:19:@13699.4]
  assign _T_15474 = _T_15473 ? _T_10366_35 : _T_15472; // @[Mux.scala 46:16:@13700.4]
  assign _T_15475 = 6'h23 == _T_11317_50; // @[Mux.scala 46:19:@13701.4]
  assign _T_15476 = _T_15475 ? _T_10366_34 : _T_15474; // @[Mux.scala 46:16:@13702.4]
  assign _T_15477 = 6'h22 == _T_11317_50; // @[Mux.scala 46:19:@13703.4]
  assign _T_15478 = _T_15477 ? _T_10366_33 : _T_15476; // @[Mux.scala 46:16:@13704.4]
  assign _T_15479 = 6'h21 == _T_11317_50; // @[Mux.scala 46:19:@13705.4]
  assign _T_15480 = _T_15479 ? _T_10366_32 : _T_15478; // @[Mux.scala 46:16:@13706.4]
  assign _T_15481 = 6'h20 == _T_11317_50; // @[Mux.scala 46:19:@13707.4]
  assign _T_15482 = _T_15481 ? _T_10366_31 : _T_15480; // @[Mux.scala 46:16:@13708.4]
  assign _T_15483 = 6'h1f == _T_11317_50; // @[Mux.scala 46:19:@13709.4]
  assign _T_15484 = _T_15483 ? _T_10366_30 : _T_15482; // @[Mux.scala 46:16:@13710.4]
  assign _T_15485 = 6'h1e == _T_11317_50; // @[Mux.scala 46:19:@13711.4]
  assign _T_15486 = _T_15485 ? _T_10366_29 : _T_15484; // @[Mux.scala 46:16:@13712.4]
  assign _T_15487 = 6'h1d == _T_11317_50; // @[Mux.scala 46:19:@13713.4]
  assign _T_15488 = _T_15487 ? _T_10366_28 : _T_15486; // @[Mux.scala 46:16:@13714.4]
  assign _T_15489 = 6'h1c == _T_11317_50; // @[Mux.scala 46:19:@13715.4]
  assign _T_15490 = _T_15489 ? _T_10366_27 : _T_15488; // @[Mux.scala 46:16:@13716.4]
  assign _T_15491 = 6'h1b == _T_11317_50; // @[Mux.scala 46:19:@13717.4]
  assign _T_15492 = _T_15491 ? _T_10366_26 : _T_15490; // @[Mux.scala 46:16:@13718.4]
  assign _T_15493 = 6'h1a == _T_11317_50; // @[Mux.scala 46:19:@13719.4]
  assign _T_15494 = _T_15493 ? _T_10366_25 : _T_15492; // @[Mux.scala 46:16:@13720.4]
  assign _T_15495 = 6'h19 == _T_11317_50; // @[Mux.scala 46:19:@13721.4]
  assign _T_15496 = _T_15495 ? _T_10366_24 : _T_15494; // @[Mux.scala 46:16:@13722.4]
  assign _T_15497 = 6'h18 == _T_11317_50; // @[Mux.scala 46:19:@13723.4]
  assign _T_15498 = _T_15497 ? _T_10366_23 : _T_15496; // @[Mux.scala 46:16:@13724.4]
  assign _T_15499 = 6'h17 == _T_11317_50; // @[Mux.scala 46:19:@13725.4]
  assign _T_15500 = _T_15499 ? _T_10366_22 : _T_15498; // @[Mux.scala 46:16:@13726.4]
  assign _T_15501 = 6'h16 == _T_11317_50; // @[Mux.scala 46:19:@13727.4]
  assign _T_15502 = _T_15501 ? _T_10366_21 : _T_15500; // @[Mux.scala 46:16:@13728.4]
  assign _T_15503 = 6'h15 == _T_11317_50; // @[Mux.scala 46:19:@13729.4]
  assign _T_15504 = _T_15503 ? _T_10366_20 : _T_15502; // @[Mux.scala 46:16:@13730.4]
  assign _T_15505 = 6'h14 == _T_11317_50; // @[Mux.scala 46:19:@13731.4]
  assign _T_15506 = _T_15505 ? _T_10366_19 : _T_15504; // @[Mux.scala 46:16:@13732.4]
  assign _T_15507 = 6'h13 == _T_11317_50; // @[Mux.scala 46:19:@13733.4]
  assign _T_15508 = _T_15507 ? _T_10366_18 : _T_15506; // @[Mux.scala 46:16:@13734.4]
  assign _T_15509 = 6'h12 == _T_11317_50; // @[Mux.scala 46:19:@13735.4]
  assign _T_15510 = _T_15509 ? _T_10366_17 : _T_15508; // @[Mux.scala 46:16:@13736.4]
  assign _T_15511 = 6'h11 == _T_11317_50; // @[Mux.scala 46:19:@13737.4]
  assign _T_15512 = _T_15511 ? _T_10366_16 : _T_15510; // @[Mux.scala 46:16:@13738.4]
  assign _T_15513 = 6'h10 == _T_11317_50; // @[Mux.scala 46:19:@13739.4]
  assign _T_15514 = _T_15513 ? _T_10366_15 : _T_15512; // @[Mux.scala 46:16:@13740.4]
  assign _T_15515 = 6'hf == _T_11317_50; // @[Mux.scala 46:19:@13741.4]
  assign _T_15516 = _T_15515 ? _T_10366_14 : _T_15514; // @[Mux.scala 46:16:@13742.4]
  assign _T_15517 = 6'he == _T_11317_50; // @[Mux.scala 46:19:@13743.4]
  assign _T_15518 = _T_15517 ? _T_10366_13 : _T_15516; // @[Mux.scala 46:16:@13744.4]
  assign _T_15519 = 6'hd == _T_11317_50; // @[Mux.scala 46:19:@13745.4]
  assign _T_15520 = _T_15519 ? _T_10366_12 : _T_15518; // @[Mux.scala 46:16:@13746.4]
  assign _T_15521 = 6'hc == _T_11317_50; // @[Mux.scala 46:19:@13747.4]
  assign _T_15522 = _T_15521 ? _T_10366_11 : _T_15520; // @[Mux.scala 46:16:@13748.4]
  assign _T_15523 = 6'hb == _T_11317_50; // @[Mux.scala 46:19:@13749.4]
  assign _T_15524 = _T_15523 ? _T_10366_10 : _T_15522; // @[Mux.scala 46:16:@13750.4]
  assign _T_15525 = 6'ha == _T_11317_50; // @[Mux.scala 46:19:@13751.4]
  assign _T_15526 = _T_15525 ? _T_10366_9 : _T_15524; // @[Mux.scala 46:16:@13752.4]
  assign _T_15527 = 6'h9 == _T_11317_50; // @[Mux.scala 46:19:@13753.4]
  assign _T_15528 = _T_15527 ? _T_10366_8 : _T_15526; // @[Mux.scala 46:16:@13754.4]
  assign _T_15529 = 6'h8 == _T_11317_50; // @[Mux.scala 46:19:@13755.4]
  assign _T_15530 = _T_15529 ? _T_10366_7 : _T_15528; // @[Mux.scala 46:16:@13756.4]
  assign _T_15531 = 6'h7 == _T_11317_50; // @[Mux.scala 46:19:@13757.4]
  assign _T_15532 = _T_15531 ? _T_10366_6 : _T_15530; // @[Mux.scala 46:16:@13758.4]
  assign _T_15533 = 6'h6 == _T_11317_50; // @[Mux.scala 46:19:@13759.4]
  assign _T_15534 = _T_15533 ? _T_10366_5 : _T_15532; // @[Mux.scala 46:16:@13760.4]
  assign _T_15535 = 6'h5 == _T_11317_50; // @[Mux.scala 46:19:@13761.4]
  assign _T_15536 = _T_15535 ? _T_10366_4 : _T_15534; // @[Mux.scala 46:16:@13762.4]
  assign _T_15537 = 6'h4 == _T_11317_50; // @[Mux.scala 46:19:@13763.4]
  assign _T_15538 = _T_15537 ? _T_10366_3 : _T_15536; // @[Mux.scala 46:16:@13764.4]
  assign _T_15539 = 6'h3 == _T_11317_50; // @[Mux.scala 46:19:@13765.4]
  assign _T_15540 = _T_15539 ? _T_10366_2 : _T_15538; // @[Mux.scala 46:16:@13766.4]
  assign _T_15541 = 6'h2 == _T_11317_50; // @[Mux.scala 46:19:@13767.4]
  assign _T_15542 = _T_15541 ? _T_10366_1 : _T_15540; // @[Mux.scala 46:16:@13768.4]
  assign _T_15543 = 6'h1 == _T_11317_50; // @[Mux.scala 46:19:@13769.4]
  assign _T_15544 = _T_15543 ? _T_10366_0 : _T_15542; // @[Mux.scala 46:16:@13770.4]
  assign _T_15598 = 6'h34 == _T_11317_51; // @[Mux.scala 46:19:@13772.4]
  assign _T_15599 = _T_15598 ? _T_10366_51 : 8'h0; // @[Mux.scala 46:16:@13773.4]
  assign _T_15600 = 6'h33 == _T_11317_51; // @[Mux.scala 46:19:@13774.4]
  assign _T_15601 = _T_15600 ? _T_10366_50 : _T_15599; // @[Mux.scala 46:16:@13775.4]
  assign _T_15602 = 6'h32 == _T_11317_51; // @[Mux.scala 46:19:@13776.4]
  assign _T_15603 = _T_15602 ? _T_10366_49 : _T_15601; // @[Mux.scala 46:16:@13777.4]
  assign _T_15604 = 6'h31 == _T_11317_51; // @[Mux.scala 46:19:@13778.4]
  assign _T_15605 = _T_15604 ? _T_10366_48 : _T_15603; // @[Mux.scala 46:16:@13779.4]
  assign _T_15606 = 6'h30 == _T_11317_51; // @[Mux.scala 46:19:@13780.4]
  assign _T_15607 = _T_15606 ? _T_10366_47 : _T_15605; // @[Mux.scala 46:16:@13781.4]
  assign _T_15608 = 6'h2f == _T_11317_51; // @[Mux.scala 46:19:@13782.4]
  assign _T_15609 = _T_15608 ? _T_10366_46 : _T_15607; // @[Mux.scala 46:16:@13783.4]
  assign _T_15610 = 6'h2e == _T_11317_51; // @[Mux.scala 46:19:@13784.4]
  assign _T_15611 = _T_15610 ? _T_10366_45 : _T_15609; // @[Mux.scala 46:16:@13785.4]
  assign _T_15612 = 6'h2d == _T_11317_51; // @[Mux.scala 46:19:@13786.4]
  assign _T_15613 = _T_15612 ? _T_10366_44 : _T_15611; // @[Mux.scala 46:16:@13787.4]
  assign _T_15614 = 6'h2c == _T_11317_51; // @[Mux.scala 46:19:@13788.4]
  assign _T_15615 = _T_15614 ? _T_10366_43 : _T_15613; // @[Mux.scala 46:16:@13789.4]
  assign _T_15616 = 6'h2b == _T_11317_51; // @[Mux.scala 46:19:@13790.4]
  assign _T_15617 = _T_15616 ? _T_10366_42 : _T_15615; // @[Mux.scala 46:16:@13791.4]
  assign _T_15618 = 6'h2a == _T_11317_51; // @[Mux.scala 46:19:@13792.4]
  assign _T_15619 = _T_15618 ? _T_10366_41 : _T_15617; // @[Mux.scala 46:16:@13793.4]
  assign _T_15620 = 6'h29 == _T_11317_51; // @[Mux.scala 46:19:@13794.4]
  assign _T_15621 = _T_15620 ? _T_10366_40 : _T_15619; // @[Mux.scala 46:16:@13795.4]
  assign _T_15622 = 6'h28 == _T_11317_51; // @[Mux.scala 46:19:@13796.4]
  assign _T_15623 = _T_15622 ? _T_10366_39 : _T_15621; // @[Mux.scala 46:16:@13797.4]
  assign _T_15624 = 6'h27 == _T_11317_51; // @[Mux.scala 46:19:@13798.4]
  assign _T_15625 = _T_15624 ? _T_10366_38 : _T_15623; // @[Mux.scala 46:16:@13799.4]
  assign _T_15626 = 6'h26 == _T_11317_51; // @[Mux.scala 46:19:@13800.4]
  assign _T_15627 = _T_15626 ? _T_10366_37 : _T_15625; // @[Mux.scala 46:16:@13801.4]
  assign _T_15628 = 6'h25 == _T_11317_51; // @[Mux.scala 46:19:@13802.4]
  assign _T_15629 = _T_15628 ? _T_10366_36 : _T_15627; // @[Mux.scala 46:16:@13803.4]
  assign _T_15630 = 6'h24 == _T_11317_51; // @[Mux.scala 46:19:@13804.4]
  assign _T_15631 = _T_15630 ? _T_10366_35 : _T_15629; // @[Mux.scala 46:16:@13805.4]
  assign _T_15632 = 6'h23 == _T_11317_51; // @[Mux.scala 46:19:@13806.4]
  assign _T_15633 = _T_15632 ? _T_10366_34 : _T_15631; // @[Mux.scala 46:16:@13807.4]
  assign _T_15634 = 6'h22 == _T_11317_51; // @[Mux.scala 46:19:@13808.4]
  assign _T_15635 = _T_15634 ? _T_10366_33 : _T_15633; // @[Mux.scala 46:16:@13809.4]
  assign _T_15636 = 6'h21 == _T_11317_51; // @[Mux.scala 46:19:@13810.4]
  assign _T_15637 = _T_15636 ? _T_10366_32 : _T_15635; // @[Mux.scala 46:16:@13811.4]
  assign _T_15638 = 6'h20 == _T_11317_51; // @[Mux.scala 46:19:@13812.4]
  assign _T_15639 = _T_15638 ? _T_10366_31 : _T_15637; // @[Mux.scala 46:16:@13813.4]
  assign _T_15640 = 6'h1f == _T_11317_51; // @[Mux.scala 46:19:@13814.4]
  assign _T_15641 = _T_15640 ? _T_10366_30 : _T_15639; // @[Mux.scala 46:16:@13815.4]
  assign _T_15642 = 6'h1e == _T_11317_51; // @[Mux.scala 46:19:@13816.4]
  assign _T_15643 = _T_15642 ? _T_10366_29 : _T_15641; // @[Mux.scala 46:16:@13817.4]
  assign _T_15644 = 6'h1d == _T_11317_51; // @[Mux.scala 46:19:@13818.4]
  assign _T_15645 = _T_15644 ? _T_10366_28 : _T_15643; // @[Mux.scala 46:16:@13819.4]
  assign _T_15646 = 6'h1c == _T_11317_51; // @[Mux.scala 46:19:@13820.4]
  assign _T_15647 = _T_15646 ? _T_10366_27 : _T_15645; // @[Mux.scala 46:16:@13821.4]
  assign _T_15648 = 6'h1b == _T_11317_51; // @[Mux.scala 46:19:@13822.4]
  assign _T_15649 = _T_15648 ? _T_10366_26 : _T_15647; // @[Mux.scala 46:16:@13823.4]
  assign _T_15650 = 6'h1a == _T_11317_51; // @[Mux.scala 46:19:@13824.4]
  assign _T_15651 = _T_15650 ? _T_10366_25 : _T_15649; // @[Mux.scala 46:16:@13825.4]
  assign _T_15652 = 6'h19 == _T_11317_51; // @[Mux.scala 46:19:@13826.4]
  assign _T_15653 = _T_15652 ? _T_10366_24 : _T_15651; // @[Mux.scala 46:16:@13827.4]
  assign _T_15654 = 6'h18 == _T_11317_51; // @[Mux.scala 46:19:@13828.4]
  assign _T_15655 = _T_15654 ? _T_10366_23 : _T_15653; // @[Mux.scala 46:16:@13829.4]
  assign _T_15656 = 6'h17 == _T_11317_51; // @[Mux.scala 46:19:@13830.4]
  assign _T_15657 = _T_15656 ? _T_10366_22 : _T_15655; // @[Mux.scala 46:16:@13831.4]
  assign _T_15658 = 6'h16 == _T_11317_51; // @[Mux.scala 46:19:@13832.4]
  assign _T_15659 = _T_15658 ? _T_10366_21 : _T_15657; // @[Mux.scala 46:16:@13833.4]
  assign _T_15660 = 6'h15 == _T_11317_51; // @[Mux.scala 46:19:@13834.4]
  assign _T_15661 = _T_15660 ? _T_10366_20 : _T_15659; // @[Mux.scala 46:16:@13835.4]
  assign _T_15662 = 6'h14 == _T_11317_51; // @[Mux.scala 46:19:@13836.4]
  assign _T_15663 = _T_15662 ? _T_10366_19 : _T_15661; // @[Mux.scala 46:16:@13837.4]
  assign _T_15664 = 6'h13 == _T_11317_51; // @[Mux.scala 46:19:@13838.4]
  assign _T_15665 = _T_15664 ? _T_10366_18 : _T_15663; // @[Mux.scala 46:16:@13839.4]
  assign _T_15666 = 6'h12 == _T_11317_51; // @[Mux.scala 46:19:@13840.4]
  assign _T_15667 = _T_15666 ? _T_10366_17 : _T_15665; // @[Mux.scala 46:16:@13841.4]
  assign _T_15668 = 6'h11 == _T_11317_51; // @[Mux.scala 46:19:@13842.4]
  assign _T_15669 = _T_15668 ? _T_10366_16 : _T_15667; // @[Mux.scala 46:16:@13843.4]
  assign _T_15670 = 6'h10 == _T_11317_51; // @[Mux.scala 46:19:@13844.4]
  assign _T_15671 = _T_15670 ? _T_10366_15 : _T_15669; // @[Mux.scala 46:16:@13845.4]
  assign _T_15672 = 6'hf == _T_11317_51; // @[Mux.scala 46:19:@13846.4]
  assign _T_15673 = _T_15672 ? _T_10366_14 : _T_15671; // @[Mux.scala 46:16:@13847.4]
  assign _T_15674 = 6'he == _T_11317_51; // @[Mux.scala 46:19:@13848.4]
  assign _T_15675 = _T_15674 ? _T_10366_13 : _T_15673; // @[Mux.scala 46:16:@13849.4]
  assign _T_15676 = 6'hd == _T_11317_51; // @[Mux.scala 46:19:@13850.4]
  assign _T_15677 = _T_15676 ? _T_10366_12 : _T_15675; // @[Mux.scala 46:16:@13851.4]
  assign _T_15678 = 6'hc == _T_11317_51; // @[Mux.scala 46:19:@13852.4]
  assign _T_15679 = _T_15678 ? _T_10366_11 : _T_15677; // @[Mux.scala 46:16:@13853.4]
  assign _T_15680 = 6'hb == _T_11317_51; // @[Mux.scala 46:19:@13854.4]
  assign _T_15681 = _T_15680 ? _T_10366_10 : _T_15679; // @[Mux.scala 46:16:@13855.4]
  assign _T_15682 = 6'ha == _T_11317_51; // @[Mux.scala 46:19:@13856.4]
  assign _T_15683 = _T_15682 ? _T_10366_9 : _T_15681; // @[Mux.scala 46:16:@13857.4]
  assign _T_15684 = 6'h9 == _T_11317_51; // @[Mux.scala 46:19:@13858.4]
  assign _T_15685 = _T_15684 ? _T_10366_8 : _T_15683; // @[Mux.scala 46:16:@13859.4]
  assign _T_15686 = 6'h8 == _T_11317_51; // @[Mux.scala 46:19:@13860.4]
  assign _T_15687 = _T_15686 ? _T_10366_7 : _T_15685; // @[Mux.scala 46:16:@13861.4]
  assign _T_15688 = 6'h7 == _T_11317_51; // @[Mux.scala 46:19:@13862.4]
  assign _T_15689 = _T_15688 ? _T_10366_6 : _T_15687; // @[Mux.scala 46:16:@13863.4]
  assign _T_15690 = 6'h6 == _T_11317_51; // @[Mux.scala 46:19:@13864.4]
  assign _T_15691 = _T_15690 ? _T_10366_5 : _T_15689; // @[Mux.scala 46:16:@13865.4]
  assign _T_15692 = 6'h5 == _T_11317_51; // @[Mux.scala 46:19:@13866.4]
  assign _T_15693 = _T_15692 ? _T_10366_4 : _T_15691; // @[Mux.scala 46:16:@13867.4]
  assign _T_15694 = 6'h4 == _T_11317_51; // @[Mux.scala 46:19:@13868.4]
  assign _T_15695 = _T_15694 ? _T_10366_3 : _T_15693; // @[Mux.scala 46:16:@13869.4]
  assign _T_15696 = 6'h3 == _T_11317_51; // @[Mux.scala 46:19:@13870.4]
  assign _T_15697 = _T_15696 ? _T_10366_2 : _T_15695; // @[Mux.scala 46:16:@13871.4]
  assign _T_15698 = 6'h2 == _T_11317_51; // @[Mux.scala 46:19:@13872.4]
  assign _T_15699 = _T_15698 ? _T_10366_1 : _T_15697; // @[Mux.scala 46:16:@13873.4]
  assign _T_15700 = 6'h1 == _T_11317_51; // @[Mux.scala 46:19:@13874.4]
  assign _T_15701 = _T_15700 ? _T_10366_0 : _T_15699; // @[Mux.scala 46:16:@13875.4]
  assign _T_15756 = 6'h35 == _T_11317_52; // @[Mux.scala 46:19:@13877.4]
  assign _T_15757 = _T_15756 ? _T_10366_52 : 8'h0; // @[Mux.scala 46:16:@13878.4]
  assign _T_15758 = 6'h34 == _T_11317_52; // @[Mux.scala 46:19:@13879.4]
  assign _T_15759 = _T_15758 ? _T_10366_51 : _T_15757; // @[Mux.scala 46:16:@13880.4]
  assign _T_15760 = 6'h33 == _T_11317_52; // @[Mux.scala 46:19:@13881.4]
  assign _T_15761 = _T_15760 ? _T_10366_50 : _T_15759; // @[Mux.scala 46:16:@13882.4]
  assign _T_15762 = 6'h32 == _T_11317_52; // @[Mux.scala 46:19:@13883.4]
  assign _T_15763 = _T_15762 ? _T_10366_49 : _T_15761; // @[Mux.scala 46:16:@13884.4]
  assign _T_15764 = 6'h31 == _T_11317_52; // @[Mux.scala 46:19:@13885.4]
  assign _T_15765 = _T_15764 ? _T_10366_48 : _T_15763; // @[Mux.scala 46:16:@13886.4]
  assign _T_15766 = 6'h30 == _T_11317_52; // @[Mux.scala 46:19:@13887.4]
  assign _T_15767 = _T_15766 ? _T_10366_47 : _T_15765; // @[Mux.scala 46:16:@13888.4]
  assign _T_15768 = 6'h2f == _T_11317_52; // @[Mux.scala 46:19:@13889.4]
  assign _T_15769 = _T_15768 ? _T_10366_46 : _T_15767; // @[Mux.scala 46:16:@13890.4]
  assign _T_15770 = 6'h2e == _T_11317_52; // @[Mux.scala 46:19:@13891.4]
  assign _T_15771 = _T_15770 ? _T_10366_45 : _T_15769; // @[Mux.scala 46:16:@13892.4]
  assign _T_15772 = 6'h2d == _T_11317_52; // @[Mux.scala 46:19:@13893.4]
  assign _T_15773 = _T_15772 ? _T_10366_44 : _T_15771; // @[Mux.scala 46:16:@13894.4]
  assign _T_15774 = 6'h2c == _T_11317_52; // @[Mux.scala 46:19:@13895.4]
  assign _T_15775 = _T_15774 ? _T_10366_43 : _T_15773; // @[Mux.scala 46:16:@13896.4]
  assign _T_15776 = 6'h2b == _T_11317_52; // @[Mux.scala 46:19:@13897.4]
  assign _T_15777 = _T_15776 ? _T_10366_42 : _T_15775; // @[Mux.scala 46:16:@13898.4]
  assign _T_15778 = 6'h2a == _T_11317_52; // @[Mux.scala 46:19:@13899.4]
  assign _T_15779 = _T_15778 ? _T_10366_41 : _T_15777; // @[Mux.scala 46:16:@13900.4]
  assign _T_15780 = 6'h29 == _T_11317_52; // @[Mux.scala 46:19:@13901.4]
  assign _T_15781 = _T_15780 ? _T_10366_40 : _T_15779; // @[Mux.scala 46:16:@13902.4]
  assign _T_15782 = 6'h28 == _T_11317_52; // @[Mux.scala 46:19:@13903.4]
  assign _T_15783 = _T_15782 ? _T_10366_39 : _T_15781; // @[Mux.scala 46:16:@13904.4]
  assign _T_15784 = 6'h27 == _T_11317_52; // @[Mux.scala 46:19:@13905.4]
  assign _T_15785 = _T_15784 ? _T_10366_38 : _T_15783; // @[Mux.scala 46:16:@13906.4]
  assign _T_15786 = 6'h26 == _T_11317_52; // @[Mux.scala 46:19:@13907.4]
  assign _T_15787 = _T_15786 ? _T_10366_37 : _T_15785; // @[Mux.scala 46:16:@13908.4]
  assign _T_15788 = 6'h25 == _T_11317_52; // @[Mux.scala 46:19:@13909.4]
  assign _T_15789 = _T_15788 ? _T_10366_36 : _T_15787; // @[Mux.scala 46:16:@13910.4]
  assign _T_15790 = 6'h24 == _T_11317_52; // @[Mux.scala 46:19:@13911.4]
  assign _T_15791 = _T_15790 ? _T_10366_35 : _T_15789; // @[Mux.scala 46:16:@13912.4]
  assign _T_15792 = 6'h23 == _T_11317_52; // @[Mux.scala 46:19:@13913.4]
  assign _T_15793 = _T_15792 ? _T_10366_34 : _T_15791; // @[Mux.scala 46:16:@13914.4]
  assign _T_15794 = 6'h22 == _T_11317_52; // @[Mux.scala 46:19:@13915.4]
  assign _T_15795 = _T_15794 ? _T_10366_33 : _T_15793; // @[Mux.scala 46:16:@13916.4]
  assign _T_15796 = 6'h21 == _T_11317_52; // @[Mux.scala 46:19:@13917.4]
  assign _T_15797 = _T_15796 ? _T_10366_32 : _T_15795; // @[Mux.scala 46:16:@13918.4]
  assign _T_15798 = 6'h20 == _T_11317_52; // @[Mux.scala 46:19:@13919.4]
  assign _T_15799 = _T_15798 ? _T_10366_31 : _T_15797; // @[Mux.scala 46:16:@13920.4]
  assign _T_15800 = 6'h1f == _T_11317_52; // @[Mux.scala 46:19:@13921.4]
  assign _T_15801 = _T_15800 ? _T_10366_30 : _T_15799; // @[Mux.scala 46:16:@13922.4]
  assign _T_15802 = 6'h1e == _T_11317_52; // @[Mux.scala 46:19:@13923.4]
  assign _T_15803 = _T_15802 ? _T_10366_29 : _T_15801; // @[Mux.scala 46:16:@13924.4]
  assign _T_15804 = 6'h1d == _T_11317_52; // @[Mux.scala 46:19:@13925.4]
  assign _T_15805 = _T_15804 ? _T_10366_28 : _T_15803; // @[Mux.scala 46:16:@13926.4]
  assign _T_15806 = 6'h1c == _T_11317_52; // @[Mux.scala 46:19:@13927.4]
  assign _T_15807 = _T_15806 ? _T_10366_27 : _T_15805; // @[Mux.scala 46:16:@13928.4]
  assign _T_15808 = 6'h1b == _T_11317_52; // @[Mux.scala 46:19:@13929.4]
  assign _T_15809 = _T_15808 ? _T_10366_26 : _T_15807; // @[Mux.scala 46:16:@13930.4]
  assign _T_15810 = 6'h1a == _T_11317_52; // @[Mux.scala 46:19:@13931.4]
  assign _T_15811 = _T_15810 ? _T_10366_25 : _T_15809; // @[Mux.scala 46:16:@13932.4]
  assign _T_15812 = 6'h19 == _T_11317_52; // @[Mux.scala 46:19:@13933.4]
  assign _T_15813 = _T_15812 ? _T_10366_24 : _T_15811; // @[Mux.scala 46:16:@13934.4]
  assign _T_15814 = 6'h18 == _T_11317_52; // @[Mux.scala 46:19:@13935.4]
  assign _T_15815 = _T_15814 ? _T_10366_23 : _T_15813; // @[Mux.scala 46:16:@13936.4]
  assign _T_15816 = 6'h17 == _T_11317_52; // @[Mux.scala 46:19:@13937.4]
  assign _T_15817 = _T_15816 ? _T_10366_22 : _T_15815; // @[Mux.scala 46:16:@13938.4]
  assign _T_15818 = 6'h16 == _T_11317_52; // @[Mux.scala 46:19:@13939.4]
  assign _T_15819 = _T_15818 ? _T_10366_21 : _T_15817; // @[Mux.scala 46:16:@13940.4]
  assign _T_15820 = 6'h15 == _T_11317_52; // @[Mux.scala 46:19:@13941.4]
  assign _T_15821 = _T_15820 ? _T_10366_20 : _T_15819; // @[Mux.scala 46:16:@13942.4]
  assign _T_15822 = 6'h14 == _T_11317_52; // @[Mux.scala 46:19:@13943.4]
  assign _T_15823 = _T_15822 ? _T_10366_19 : _T_15821; // @[Mux.scala 46:16:@13944.4]
  assign _T_15824 = 6'h13 == _T_11317_52; // @[Mux.scala 46:19:@13945.4]
  assign _T_15825 = _T_15824 ? _T_10366_18 : _T_15823; // @[Mux.scala 46:16:@13946.4]
  assign _T_15826 = 6'h12 == _T_11317_52; // @[Mux.scala 46:19:@13947.4]
  assign _T_15827 = _T_15826 ? _T_10366_17 : _T_15825; // @[Mux.scala 46:16:@13948.4]
  assign _T_15828 = 6'h11 == _T_11317_52; // @[Mux.scala 46:19:@13949.4]
  assign _T_15829 = _T_15828 ? _T_10366_16 : _T_15827; // @[Mux.scala 46:16:@13950.4]
  assign _T_15830 = 6'h10 == _T_11317_52; // @[Mux.scala 46:19:@13951.4]
  assign _T_15831 = _T_15830 ? _T_10366_15 : _T_15829; // @[Mux.scala 46:16:@13952.4]
  assign _T_15832 = 6'hf == _T_11317_52; // @[Mux.scala 46:19:@13953.4]
  assign _T_15833 = _T_15832 ? _T_10366_14 : _T_15831; // @[Mux.scala 46:16:@13954.4]
  assign _T_15834 = 6'he == _T_11317_52; // @[Mux.scala 46:19:@13955.4]
  assign _T_15835 = _T_15834 ? _T_10366_13 : _T_15833; // @[Mux.scala 46:16:@13956.4]
  assign _T_15836 = 6'hd == _T_11317_52; // @[Mux.scala 46:19:@13957.4]
  assign _T_15837 = _T_15836 ? _T_10366_12 : _T_15835; // @[Mux.scala 46:16:@13958.4]
  assign _T_15838 = 6'hc == _T_11317_52; // @[Mux.scala 46:19:@13959.4]
  assign _T_15839 = _T_15838 ? _T_10366_11 : _T_15837; // @[Mux.scala 46:16:@13960.4]
  assign _T_15840 = 6'hb == _T_11317_52; // @[Mux.scala 46:19:@13961.4]
  assign _T_15841 = _T_15840 ? _T_10366_10 : _T_15839; // @[Mux.scala 46:16:@13962.4]
  assign _T_15842 = 6'ha == _T_11317_52; // @[Mux.scala 46:19:@13963.4]
  assign _T_15843 = _T_15842 ? _T_10366_9 : _T_15841; // @[Mux.scala 46:16:@13964.4]
  assign _T_15844 = 6'h9 == _T_11317_52; // @[Mux.scala 46:19:@13965.4]
  assign _T_15845 = _T_15844 ? _T_10366_8 : _T_15843; // @[Mux.scala 46:16:@13966.4]
  assign _T_15846 = 6'h8 == _T_11317_52; // @[Mux.scala 46:19:@13967.4]
  assign _T_15847 = _T_15846 ? _T_10366_7 : _T_15845; // @[Mux.scala 46:16:@13968.4]
  assign _T_15848 = 6'h7 == _T_11317_52; // @[Mux.scala 46:19:@13969.4]
  assign _T_15849 = _T_15848 ? _T_10366_6 : _T_15847; // @[Mux.scala 46:16:@13970.4]
  assign _T_15850 = 6'h6 == _T_11317_52; // @[Mux.scala 46:19:@13971.4]
  assign _T_15851 = _T_15850 ? _T_10366_5 : _T_15849; // @[Mux.scala 46:16:@13972.4]
  assign _T_15852 = 6'h5 == _T_11317_52; // @[Mux.scala 46:19:@13973.4]
  assign _T_15853 = _T_15852 ? _T_10366_4 : _T_15851; // @[Mux.scala 46:16:@13974.4]
  assign _T_15854 = 6'h4 == _T_11317_52; // @[Mux.scala 46:19:@13975.4]
  assign _T_15855 = _T_15854 ? _T_10366_3 : _T_15853; // @[Mux.scala 46:16:@13976.4]
  assign _T_15856 = 6'h3 == _T_11317_52; // @[Mux.scala 46:19:@13977.4]
  assign _T_15857 = _T_15856 ? _T_10366_2 : _T_15855; // @[Mux.scala 46:16:@13978.4]
  assign _T_15858 = 6'h2 == _T_11317_52; // @[Mux.scala 46:19:@13979.4]
  assign _T_15859 = _T_15858 ? _T_10366_1 : _T_15857; // @[Mux.scala 46:16:@13980.4]
  assign _T_15860 = 6'h1 == _T_11317_52; // @[Mux.scala 46:19:@13981.4]
  assign _T_15861 = _T_15860 ? _T_10366_0 : _T_15859; // @[Mux.scala 46:16:@13982.4]
  assign _T_15917 = 6'h36 == _T_11317_53; // @[Mux.scala 46:19:@13984.4]
  assign _T_15918 = _T_15917 ? _T_10366_53 : 8'h0; // @[Mux.scala 46:16:@13985.4]
  assign _T_15919 = 6'h35 == _T_11317_53; // @[Mux.scala 46:19:@13986.4]
  assign _T_15920 = _T_15919 ? _T_10366_52 : _T_15918; // @[Mux.scala 46:16:@13987.4]
  assign _T_15921 = 6'h34 == _T_11317_53; // @[Mux.scala 46:19:@13988.4]
  assign _T_15922 = _T_15921 ? _T_10366_51 : _T_15920; // @[Mux.scala 46:16:@13989.4]
  assign _T_15923 = 6'h33 == _T_11317_53; // @[Mux.scala 46:19:@13990.4]
  assign _T_15924 = _T_15923 ? _T_10366_50 : _T_15922; // @[Mux.scala 46:16:@13991.4]
  assign _T_15925 = 6'h32 == _T_11317_53; // @[Mux.scala 46:19:@13992.4]
  assign _T_15926 = _T_15925 ? _T_10366_49 : _T_15924; // @[Mux.scala 46:16:@13993.4]
  assign _T_15927 = 6'h31 == _T_11317_53; // @[Mux.scala 46:19:@13994.4]
  assign _T_15928 = _T_15927 ? _T_10366_48 : _T_15926; // @[Mux.scala 46:16:@13995.4]
  assign _T_15929 = 6'h30 == _T_11317_53; // @[Mux.scala 46:19:@13996.4]
  assign _T_15930 = _T_15929 ? _T_10366_47 : _T_15928; // @[Mux.scala 46:16:@13997.4]
  assign _T_15931 = 6'h2f == _T_11317_53; // @[Mux.scala 46:19:@13998.4]
  assign _T_15932 = _T_15931 ? _T_10366_46 : _T_15930; // @[Mux.scala 46:16:@13999.4]
  assign _T_15933 = 6'h2e == _T_11317_53; // @[Mux.scala 46:19:@14000.4]
  assign _T_15934 = _T_15933 ? _T_10366_45 : _T_15932; // @[Mux.scala 46:16:@14001.4]
  assign _T_15935 = 6'h2d == _T_11317_53; // @[Mux.scala 46:19:@14002.4]
  assign _T_15936 = _T_15935 ? _T_10366_44 : _T_15934; // @[Mux.scala 46:16:@14003.4]
  assign _T_15937 = 6'h2c == _T_11317_53; // @[Mux.scala 46:19:@14004.4]
  assign _T_15938 = _T_15937 ? _T_10366_43 : _T_15936; // @[Mux.scala 46:16:@14005.4]
  assign _T_15939 = 6'h2b == _T_11317_53; // @[Mux.scala 46:19:@14006.4]
  assign _T_15940 = _T_15939 ? _T_10366_42 : _T_15938; // @[Mux.scala 46:16:@14007.4]
  assign _T_15941 = 6'h2a == _T_11317_53; // @[Mux.scala 46:19:@14008.4]
  assign _T_15942 = _T_15941 ? _T_10366_41 : _T_15940; // @[Mux.scala 46:16:@14009.4]
  assign _T_15943 = 6'h29 == _T_11317_53; // @[Mux.scala 46:19:@14010.4]
  assign _T_15944 = _T_15943 ? _T_10366_40 : _T_15942; // @[Mux.scala 46:16:@14011.4]
  assign _T_15945 = 6'h28 == _T_11317_53; // @[Mux.scala 46:19:@14012.4]
  assign _T_15946 = _T_15945 ? _T_10366_39 : _T_15944; // @[Mux.scala 46:16:@14013.4]
  assign _T_15947 = 6'h27 == _T_11317_53; // @[Mux.scala 46:19:@14014.4]
  assign _T_15948 = _T_15947 ? _T_10366_38 : _T_15946; // @[Mux.scala 46:16:@14015.4]
  assign _T_15949 = 6'h26 == _T_11317_53; // @[Mux.scala 46:19:@14016.4]
  assign _T_15950 = _T_15949 ? _T_10366_37 : _T_15948; // @[Mux.scala 46:16:@14017.4]
  assign _T_15951 = 6'h25 == _T_11317_53; // @[Mux.scala 46:19:@14018.4]
  assign _T_15952 = _T_15951 ? _T_10366_36 : _T_15950; // @[Mux.scala 46:16:@14019.4]
  assign _T_15953 = 6'h24 == _T_11317_53; // @[Mux.scala 46:19:@14020.4]
  assign _T_15954 = _T_15953 ? _T_10366_35 : _T_15952; // @[Mux.scala 46:16:@14021.4]
  assign _T_15955 = 6'h23 == _T_11317_53; // @[Mux.scala 46:19:@14022.4]
  assign _T_15956 = _T_15955 ? _T_10366_34 : _T_15954; // @[Mux.scala 46:16:@14023.4]
  assign _T_15957 = 6'h22 == _T_11317_53; // @[Mux.scala 46:19:@14024.4]
  assign _T_15958 = _T_15957 ? _T_10366_33 : _T_15956; // @[Mux.scala 46:16:@14025.4]
  assign _T_15959 = 6'h21 == _T_11317_53; // @[Mux.scala 46:19:@14026.4]
  assign _T_15960 = _T_15959 ? _T_10366_32 : _T_15958; // @[Mux.scala 46:16:@14027.4]
  assign _T_15961 = 6'h20 == _T_11317_53; // @[Mux.scala 46:19:@14028.4]
  assign _T_15962 = _T_15961 ? _T_10366_31 : _T_15960; // @[Mux.scala 46:16:@14029.4]
  assign _T_15963 = 6'h1f == _T_11317_53; // @[Mux.scala 46:19:@14030.4]
  assign _T_15964 = _T_15963 ? _T_10366_30 : _T_15962; // @[Mux.scala 46:16:@14031.4]
  assign _T_15965 = 6'h1e == _T_11317_53; // @[Mux.scala 46:19:@14032.4]
  assign _T_15966 = _T_15965 ? _T_10366_29 : _T_15964; // @[Mux.scala 46:16:@14033.4]
  assign _T_15967 = 6'h1d == _T_11317_53; // @[Mux.scala 46:19:@14034.4]
  assign _T_15968 = _T_15967 ? _T_10366_28 : _T_15966; // @[Mux.scala 46:16:@14035.4]
  assign _T_15969 = 6'h1c == _T_11317_53; // @[Mux.scala 46:19:@14036.4]
  assign _T_15970 = _T_15969 ? _T_10366_27 : _T_15968; // @[Mux.scala 46:16:@14037.4]
  assign _T_15971 = 6'h1b == _T_11317_53; // @[Mux.scala 46:19:@14038.4]
  assign _T_15972 = _T_15971 ? _T_10366_26 : _T_15970; // @[Mux.scala 46:16:@14039.4]
  assign _T_15973 = 6'h1a == _T_11317_53; // @[Mux.scala 46:19:@14040.4]
  assign _T_15974 = _T_15973 ? _T_10366_25 : _T_15972; // @[Mux.scala 46:16:@14041.4]
  assign _T_15975 = 6'h19 == _T_11317_53; // @[Mux.scala 46:19:@14042.4]
  assign _T_15976 = _T_15975 ? _T_10366_24 : _T_15974; // @[Mux.scala 46:16:@14043.4]
  assign _T_15977 = 6'h18 == _T_11317_53; // @[Mux.scala 46:19:@14044.4]
  assign _T_15978 = _T_15977 ? _T_10366_23 : _T_15976; // @[Mux.scala 46:16:@14045.4]
  assign _T_15979 = 6'h17 == _T_11317_53; // @[Mux.scala 46:19:@14046.4]
  assign _T_15980 = _T_15979 ? _T_10366_22 : _T_15978; // @[Mux.scala 46:16:@14047.4]
  assign _T_15981 = 6'h16 == _T_11317_53; // @[Mux.scala 46:19:@14048.4]
  assign _T_15982 = _T_15981 ? _T_10366_21 : _T_15980; // @[Mux.scala 46:16:@14049.4]
  assign _T_15983 = 6'h15 == _T_11317_53; // @[Mux.scala 46:19:@14050.4]
  assign _T_15984 = _T_15983 ? _T_10366_20 : _T_15982; // @[Mux.scala 46:16:@14051.4]
  assign _T_15985 = 6'h14 == _T_11317_53; // @[Mux.scala 46:19:@14052.4]
  assign _T_15986 = _T_15985 ? _T_10366_19 : _T_15984; // @[Mux.scala 46:16:@14053.4]
  assign _T_15987 = 6'h13 == _T_11317_53; // @[Mux.scala 46:19:@14054.4]
  assign _T_15988 = _T_15987 ? _T_10366_18 : _T_15986; // @[Mux.scala 46:16:@14055.4]
  assign _T_15989 = 6'h12 == _T_11317_53; // @[Mux.scala 46:19:@14056.4]
  assign _T_15990 = _T_15989 ? _T_10366_17 : _T_15988; // @[Mux.scala 46:16:@14057.4]
  assign _T_15991 = 6'h11 == _T_11317_53; // @[Mux.scala 46:19:@14058.4]
  assign _T_15992 = _T_15991 ? _T_10366_16 : _T_15990; // @[Mux.scala 46:16:@14059.4]
  assign _T_15993 = 6'h10 == _T_11317_53; // @[Mux.scala 46:19:@14060.4]
  assign _T_15994 = _T_15993 ? _T_10366_15 : _T_15992; // @[Mux.scala 46:16:@14061.4]
  assign _T_15995 = 6'hf == _T_11317_53; // @[Mux.scala 46:19:@14062.4]
  assign _T_15996 = _T_15995 ? _T_10366_14 : _T_15994; // @[Mux.scala 46:16:@14063.4]
  assign _T_15997 = 6'he == _T_11317_53; // @[Mux.scala 46:19:@14064.4]
  assign _T_15998 = _T_15997 ? _T_10366_13 : _T_15996; // @[Mux.scala 46:16:@14065.4]
  assign _T_15999 = 6'hd == _T_11317_53; // @[Mux.scala 46:19:@14066.4]
  assign _T_16000 = _T_15999 ? _T_10366_12 : _T_15998; // @[Mux.scala 46:16:@14067.4]
  assign _T_16001 = 6'hc == _T_11317_53; // @[Mux.scala 46:19:@14068.4]
  assign _T_16002 = _T_16001 ? _T_10366_11 : _T_16000; // @[Mux.scala 46:16:@14069.4]
  assign _T_16003 = 6'hb == _T_11317_53; // @[Mux.scala 46:19:@14070.4]
  assign _T_16004 = _T_16003 ? _T_10366_10 : _T_16002; // @[Mux.scala 46:16:@14071.4]
  assign _T_16005 = 6'ha == _T_11317_53; // @[Mux.scala 46:19:@14072.4]
  assign _T_16006 = _T_16005 ? _T_10366_9 : _T_16004; // @[Mux.scala 46:16:@14073.4]
  assign _T_16007 = 6'h9 == _T_11317_53; // @[Mux.scala 46:19:@14074.4]
  assign _T_16008 = _T_16007 ? _T_10366_8 : _T_16006; // @[Mux.scala 46:16:@14075.4]
  assign _T_16009 = 6'h8 == _T_11317_53; // @[Mux.scala 46:19:@14076.4]
  assign _T_16010 = _T_16009 ? _T_10366_7 : _T_16008; // @[Mux.scala 46:16:@14077.4]
  assign _T_16011 = 6'h7 == _T_11317_53; // @[Mux.scala 46:19:@14078.4]
  assign _T_16012 = _T_16011 ? _T_10366_6 : _T_16010; // @[Mux.scala 46:16:@14079.4]
  assign _T_16013 = 6'h6 == _T_11317_53; // @[Mux.scala 46:19:@14080.4]
  assign _T_16014 = _T_16013 ? _T_10366_5 : _T_16012; // @[Mux.scala 46:16:@14081.4]
  assign _T_16015 = 6'h5 == _T_11317_53; // @[Mux.scala 46:19:@14082.4]
  assign _T_16016 = _T_16015 ? _T_10366_4 : _T_16014; // @[Mux.scala 46:16:@14083.4]
  assign _T_16017 = 6'h4 == _T_11317_53; // @[Mux.scala 46:19:@14084.4]
  assign _T_16018 = _T_16017 ? _T_10366_3 : _T_16016; // @[Mux.scala 46:16:@14085.4]
  assign _T_16019 = 6'h3 == _T_11317_53; // @[Mux.scala 46:19:@14086.4]
  assign _T_16020 = _T_16019 ? _T_10366_2 : _T_16018; // @[Mux.scala 46:16:@14087.4]
  assign _T_16021 = 6'h2 == _T_11317_53; // @[Mux.scala 46:19:@14088.4]
  assign _T_16022 = _T_16021 ? _T_10366_1 : _T_16020; // @[Mux.scala 46:16:@14089.4]
  assign _T_16023 = 6'h1 == _T_11317_53; // @[Mux.scala 46:19:@14090.4]
  assign _T_16024 = _T_16023 ? _T_10366_0 : _T_16022; // @[Mux.scala 46:16:@14091.4]
  assign _T_16081 = 6'h37 == _T_11317_54; // @[Mux.scala 46:19:@14093.4]
  assign _T_16082 = _T_16081 ? _T_10366_54 : 8'h0; // @[Mux.scala 46:16:@14094.4]
  assign _T_16083 = 6'h36 == _T_11317_54; // @[Mux.scala 46:19:@14095.4]
  assign _T_16084 = _T_16083 ? _T_10366_53 : _T_16082; // @[Mux.scala 46:16:@14096.4]
  assign _T_16085 = 6'h35 == _T_11317_54; // @[Mux.scala 46:19:@14097.4]
  assign _T_16086 = _T_16085 ? _T_10366_52 : _T_16084; // @[Mux.scala 46:16:@14098.4]
  assign _T_16087 = 6'h34 == _T_11317_54; // @[Mux.scala 46:19:@14099.4]
  assign _T_16088 = _T_16087 ? _T_10366_51 : _T_16086; // @[Mux.scala 46:16:@14100.4]
  assign _T_16089 = 6'h33 == _T_11317_54; // @[Mux.scala 46:19:@14101.4]
  assign _T_16090 = _T_16089 ? _T_10366_50 : _T_16088; // @[Mux.scala 46:16:@14102.4]
  assign _T_16091 = 6'h32 == _T_11317_54; // @[Mux.scala 46:19:@14103.4]
  assign _T_16092 = _T_16091 ? _T_10366_49 : _T_16090; // @[Mux.scala 46:16:@14104.4]
  assign _T_16093 = 6'h31 == _T_11317_54; // @[Mux.scala 46:19:@14105.4]
  assign _T_16094 = _T_16093 ? _T_10366_48 : _T_16092; // @[Mux.scala 46:16:@14106.4]
  assign _T_16095 = 6'h30 == _T_11317_54; // @[Mux.scala 46:19:@14107.4]
  assign _T_16096 = _T_16095 ? _T_10366_47 : _T_16094; // @[Mux.scala 46:16:@14108.4]
  assign _T_16097 = 6'h2f == _T_11317_54; // @[Mux.scala 46:19:@14109.4]
  assign _T_16098 = _T_16097 ? _T_10366_46 : _T_16096; // @[Mux.scala 46:16:@14110.4]
  assign _T_16099 = 6'h2e == _T_11317_54; // @[Mux.scala 46:19:@14111.4]
  assign _T_16100 = _T_16099 ? _T_10366_45 : _T_16098; // @[Mux.scala 46:16:@14112.4]
  assign _T_16101 = 6'h2d == _T_11317_54; // @[Mux.scala 46:19:@14113.4]
  assign _T_16102 = _T_16101 ? _T_10366_44 : _T_16100; // @[Mux.scala 46:16:@14114.4]
  assign _T_16103 = 6'h2c == _T_11317_54; // @[Mux.scala 46:19:@14115.4]
  assign _T_16104 = _T_16103 ? _T_10366_43 : _T_16102; // @[Mux.scala 46:16:@14116.4]
  assign _T_16105 = 6'h2b == _T_11317_54; // @[Mux.scala 46:19:@14117.4]
  assign _T_16106 = _T_16105 ? _T_10366_42 : _T_16104; // @[Mux.scala 46:16:@14118.4]
  assign _T_16107 = 6'h2a == _T_11317_54; // @[Mux.scala 46:19:@14119.4]
  assign _T_16108 = _T_16107 ? _T_10366_41 : _T_16106; // @[Mux.scala 46:16:@14120.4]
  assign _T_16109 = 6'h29 == _T_11317_54; // @[Mux.scala 46:19:@14121.4]
  assign _T_16110 = _T_16109 ? _T_10366_40 : _T_16108; // @[Mux.scala 46:16:@14122.4]
  assign _T_16111 = 6'h28 == _T_11317_54; // @[Mux.scala 46:19:@14123.4]
  assign _T_16112 = _T_16111 ? _T_10366_39 : _T_16110; // @[Mux.scala 46:16:@14124.4]
  assign _T_16113 = 6'h27 == _T_11317_54; // @[Mux.scala 46:19:@14125.4]
  assign _T_16114 = _T_16113 ? _T_10366_38 : _T_16112; // @[Mux.scala 46:16:@14126.4]
  assign _T_16115 = 6'h26 == _T_11317_54; // @[Mux.scala 46:19:@14127.4]
  assign _T_16116 = _T_16115 ? _T_10366_37 : _T_16114; // @[Mux.scala 46:16:@14128.4]
  assign _T_16117 = 6'h25 == _T_11317_54; // @[Mux.scala 46:19:@14129.4]
  assign _T_16118 = _T_16117 ? _T_10366_36 : _T_16116; // @[Mux.scala 46:16:@14130.4]
  assign _T_16119 = 6'h24 == _T_11317_54; // @[Mux.scala 46:19:@14131.4]
  assign _T_16120 = _T_16119 ? _T_10366_35 : _T_16118; // @[Mux.scala 46:16:@14132.4]
  assign _T_16121 = 6'h23 == _T_11317_54; // @[Mux.scala 46:19:@14133.4]
  assign _T_16122 = _T_16121 ? _T_10366_34 : _T_16120; // @[Mux.scala 46:16:@14134.4]
  assign _T_16123 = 6'h22 == _T_11317_54; // @[Mux.scala 46:19:@14135.4]
  assign _T_16124 = _T_16123 ? _T_10366_33 : _T_16122; // @[Mux.scala 46:16:@14136.4]
  assign _T_16125 = 6'h21 == _T_11317_54; // @[Mux.scala 46:19:@14137.4]
  assign _T_16126 = _T_16125 ? _T_10366_32 : _T_16124; // @[Mux.scala 46:16:@14138.4]
  assign _T_16127 = 6'h20 == _T_11317_54; // @[Mux.scala 46:19:@14139.4]
  assign _T_16128 = _T_16127 ? _T_10366_31 : _T_16126; // @[Mux.scala 46:16:@14140.4]
  assign _T_16129 = 6'h1f == _T_11317_54; // @[Mux.scala 46:19:@14141.4]
  assign _T_16130 = _T_16129 ? _T_10366_30 : _T_16128; // @[Mux.scala 46:16:@14142.4]
  assign _T_16131 = 6'h1e == _T_11317_54; // @[Mux.scala 46:19:@14143.4]
  assign _T_16132 = _T_16131 ? _T_10366_29 : _T_16130; // @[Mux.scala 46:16:@14144.4]
  assign _T_16133 = 6'h1d == _T_11317_54; // @[Mux.scala 46:19:@14145.4]
  assign _T_16134 = _T_16133 ? _T_10366_28 : _T_16132; // @[Mux.scala 46:16:@14146.4]
  assign _T_16135 = 6'h1c == _T_11317_54; // @[Mux.scala 46:19:@14147.4]
  assign _T_16136 = _T_16135 ? _T_10366_27 : _T_16134; // @[Mux.scala 46:16:@14148.4]
  assign _T_16137 = 6'h1b == _T_11317_54; // @[Mux.scala 46:19:@14149.4]
  assign _T_16138 = _T_16137 ? _T_10366_26 : _T_16136; // @[Mux.scala 46:16:@14150.4]
  assign _T_16139 = 6'h1a == _T_11317_54; // @[Mux.scala 46:19:@14151.4]
  assign _T_16140 = _T_16139 ? _T_10366_25 : _T_16138; // @[Mux.scala 46:16:@14152.4]
  assign _T_16141 = 6'h19 == _T_11317_54; // @[Mux.scala 46:19:@14153.4]
  assign _T_16142 = _T_16141 ? _T_10366_24 : _T_16140; // @[Mux.scala 46:16:@14154.4]
  assign _T_16143 = 6'h18 == _T_11317_54; // @[Mux.scala 46:19:@14155.4]
  assign _T_16144 = _T_16143 ? _T_10366_23 : _T_16142; // @[Mux.scala 46:16:@14156.4]
  assign _T_16145 = 6'h17 == _T_11317_54; // @[Mux.scala 46:19:@14157.4]
  assign _T_16146 = _T_16145 ? _T_10366_22 : _T_16144; // @[Mux.scala 46:16:@14158.4]
  assign _T_16147 = 6'h16 == _T_11317_54; // @[Mux.scala 46:19:@14159.4]
  assign _T_16148 = _T_16147 ? _T_10366_21 : _T_16146; // @[Mux.scala 46:16:@14160.4]
  assign _T_16149 = 6'h15 == _T_11317_54; // @[Mux.scala 46:19:@14161.4]
  assign _T_16150 = _T_16149 ? _T_10366_20 : _T_16148; // @[Mux.scala 46:16:@14162.4]
  assign _T_16151 = 6'h14 == _T_11317_54; // @[Mux.scala 46:19:@14163.4]
  assign _T_16152 = _T_16151 ? _T_10366_19 : _T_16150; // @[Mux.scala 46:16:@14164.4]
  assign _T_16153 = 6'h13 == _T_11317_54; // @[Mux.scala 46:19:@14165.4]
  assign _T_16154 = _T_16153 ? _T_10366_18 : _T_16152; // @[Mux.scala 46:16:@14166.4]
  assign _T_16155 = 6'h12 == _T_11317_54; // @[Mux.scala 46:19:@14167.4]
  assign _T_16156 = _T_16155 ? _T_10366_17 : _T_16154; // @[Mux.scala 46:16:@14168.4]
  assign _T_16157 = 6'h11 == _T_11317_54; // @[Mux.scala 46:19:@14169.4]
  assign _T_16158 = _T_16157 ? _T_10366_16 : _T_16156; // @[Mux.scala 46:16:@14170.4]
  assign _T_16159 = 6'h10 == _T_11317_54; // @[Mux.scala 46:19:@14171.4]
  assign _T_16160 = _T_16159 ? _T_10366_15 : _T_16158; // @[Mux.scala 46:16:@14172.4]
  assign _T_16161 = 6'hf == _T_11317_54; // @[Mux.scala 46:19:@14173.4]
  assign _T_16162 = _T_16161 ? _T_10366_14 : _T_16160; // @[Mux.scala 46:16:@14174.4]
  assign _T_16163 = 6'he == _T_11317_54; // @[Mux.scala 46:19:@14175.4]
  assign _T_16164 = _T_16163 ? _T_10366_13 : _T_16162; // @[Mux.scala 46:16:@14176.4]
  assign _T_16165 = 6'hd == _T_11317_54; // @[Mux.scala 46:19:@14177.4]
  assign _T_16166 = _T_16165 ? _T_10366_12 : _T_16164; // @[Mux.scala 46:16:@14178.4]
  assign _T_16167 = 6'hc == _T_11317_54; // @[Mux.scala 46:19:@14179.4]
  assign _T_16168 = _T_16167 ? _T_10366_11 : _T_16166; // @[Mux.scala 46:16:@14180.4]
  assign _T_16169 = 6'hb == _T_11317_54; // @[Mux.scala 46:19:@14181.4]
  assign _T_16170 = _T_16169 ? _T_10366_10 : _T_16168; // @[Mux.scala 46:16:@14182.4]
  assign _T_16171 = 6'ha == _T_11317_54; // @[Mux.scala 46:19:@14183.4]
  assign _T_16172 = _T_16171 ? _T_10366_9 : _T_16170; // @[Mux.scala 46:16:@14184.4]
  assign _T_16173 = 6'h9 == _T_11317_54; // @[Mux.scala 46:19:@14185.4]
  assign _T_16174 = _T_16173 ? _T_10366_8 : _T_16172; // @[Mux.scala 46:16:@14186.4]
  assign _T_16175 = 6'h8 == _T_11317_54; // @[Mux.scala 46:19:@14187.4]
  assign _T_16176 = _T_16175 ? _T_10366_7 : _T_16174; // @[Mux.scala 46:16:@14188.4]
  assign _T_16177 = 6'h7 == _T_11317_54; // @[Mux.scala 46:19:@14189.4]
  assign _T_16178 = _T_16177 ? _T_10366_6 : _T_16176; // @[Mux.scala 46:16:@14190.4]
  assign _T_16179 = 6'h6 == _T_11317_54; // @[Mux.scala 46:19:@14191.4]
  assign _T_16180 = _T_16179 ? _T_10366_5 : _T_16178; // @[Mux.scala 46:16:@14192.4]
  assign _T_16181 = 6'h5 == _T_11317_54; // @[Mux.scala 46:19:@14193.4]
  assign _T_16182 = _T_16181 ? _T_10366_4 : _T_16180; // @[Mux.scala 46:16:@14194.4]
  assign _T_16183 = 6'h4 == _T_11317_54; // @[Mux.scala 46:19:@14195.4]
  assign _T_16184 = _T_16183 ? _T_10366_3 : _T_16182; // @[Mux.scala 46:16:@14196.4]
  assign _T_16185 = 6'h3 == _T_11317_54; // @[Mux.scala 46:19:@14197.4]
  assign _T_16186 = _T_16185 ? _T_10366_2 : _T_16184; // @[Mux.scala 46:16:@14198.4]
  assign _T_16187 = 6'h2 == _T_11317_54; // @[Mux.scala 46:19:@14199.4]
  assign _T_16188 = _T_16187 ? _T_10366_1 : _T_16186; // @[Mux.scala 46:16:@14200.4]
  assign _T_16189 = 6'h1 == _T_11317_54; // @[Mux.scala 46:19:@14201.4]
  assign _T_16190 = _T_16189 ? _T_10366_0 : _T_16188; // @[Mux.scala 46:16:@14202.4]
  assign _T_16248 = 6'h38 == _T_11317_55; // @[Mux.scala 46:19:@14204.4]
  assign _T_16249 = _T_16248 ? _T_10366_55 : 8'h0; // @[Mux.scala 46:16:@14205.4]
  assign _T_16250 = 6'h37 == _T_11317_55; // @[Mux.scala 46:19:@14206.4]
  assign _T_16251 = _T_16250 ? _T_10366_54 : _T_16249; // @[Mux.scala 46:16:@14207.4]
  assign _T_16252 = 6'h36 == _T_11317_55; // @[Mux.scala 46:19:@14208.4]
  assign _T_16253 = _T_16252 ? _T_10366_53 : _T_16251; // @[Mux.scala 46:16:@14209.4]
  assign _T_16254 = 6'h35 == _T_11317_55; // @[Mux.scala 46:19:@14210.4]
  assign _T_16255 = _T_16254 ? _T_10366_52 : _T_16253; // @[Mux.scala 46:16:@14211.4]
  assign _T_16256 = 6'h34 == _T_11317_55; // @[Mux.scala 46:19:@14212.4]
  assign _T_16257 = _T_16256 ? _T_10366_51 : _T_16255; // @[Mux.scala 46:16:@14213.4]
  assign _T_16258 = 6'h33 == _T_11317_55; // @[Mux.scala 46:19:@14214.4]
  assign _T_16259 = _T_16258 ? _T_10366_50 : _T_16257; // @[Mux.scala 46:16:@14215.4]
  assign _T_16260 = 6'h32 == _T_11317_55; // @[Mux.scala 46:19:@14216.4]
  assign _T_16261 = _T_16260 ? _T_10366_49 : _T_16259; // @[Mux.scala 46:16:@14217.4]
  assign _T_16262 = 6'h31 == _T_11317_55; // @[Mux.scala 46:19:@14218.4]
  assign _T_16263 = _T_16262 ? _T_10366_48 : _T_16261; // @[Mux.scala 46:16:@14219.4]
  assign _T_16264 = 6'h30 == _T_11317_55; // @[Mux.scala 46:19:@14220.4]
  assign _T_16265 = _T_16264 ? _T_10366_47 : _T_16263; // @[Mux.scala 46:16:@14221.4]
  assign _T_16266 = 6'h2f == _T_11317_55; // @[Mux.scala 46:19:@14222.4]
  assign _T_16267 = _T_16266 ? _T_10366_46 : _T_16265; // @[Mux.scala 46:16:@14223.4]
  assign _T_16268 = 6'h2e == _T_11317_55; // @[Mux.scala 46:19:@14224.4]
  assign _T_16269 = _T_16268 ? _T_10366_45 : _T_16267; // @[Mux.scala 46:16:@14225.4]
  assign _T_16270 = 6'h2d == _T_11317_55; // @[Mux.scala 46:19:@14226.4]
  assign _T_16271 = _T_16270 ? _T_10366_44 : _T_16269; // @[Mux.scala 46:16:@14227.4]
  assign _T_16272 = 6'h2c == _T_11317_55; // @[Mux.scala 46:19:@14228.4]
  assign _T_16273 = _T_16272 ? _T_10366_43 : _T_16271; // @[Mux.scala 46:16:@14229.4]
  assign _T_16274 = 6'h2b == _T_11317_55; // @[Mux.scala 46:19:@14230.4]
  assign _T_16275 = _T_16274 ? _T_10366_42 : _T_16273; // @[Mux.scala 46:16:@14231.4]
  assign _T_16276 = 6'h2a == _T_11317_55; // @[Mux.scala 46:19:@14232.4]
  assign _T_16277 = _T_16276 ? _T_10366_41 : _T_16275; // @[Mux.scala 46:16:@14233.4]
  assign _T_16278 = 6'h29 == _T_11317_55; // @[Mux.scala 46:19:@14234.4]
  assign _T_16279 = _T_16278 ? _T_10366_40 : _T_16277; // @[Mux.scala 46:16:@14235.4]
  assign _T_16280 = 6'h28 == _T_11317_55; // @[Mux.scala 46:19:@14236.4]
  assign _T_16281 = _T_16280 ? _T_10366_39 : _T_16279; // @[Mux.scala 46:16:@14237.4]
  assign _T_16282 = 6'h27 == _T_11317_55; // @[Mux.scala 46:19:@14238.4]
  assign _T_16283 = _T_16282 ? _T_10366_38 : _T_16281; // @[Mux.scala 46:16:@14239.4]
  assign _T_16284 = 6'h26 == _T_11317_55; // @[Mux.scala 46:19:@14240.4]
  assign _T_16285 = _T_16284 ? _T_10366_37 : _T_16283; // @[Mux.scala 46:16:@14241.4]
  assign _T_16286 = 6'h25 == _T_11317_55; // @[Mux.scala 46:19:@14242.4]
  assign _T_16287 = _T_16286 ? _T_10366_36 : _T_16285; // @[Mux.scala 46:16:@14243.4]
  assign _T_16288 = 6'h24 == _T_11317_55; // @[Mux.scala 46:19:@14244.4]
  assign _T_16289 = _T_16288 ? _T_10366_35 : _T_16287; // @[Mux.scala 46:16:@14245.4]
  assign _T_16290 = 6'h23 == _T_11317_55; // @[Mux.scala 46:19:@14246.4]
  assign _T_16291 = _T_16290 ? _T_10366_34 : _T_16289; // @[Mux.scala 46:16:@14247.4]
  assign _T_16292 = 6'h22 == _T_11317_55; // @[Mux.scala 46:19:@14248.4]
  assign _T_16293 = _T_16292 ? _T_10366_33 : _T_16291; // @[Mux.scala 46:16:@14249.4]
  assign _T_16294 = 6'h21 == _T_11317_55; // @[Mux.scala 46:19:@14250.4]
  assign _T_16295 = _T_16294 ? _T_10366_32 : _T_16293; // @[Mux.scala 46:16:@14251.4]
  assign _T_16296 = 6'h20 == _T_11317_55; // @[Mux.scala 46:19:@14252.4]
  assign _T_16297 = _T_16296 ? _T_10366_31 : _T_16295; // @[Mux.scala 46:16:@14253.4]
  assign _T_16298 = 6'h1f == _T_11317_55; // @[Mux.scala 46:19:@14254.4]
  assign _T_16299 = _T_16298 ? _T_10366_30 : _T_16297; // @[Mux.scala 46:16:@14255.4]
  assign _T_16300 = 6'h1e == _T_11317_55; // @[Mux.scala 46:19:@14256.4]
  assign _T_16301 = _T_16300 ? _T_10366_29 : _T_16299; // @[Mux.scala 46:16:@14257.4]
  assign _T_16302 = 6'h1d == _T_11317_55; // @[Mux.scala 46:19:@14258.4]
  assign _T_16303 = _T_16302 ? _T_10366_28 : _T_16301; // @[Mux.scala 46:16:@14259.4]
  assign _T_16304 = 6'h1c == _T_11317_55; // @[Mux.scala 46:19:@14260.4]
  assign _T_16305 = _T_16304 ? _T_10366_27 : _T_16303; // @[Mux.scala 46:16:@14261.4]
  assign _T_16306 = 6'h1b == _T_11317_55; // @[Mux.scala 46:19:@14262.4]
  assign _T_16307 = _T_16306 ? _T_10366_26 : _T_16305; // @[Mux.scala 46:16:@14263.4]
  assign _T_16308 = 6'h1a == _T_11317_55; // @[Mux.scala 46:19:@14264.4]
  assign _T_16309 = _T_16308 ? _T_10366_25 : _T_16307; // @[Mux.scala 46:16:@14265.4]
  assign _T_16310 = 6'h19 == _T_11317_55; // @[Mux.scala 46:19:@14266.4]
  assign _T_16311 = _T_16310 ? _T_10366_24 : _T_16309; // @[Mux.scala 46:16:@14267.4]
  assign _T_16312 = 6'h18 == _T_11317_55; // @[Mux.scala 46:19:@14268.4]
  assign _T_16313 = _T_16312 ? _T_10366_23 : _T_16311; // @[Mux.scala 46:16:@14269.4]
  assign _T_16314 = 6'h17 == _T_11317_55; // @[Mux.scala 46:19:@14270.4]
  assign _T_16315 = _T_16314 ? _T_10366_22 : _T_16313; // @[Mux.scala 46:16:@14271.4]
  assign _T_16316 = 6'h16 == _T_11317_55; // @[Mux.scala 46:19:@14272.4]
  assign _T_16317 = _T_16316 ? _T_10366_21 : _T_16315; // @[Mux.scala 46:16:@14273.4]
  assign _T_16318 = 6'h15 == _T_11317_55; // @[Mux.scala 46:19:@14274.4]
  assign _T_16319 = _T_16318 ? _T_10366_20 : _T_16317; // @[Mux.scala 46:16:@14275.4]
  assign _T_16320 = 6'h14 == _T_11317_55; // @[Mux.scala 46:19:@14276.4]
  assign _T_16321 = _T_16320 ? _T_10366_19 : _T_16319; // @[Mux.scala 46:16:@14277.4]
  assign _T_16322 = 6'h13 == _T_11317_55; // @[Mux.scala 46:19:@14278.4]
  assign _T_16323 = _T_16322 ? _T_10366_18 : _T_16321; // @[Mux.scala 46:16:@14279.4]
  assign _T_16324 = 6'h12 == _T_11317_55; // @[Mux.scala 46:19:@14280.4]
  assign _T_16325 = _T_16324 ? _T_10366_17 : _T_16323; // @[Mux.scala 46:16:@14281.4]
  assign _T_16326 = 6'h11 == _T_11317_55; // @[Mux.scala 46:19:@14282.4]
  assign _T_16327 = _T_16326 ? _T_10366_16 : _T_16325; // @[Mux.scala 46:16:@14283.4]
  assign _T_16328 = 6'h10 == _T_11317_55; // @[Mux.scala 46:19:@14284.4]
  assign _T_16329 = _T_16328 ? _T_10366_15 : _T_16327; // @[Mux.scala 46:16:@14285.4]
  assign _T_16330 = 6'hf == _T_11317_55; // @[Mux.scala 46:19:@14286.4]
  assign _T_16331 = _T_16330 ? _T_10366_14 : _T_16329; // @[Mux.scala 46:16:@14287.4]
  assign _T_16332 = 6'he == _T_11317_55; // @[Mux.scala 46:19:@14288.4]
  assign _T_16333 = _T_16332 ? _T_10366_13 : _T_16331; // @[Mux.scala 46:16:@14289.4]
  assign _T_16334 = 6'hd == _T_11317_55; // @[Mux.scala 46:19:@14290.4]
  assign _T_16335 = _T_16334 ? _T_10366_12 : _T_16333; // @[Mux.scala 46:16:@14291.4]
  assign _T_16336 = 6'hc == _T_11317_55; // @[Mux.scala 46:19:@14292.4]
  assign _T_16337 = _T_16336 ? _T_10366_11 : _T_16335; // @[Mux.scala 46:16:@14293.4]
  assign _T_16338 = 6'hb == _T_11317_55; // @[Mux.scala 46:19:@14294.4]
  assign _T_16339 = _T_16338 ? _T_10366_10 : _T_16337; // @[Mux.scala 46:16:@14295.4]
  assign _T_16340 = 6'ha == _T_11317_55; // @[Mux.scala 46:19:@14296.4]
  assign _T_16341 = _T_16340 ? _T_10366_9 : _T_16339; // @[Mux.scala 46:16:@14297.4]
  assign _T_16342 = 6'h9 == _T_11317_55; // @[Mux.scala 46:19:@14298.4]
  assign _T_16343 = _T_16342 ? _T_10366_8 : _T_16341; // @[Mux.scala 46:16:@14299.4]
  assign _T_16344 = 6'h8 == _T_11317_55; // @[Mux.scala 46:19:@14300.4]
  assign _T_16345 = _T_16344 ? _T_10366_7 : _T_16343; // @[Mux.scala 46:16:@14301.4]
  assign _T_16346 = 6'h7 == _T_11317_55; // @[Mux.scala 46:19:@14302.4]
  assign _T_16347 = _T_16346 ? _T_10366_6 : _T_16345; // @[Mux.scala 46:16:@14303.4]
  assign _T_16348 = 6'h6 == _T_11317_55; // @[Mux.scala 46:19:@14304.4]
  assign _T_16349 = _T_16348 ? _T_10366_5 : _T_16347; // @[Mux.scala 46:16:@14305.4]
  assign _T_16350 = 6'h5 == _T_11317_55; // @[Mux.scala 46:19:@14306.4]
  assign _T_16351 = _T_16350 ? _T_10366_4 : _T_16349; // @[Mux.scala 46:16:@14307.4]
  assign _T_16352 = 6'h4 == _T_11317_55; // @[Mux.scala 46:19:@14308.4]
  assign _T_16353 = _T_16352 ? _T_10366_3 : _T_16351; // @[Mux.scala 46:16:@14309.4]
  assign _T_16354 = 6'h3 == _T_11317_55; // @[Mux.scala 46:19:@14310.4]
  assign _T_16355 = _T_16354 ? _T_10366_2 : _T_16353; // @[Mux.scala 46:16:@14311.4]
  assign _T_16356 = 6'h2 == _T_11317_55; // @[Mux.scala 46:19:@14312.4]
  assign _T_16357 = _T_16356 ? _T_10366_1 : _T_16355; // @[Mux.scala 46:16:@14313.4]
  assign _T_16358 = 6'h1 == _T_11317_55; // @[Mux.scala 46:19:@14314.4]
  assign _T_16359 = _T_16358 ? _T_10366_0 : _T_16357; // @[Mux.scala 46:16:@14315.4]
  assign _T_16418 = 6'h39 == _T_11317_56; // @[Mux.scala 46:19:@14317.4]
  assign _T_16419 = _T_16418 ? _T_10366_56 : 8'h0; // @[Mux.scala 46:16:@14318.4]
  assign _T_16420 = 6'h38 == _T_11317_56; // @[Mux.scala 46:19:@14319.4]
  assign _T_16421 = _T_16420 ? _T_10366_55 : _T_16419; // @[Mux.scala 46:16:@14320.4]
  assign _T_16422 = 6'h37 == _T_11317_56; // @[Mux.scala 46:19:@14321.4]
  assign _T_16423 = _T_16422 ? _T_10366_54 : _T_16421; // @[Mux.scala 46:16:@14322.4]
  assign _T_16424 = 6'h36 == _T_11317_56; // @[Mux.scala 46:19:@14323.4]
  assign _T_16425 = _T_16424 ? _T_10366_53 : _T_16423; // @[Mux.scala 46:16:@14324.4]
  assign _T_16426 = 6'h35 == _T_11317_56; // @[Mux.scala 46:19:@14325.4]
  assign _T_16427 = _T_16426 ? _T_10366_52 : _T_16425; // @[Mux.scala 46:16:@14326.4]
  assign _T_16428 = 6'h34 == _T_11317_56; // @[Mux.scala 46:19:@14327.4]
  assign _T_16429 = _T_16428 ? _T_10366_51 : _T_16427; // @[Mux.scala 46:16:@14328.4]
  assign _T_16430 = 6'h33 == _T_11317_56; // @[Mux.scala 46:19:@14329.4]
  assign _T_16431 = _T_16430 ? _T_10366_50 : _T_16429; // @[Mux.scala 46:16:@14330.4]
  assign _T_16432 = 6'h32 == _T_11317_56; // @[Mux.scala 46:19:@14331.4]
  assign _T_16433 = _T_16432 ? _T_10366_49 : _T_16431; // @[Mux.scala 46:16:@14332.4]
  assign _T_16434 = 6'h31 == _T_11317_56; // @[Mux.scala 46:19:@14333.4]
  assign _T_16435 = _T_16434 ? _T_10366_48 : _T_16433; // @[Mux.scala 46:16:@14334.4]
  assign _T_16436 = 6'h30 == _T_11317_56; // @[Mux.scala 46:19:@14335.4]
  assign _T_16437 = _T_16436 ? _T_10366_47 : _T_16435; // @[Mux.scala 46:16:@14336.4]
  assign _T_16438 = 6'h2f == _T_11317_56; // @[Mux.scala 46:19:@14337.4]
  assign _T_16439 = _T_16438 ? _T_10366_46 : _T_16437; // @[Mux.scala 46:16:@14338.4]
  assign _T_16440 = 6'h2e == _T_11317_56; // @[Mux.scala 46:19:@14339.4]
  assign _T_16441 = _T_16440 ? _T_10366_45 : _T_16439; // @[Mux.scala 46:16:@14340.4]
  assign _T_16442 = 6'h2d == _T_11317_56; // @[Mux.scala 46:19:@14341.4]
  assign _T_16443 = _T_16442 ? _T_10366_44 : _T_16441; // @[Mux.scala 46:16:@14342.4]
  assign _T_16444 = 6'h2c == _T_11317_56; // @[Mux.scala 46:19:@14343.4]
  assign _T_16445 = _T_16444 ? _T_10366_43 : _T_16443; // @[Mux.scala 46:16:@14344.4]
  assign _T_16446 = 6'h2b == _T_11317_56; // @[Mux.scala 46:19:@14345.4]
  assign _T_16447 = _T_16446 ? _T_10366_42 : _T_16445; // @[Mux.scala 46:16:@14346.4]
  assign _T_16448 = 6'h2a == _T_11317_56; // @[Mux.scala 46:19:@14347.4]
  assign _T_16449 = _T_16448 ? _T_10366_41 : _T_16447; // @[Mux.scala 46:16:@14348.4]
  assign _T_16450 = 6'h29 == _T_11317_56; // @[Mux.scala 46:19:@14349.4]
  assign _T_16451 = _T_16450 ? _T_10366_40 : _T_16449; // @[Mux.scala 46:16:@14350.4]
  assign _T_16452 = 6'h28 == _T_11317_56; // @[Mux.scala 46:19:@14351.4]
  assign _T_16453 = _T_16452 ? _T_10366_39 : _T_16451; // @[Mux.scala 46:16:@14352.4]
  assign _T_16454 = 6'h27 == _T_11317_56; // @[Mux.scala 46:19:@14353.4]
  assign _T_16455 = _T_16454 ? _T_10366_38 : _T_16453; // @[Mux.scala 46:16:@14354.4]
  assign _T_16456 = 6'h26 == _T_11317_56; // @[Mux.scala 46:19:@14355.4]
  assign _T_16457 = _T_16456 ? _T_10366_37 : _T_16455; // @[Mux.scala 46:16:@14356.4]
  assign _T_16458 = 6'h25 == _T_11317_56; // @[Mux.scala 46:19:@14357.4]
  assign _T_16459 = _T_16458 ? _T_10366_36 : _T_16457; // @[Mux.scala 46:16:@14358.4]
  assign _T_16460 = 6'h24 == _T_11317_56; // @[Mux.scala 46:19:@14359.4]
  assign _T_16461 = _T_16460 ? _T_10366_35 : _T_16459; // @[Mux.scala 46:16:@14360.4]
  assign _T_16462 = 6'h23 == _T_11317_56; // @[Mux.scala 46:19:@14361.4]
  assign _T_16463 = _T_16462 ? _T_10366_34 : _T_16461; // @[Mux.scala 46:16:@14362.4]
  assign _T_16464 = 6'h22 == _T_11317_56; // @[Mux.scala 46:19:@14363.4]
  assign _T_16465 = _T_16464 ? _T_10366_33 : _T_16463; // @[Mux.scala 46:16:@14364.4]
  assign _T_16466 = 6'h21 == _T_11317_56; // @[Mux.scala 46:19:@14365.4]
  assign _T_16467 = _T_16466 ? _T_10366_32 : _T_16465; // @[Mux.scala 46:16:@14366.4]
  assign _T_16468 = 6'h20 == _T_11317_56; // @[Mux.scala 46:19:@14367.4]
  assign _T_16469 = _T_16468 ? _T_10366_31 : _T_16467; // @[Mux.scala 46:16:@14368.4]
  assign _T_16470 = 6'h1f == _T_11317_56; // @[Mux.scala 46:19:@14369.4]
  assign _T_16471 = _T_16470 ? _T_10366_30 : _T_16469; // @[Mux.scala 46:16:@14370.4]
  assign _T_16472 = 6'h1e == _T_11317_56; // @[Mux.scala 46:19:@14371.4]
  assign _T_16473 = _T_16472 ? _T_10366_29 : _T_16471; // @[Mux.scala 46:16:@14372.4]
  assign _T_16474 = 6'h1d == _T_11317_56; // @[Mux.scala 46:19:@14373.4]
  assign _T_16475 = _T_16474 ? _T_10366_28 : _T_16473; // @[Mux.scala 46:16:@14374.4]
  assign _T_16476 = 6'h1c == _T_11317_56; // @[Mux.scala 46:19:@14375.4]
  assign _T_16477 = _T_16476 ? _T_10366_27 : _T_16475; // @[Mux.scala 46:16:@14376.4]
  assign _T_16478 = 6'h1b == _T_11317_56; // @[Mux.scala 46:19:@14377.4]
  assign _T_16479 = _T_16478 ? _T_10366_26 : _T_16477; // @[Mux.scala 46:16:@14378.4]
  assign _T_16480 = 6'h1a == _T_11317_56; // @[Mux.scala 46:19:@14379.4]
  assign _T_16481 = _T_16480 ? _T_10366_25 : _T_16479; // @[Mux.scala 46:16:@14380.4]
  assign _T_16482 = 6'h19 == _T_11317_56; // @[Mux.scala 46:19:@14381.4]
  assign _T_16483 = _T_16482 ? _T_10366_24 : _T_16481; // @[Mux.scala 46:16:@14382.4]
  assign _T_16484 = 6'h18 == _T_11317_56; // @[Mux.scala 46:19:@14383.4]
  assign _T_16485 = _T_16484 ? _T_10366_23 : _T_16483; // @[Mux.scala 46:16:@14384.4]
  assign _T_16486 = 6'h17 == _T_11317_56; // @[Mux.scala 46:19:@14385.4]
  assign _T_16487 = _T_16486 ? _T_10366_22 : _T_16485; // @[Mux.scala 46:16:@14386.4]
  assign _T_16488 = 6'h16 == _T_11317_56; // @[Mux.scala 46:19:@14387.4]
  assign _T_16489 = _T_16488 ? _T_10366_21 : _T_16487; // @[Mux.scala 46:16:@14388.4]
  assign _T_16490 = 6'h15 == _T_11317_56; // @[Mux.scala 46:19:@14389.4]
  assign _T_16491 = _T_16490 ? _T_10366_20 : _T_16489; // @[Mux.scala 46:16:@14390.4]
  assign _T_16492 = 6'h14 == _T_11317_56; // @[Mux.scala 46:19:@14391.4]
  assign _T_16493 = _T_16492 ? _T_10366_19 : _T_16491; // @[Mux.scala 46:16:@14392.4]
  assign _T_16494 = 6'h13 == _T_11317_56; // @[Mux.scala 46:19:@14393.4]
  assign _T_16495 = _T_16494 ? _T_10366_18 : _T_16493; // @[Mux.scala 46:16:@14394.4]
  assign _T_16496 = 6'h12 == _T_11317_56; // @[Mux.scala 46:19:@14395.4]
  assign _T_16497 = _T_16496 ? _T_10366_17 : _T_16495; // @[Mux.scala 46:16:@14396.4]
  assign _T_16498 = 6'h11 == _T_11317_56; // @[Mux.scala 46:19:@14397.4]
  assign _T_16499 = _T_16498 ? _T_10366_16 : _T_16497; // @[Mux.scala 46:16:@14398.4]
  assign _T_16500 = 6'h10 == _T_11317_56; // @[Mux.scala 46:19:@14399.4]
  assign _T_16501 = _T_16500 ? _T_10366_15 : _T_16499; // @[Mux.scala 46:16:@14400.4]
  assign _T_16502 = 6'hf == _T_11317_56; // @[Mux.scala 46:19:@14401.4]
  assign _T_16503 = _T_16502 ? _T_10366_14 : _T_16501; // @[Mux.scala 46:16:@14402.4]
  assign _T_16504 = 6'he == _T_11317_56; // @[Mux.scala 46:19:@14403.4]
  assign _T_16505 = _T_16504 ? _T_10366_13 : _T_16503; // @[Mux.scala 46:16:@14404.4]
  assign _T_16506 = 6'hd == _T_11317_56; // @[Mux.scala 46:19:@14405.4]
  assign _T_16507 = _T_16506 ? _T_10366_12 : _T_16505; // @[Mux.scala 46:16:@14406.4]
  assign _T_16508 = 6'hc == _T_11317_56; // @[Mux.scala 46:19:@14407.4]
  assign _T_16509 = _T_16508 ? _T_10366_11 : _T_16507; // @[Mux.scala 46:16:@14408.4]
  assign _T_16510 = 6'hb == _T_11317_56; // @[Mux.scala 46:19:@14409.4]
  assign _T_16511 = _T_16510 ? _T_10366_10 : _T_16509; // @[Mux.scala 46:16:@14410.4]
  assign _T_16512 = 6'ha == _T_11317_56; // @[Mux.scala 46:19:@14411.4]
  assign _T_16513 = _T_16512 ? _T_10366_9 : _T_16511; // @[Mux.scala 46:16:@14412.4]
  assign _T_16514 = 6'h9 == _T_11317_56; // @[Mux.scala 46:19:@14413.4]
  assign _T_16515 = _T_16514 ? _T_10366_8 : _T_16513; // @[Mux.scala 46:16:@14414.4]
  assign _T_16516 = 6'h8 == _T_11317_56; // @[Mux.scala 46:19:@14415.4]
  assign _T_16517 = _T_16516 ? _T_10366_7 : _T_16515; // @[Mux.scala 46:16:@14416.4]
  assign _T_16518 = 6'h7 == _T_11317_56; // @[Mux.scala 46:19:@14417.4]
  assign _T_16519 = _T_16518 ? _T_10366_6 : _T_16517; // @[Mux.scala 46:16:@14418.4]
  assign _T_16520 = 6'h6 == _T_11317_56; // @[Mux.scala 46:19:@14419.4]
  assign _T_16521 = _T_16520 ? _T_10366_5 : _T_16519; // @[Mux.scala 46:16:@14420.4]
  assign _T_16522 = 6'h5 == _T_11317_56; // @[Mux.scala 46:19:@14421.4]
  assign _T_16523 = _T_16522 ? _T_10366_4 : _T_16521; // @[Mux.scala 46:16:@14422.4]
  assign _T_16524 = 6'h4 == _T_11317_56; // @[Mux.scala 46:19:@14423.4]
  assign _T_16525 = _T_16524 ? _T_10366_3 : _T_16523; // @[Mux.scala 46:16:@14424.4]
  assign _T_16526 = 6'h3 == _T_11317_56; // @[Mux.scala 46:19:@14425.4]
  assign _T_16527 = _T_16526 ? _T_10366_2 : _T_16525; // @[Mux.scala 46:16:@14426.4]
  assign _T_16528 = 6'h2 == _T_11317_56; // @[Mux.scala 46:19:@14427.4]
  assign _T_16529 = _T_16528 ? _T_10366_1 : _T_16527; // @[Mux.scala 46:16:@14428.4]
  assign _T_16530 = 6'h1 == _T_11317_56; // @[Mux.scala 46:19:@14429.4]
  assign _T_16531 = _T_16530 ? _T_10366_0 : _T_16529; // @[Mux.scala 46:16:@14430.4]
  assign _T_16591 = 6'h3a == _T_11317_57; // @[Mux.scala 46:19:@14432.4]
  assign _T_16592 = _T_16591 ? _T_10366_57 : 8'h0; // @[Mux.scala 46:16:@14433.4]
  assign _T_16593 = 6'h39 == _T_11317_57; // @[Mux.scala 46:19:@14434.4]
  assign _T_16594 = _T_16593 ? _T_10366_56 : _T_16592; // @[Mux.scala 46:16:@14435.4]
  assign _T_16595 = 6'h38 == _T_11317_57; // @[Mux.scala 46:19:@14436.4]
  assign _T_16596 = _T_16595 ? _T_10366_55 : _T_16594; // @[Mux.scala 46:16:@14437.4]
  assign _T_16597 = 6'h37 == _T_11317_57; // @[Mux.scala 46:19:@14438.4]
  assign _T_16598 = _T_16597 ? _T_10366_54 : _T_16596; // @[Mux.scala 46:16:@14439.4]
  assign _T_16599 = 6'h36 == _T_11317_57; // @[Mux.scala 46:19:@14440.4]
  assign _T_16600 = _T_16599 ? _T_10366_53 : _T_16598; // @[Mux.scala 46:16:@14441.4]
  assign _T_16601 = 6'h35 == _T_11317_57; // @[Mux.scala 46:19:@14442.4]
  assign _T_16602 = _T_16601 ? _T_10366_52 : _T_16600; // @[Mux.scala 46:16:@14443.4]
  assign _T_16603 = 6'h34 == _T_11317_57; // @[Mux.scala 46:19:@14444.4]
  assign _T_16604 = _T_16603 ? _T_10366_51 : _T_16602; // @[Mux.scala 46:16:@14445.4]
  assign _T_16605 = 6'h33 == _T_11317_57; // @[Mux.scala 46:19:@14446.4]
  assign _T_16606 = _T_16605 ? _T_10366_50 : _T_16604; // @[Mux.scala 46:16:@14447.4]
  assign _T_16607 = 6'h32 == _T_11317_57; // @[Mux.scala 46:19:@14448.4]
  assign _T_16608 = _T_16607 ? _T_10366_49 : _T_16606; // @[Mux.scala 46:16:@14449.4]
  assign _T_16609 = 6'h31 == _T_11317_57; // @[Mux.scala 46:19:@14450.4]
  assign _T_16610 = _T_16609 ? _T_10366_48 : _T_16608; // @[Mux.scala 46:16:@14451.4]
  assign _T_16611 = 6'h30 == _T_11317_57; // @[Mux.scala 46:19:@14452.4]
  assign _T_16612 = _T_16611 ? _T_10366_47 : _T_16610; // @[Mux.scala 46:16:@14453.4]
  assign _T_16613 = 6'h2f == _T_11317_57; // @[Mux.scala 46:19:@14454.4]
  assign _T_16614 = _T_16613 ? _T_10366_46 : _T_16612; // @[Mux.scala 46:16:@14455.4]
  assign _T_16615 = 6'h2e == _T_11317_57; // @[Mux.scala 46:19:@14456.4]
  assign _T_16616 = _T_16615 ? _T_10366_45 : _T_16614; // @[Mux.scala 46:16:@14457.4]
  assign _T_16617 = 6'h2d == _T_11317_57; // @[Mux.scala 46:19:@14458.4]
  assign _T_16618 = _T_16617 ? _T_10366_44 : _T_16616; // @[Mux.scala 46:16:@14459.4]
  assign _T_16619 = 6'h2c == _T_11317_57; // @[Mux.scala 46:19:@14460.4]
  assign _T_16620 = _T_16619 ? _T_10366_43 : _T_16618; // @[Mux.scala 46:16:@14461.4]
  assign _T_16621 = 6'h2b == _T_11317_57; // @[Mux.scala 46:19:@14462.4]
  assign _T_16622 = _T_16621 ? _T_10366_42 : _T_16620; // @[Mux.scala 46:16:@14463.4]
  assign _T_16623 = 6'h2a == _T_11317_57; // @[Mux.scala 46:19:@14464.4]
  assign _T_16624 = _T_16623 ? _T_10366_41 : _T_16622; // @[Mux.scala 46:16:@14465.4]
  assign _T_16625 = 6'h29 == _T_11317_57; // @[Mux.scala 46:19:@14466.4]
  assign _T_16626 = _T_16625 ? _T_10366_40 : _T_16624; // @[Mux.scala 46:16:@14467.4]
  assign _T_16627 = 6'h28 == _T_11317_57; // @[Mux.scala 46:19:@14468.4]
  assign _T_16628 = _T_16627 ? _T_10366_39 : _T_16626; // @[Mux.scala 46:16:@14469.4]
  assign _T_16629 = 6'h27 == _T_11317_57; // @[Mux.scala 46:19:@14470.4]
  assign _T_16630 = _T_16629 ? _T_10366_38 : _T_16628; // @[Mux.scala 46:16:@14471.4]
  assign _T_16631 = 6'h26 == _T_11317_57; // @[Mux.scala 46:19:@14472.4]
  assign _T_16632 = _T_16631 ? _T_10366_37 : _T_16630; // @[Mux.scala 46:16:@14473.4]
  assign _T_16633 = 6'h25 == _T_11317_57; // @[Mux.scala 46:19:@14474.4]
  assign _T_16634 = _T_16633 ? _T_10366_36 : _T_16632; // @[Mux.scala 46:16:@14475.4]
  assign _T_16635 = 6'h24 == _T_11317_57; // @[Mux.scala 46:19:@14476.4]
  assign _T_16636 = _T_16635 ? _T_10366_35 : _T_16634; // @[Mux.scala 46:16:@14477.4]
  assign _T_16637 = 6'h23 == _T_11317_57; // @[Mux.scala 46:19:@14478.4]
  assign _T_16638 = _T_16637 ? _T_10366_34 : _T_16636; // @[Mux.scala 46:16:@14479.4]
  assign _T_16639 = 6'h22 == _T_11317_57; // @[Mux.scala 46:19:@14480.4]
  assign _T_16640 = _T_16639 ? _T_10366_33 : _T_16638; // @[Mux.scala 46:16:@14481.4]
  assign _T_16641 = 6'h21 == _T_11317_57; // @[Mux.scala 46:19:@14482.4]
  assign _T_16642 = _T_16641 ? _T_10366_32 : _T_16640; // @[Mux.scala 46:16:@14483.4]
  assign _T_16643 = 6'h20 == _T_11317_57; // @[Mux.scala 46:19:@14484.4]
  assign _T_16644 = _T_16643 ? _T_10366_31 : _T_16642; // @[Mux.scala 46:16:@14485.4]
  assign _T_16645 = 6'h1f == _T_11317_57; // @[Mux.scala 46:19:@14486.4]
  assign _T_16646 = _T_16645 ? _T_10366_30 : _T_16644; // @[Mux.scala 46:16:@14487.4]
  assign _T_16647 = 6'h1e == _T_11317_57; // @[Mux.scala 46:19:@14488.4]
  assign _T_16648 = _T_16647 ? _T_10366_29 : _T_16646; // @[Mux.scala 46:16:@14489.4]
  assign _T_16649 = 6'h1d == _T_11317_57; // @[Mux.scala 46:19:@14490.4]
  assign _T_16650 = _T_16649 ? _T_10366_28 : _T_16648; // @[Mux.scala 46:16:@14491.4]
  assign _T_16651 = 6'h1c == _T_11317_57; // @[Mux.scala 46:19:@14492.4]
  assign _T_16652 = _T_16651 ? _T_10366_27 : _T_16650; // @[Mux.scala 46:16:@14493.4]
  assign _T_16653 = 6'h1b == _T_11317_57; // @[Mux.scala 46:19:@14494.4]
  assign _T_16654 = _T_16653 ? _T_10366_26 : _T_16652; // @[Mux.scala 46:16:@14495.4]
  assign _T_16655 = 6'h1a == _T_11317_57; // @[Mux.scala 46:19:@14496.4]
  assign _T_16656 = _T_16655 ? _T_10366_25 : _T_16654; // @[Mux.scala 46:16:@14497.4]
  assign _T_16657 = 6'h19 == _T_11317_57; // @[Mux.scala 46:19:@14498.4]
  assign _T_16658 = _T_16657 ? _T_10366_24 : _T_16656; // @[Mux.scala 46:16:@14499.4]
  assign _T_16659 = 6'h18 == _T_11317_57; // @[Mux.scala 46:19:@14500.4]
  assign _T_16660 = _T_16659 ? _T_10366_23 : _T_16658; // @[Mux.scala 46:16:@14501.4]
  assign _T_16661 = 6'h17 == _T_11317_57; // @[Mux.scala 46:19:@14502.4]
  assign _T_16662 = _T_16661 ? _T_10366_22 : _T_16660; // @[Mux.scala 46:16:@14503.4]
  assign _T_16663 = 6'h16 == _T_11317_57; // @[Mux.scala 46:19:@14504.4]
  assign _T_16664 = _T_16663 ? _T_10366_21 : _T_16662; // @[Mux.scala 46:16:@14505.4]
  assign _T_16665 = 6'h15 == _T_11317_57; // @[Mux.scala 46:19:@14506.4]
  assign _T_16666 = _T_16665 ? _T_10366_20 : _T_16664; // @[Mux.scala 46:16:@14507.4]
  assign _T_16667 = 6'h14 == _T_11317_57; // @[Mux.scala 46:19:@14508.4]
  assign _T_16668 = _T_16667 ? _T_10366_19 : _T_16666; // @[Mux.scala 46:16:@14509.4]
  assign _T_16669 = 6'h13 == _T_11317_57; // @[Mux.scala 46:19:@14510.4]
  assign _T_16670 = _T_16669 ? _T_10366_18 : _T_16668; // @[Mux.scala 46:16:@14511.4]
  assign _T_16671 = 6'h12 == _T_11317_57; // @[Mux.scala 46:19:@14512.4]
  assign _T_16672 = _T_16671 ? _T_10366_17 : _T_16670; // @[Mux.scala 46:16:@14513.4]
  assign _T_16673 = 6'h11 == _T_11317_57; // @[Mux.scala 46:19:@14514.4]
  assign _T_16674 = _T_16673 ? _T_10366_16 : _T_16672; // @[Mux.scala 46:16:@14515.4]
  assign _T_16675 = 6'h10 == _T_11317_57; // @[Mux.scala 46:19:@14516.4]
  assign _T_16676 = _T_16675 ? _T_10366_15 : _T_16674; // @[Mux.scala 46:16:@14517.4]
  assign _T_16677 = 6'hf == _T_11317_57; // @[Mux.scala 46:19:@14518.4]
  assign _T_16678 = _T_16677 ? _T_10366_14 : _T_16676; // @[Mux.scala 46:16:@14519.4]
  assign _T_16679 = 6'he == _T_11317_57; // @[Mux.scala 46:19:@14520.4]
  assign _T_16680 = _T_16679 ? _T_10366_13 : _T_16678; // @[Mux.scala 46:16:@14521.4]
  assign _T_16681 = 6'hd == _T_11317_57; // @[Mux.scala 46:19:@14522.4]
  assign _T_16682 = _T_16681 ? _T_10366_12 : _T_16680; // @[Mux.scala 46:16:@14523.4]
  assign _T_16683 = 6'hc == _T_11317_57; // @[Mux.scala 46:19:@14524.4]
  assign _T_16684 = _T_16683 ? _T_10366_11 : _T_16682; // @[Mux.scala 46:16:@14525.4]
  assign _T_16685 = 6'hb == _T_11317_57; // @[Mux.scala 46:19:@14526.4]
  assign _T_16686 = _T_16685 ? _T_10366_10 : _T_16684; // @[Mux.scala 46:16:@14527.4]
  assign _T_16687 = 6'ha == _T_11317_57; // @[Mux.scala 46:19:@14528.4]
  assign _T_16688 = _T_16687 ? _T_10366_9 : _T_16686; // @[Mux.scala 46:16:@14529.4]
  assign _T_16689 = 6'h9 == _T_11317_57; // @[Mux.scala 46:19:@14530.4]
  assign _T_16690 = _T_16689 ? _T_10366_8 : _T_16688; // @[Mux.scala 46:16:@14531.4]
  assign _T_16691 = 6'h8 == _T_11317_57; // @[Mux.scala 46:19:@14532.4]
  assign _T_16692 = _T_16691 ? _T_10366_7 : _T_16690; // @[Mux.scala 46:16:@14533.4]
  assign _T_16693 = 6'h7 == _T_11317_57; // @[Mux.scala 46:19:@14534.4]
  assign _T_16694 = _T_16693 ? _T_10366_6 : _T_16692; // @[Mux.scala 46:16:@14535.4]
  assign _T_16695 = 6'h6 == _T_11317_57; // @[Mux.scala 46:19:@14536.4]
  assign _T_16696 = _T_16695 ? _T_10366_5 : _T_16694; // @[Mux.scala 46:16:@14537.4]
  assign _T_16697 = 6'h5 == _T_11317_57; // @[Mux.scala 46:19:@14538.4]
  assign _T_16698 = _T_16697 ? _T_10366_4 : _T_16696; // @[Mux.scala 46:16:@14539.4]
  assign _T_16699 = 6'h4 == _T_11317_57; // @[Mux.scala 46:19:@14540.4]
  assign _T_16700 = _T_16699 ? _T_10366_3 : _T_16698; // @[Mux.scala 46:16:@14541.4]
  assign _T_16701 = 6'h3 == _T_11317_57; // @[Mux.scala 46:19:@14542.4]
  assign _T_16702 = _T_16701 ? _T_10366_2 : _T_16700; // @[Mux.scala 46:16:@14543.4]
  assign _T_16703 = 6'h2 == _T_11317_57; // @[Mux.scala 46:19:@14544.4]
  assign _T_16704 = _T_16703 ? _T_10366_1 : _T_16702; // @[Mux.scala 46:16:@14545.4]
  assign _T_16705 = 6'h1 == _T_11317_57; // @[Mux.scala 46:19:@14546.4]
  assign _T_16706 = _T_16705 ? _T_10366_0 : _T_16704; // @[Mux.scala 46:16:@14547.4]
  assign _T_16767 = 6'h3b == _T_11317_58; // @[Mux.scala 46:19:@14549.4]
  assign _T_16768 = _T_16767 ? _T_10366_58 : 8'h0; // @[Mux.scala 46:16:@14550.4]
  assign _T_16769 = 6'h3a == _T_11317_58; // @[Mux.scala 46:19:@14551.4]
  assign _T_16770 = _T_16769 ? _T_10366_57 : _T_16768; // @[Mux.scala 46:16:@14552.4]
  assign _T_16771 = 6'h39 == _T_11317_58; // @[Mux.scala 46:19:@14553.4]
  assign _T_16772 = _T_16771 ? _T_10366_56 : _T_16770; // @[Mux.scala 46:16:@14554.4]
  assign _T_16773 = 6'h38 == _T_11317_58; // @[Mux.scala 46:19:@14555.4]
  assign _T_16774 = _T_16773 ? _T_10366_55 : _T_16772; // @[Mux.scala 46:16:@14556.4]
  assign _T_16775 = 6'h37 == _T_11317_58; // @[Mux.scala 46:19:@14557.4]
  assign _T_16776 = _T_16775 ? _T_10366_54 : _T_16774; // @[Mux.scala 46:16:@14558.4]
  assign _T_16777 = 6'h36 == _T_11317_58; // @[Mux.scala 46:19:@14559.4]
  assign _T_16778 = _T_16777 ? _T_10366_53 : _T_16776; // @[Mux.scala 46:16:@14560.4]
  assign _T_16779 = 6'h35 == _T_11317_58; // @[Mux.scala 46:19:@14561.4]
  assign _T_16780 = _T_16779 ? _T_10366_52 : _T_16778; // @[Mux.scala 46:16:@14562.4]
  assign _T_16781 = 6'h34 == _T_11317_58; // @[Mux.scala 46:19:@14563.4]
  assign _T_16782 = _T_16781 ? _T_10366_51 : _T_16780; // @[Mux.scala 46:16:@14564.4]
  assign _T_16783 = 6'h33 == _T_11317_58; // @[Mux.scala 46:19:@14565.4]
  assign _T_16784 = _T_16783 ? _T_10366_50 : _T_16782; // @[Mux.scala 46:16:@14566.4]
  assign _T_16785 = 6'h32 == _T_11317_58; // @[Mux.scala 46:19:@14567.4]
  assign _T_16786 = _T_16785 ? _T_10366_49 : _T_16784; // @[Mux.scala 46:16:@14568.4]
  assign _T_16787 = 6'h31 == _T_11317_58; // @[Mux.scala 46:19:@14569.4]
  assign _T_16788 = _T_16787 ? _T_10366_48 : _T_16786; // @[Mux.scala 46:16:@14570.4]
  assign _T_16789 = 6'h30 == _T_11317_58; // @[Mux.scala 46:19:@14571.4]
  assign _T_16790 = _T_16789 ? _T_10366_47 : _T_16788; // @[Mux.scala 46:16:@14572.4]
  assign _T_16791 = 6'h2f == _T_11317_58; // @[Mux.scala 46:19:@14573.4]
  assign _T_16792 = _T_16791 ? _T_10366_46 : _T_16790; // @[Mux.scala 46:16:@14574.4]
  assign _T_16793 = 6'h2e == _T_11317_58; // @[Mux.scala 46:19:@14575.4]
  assign _T_16794 = _T_16793 ? _T_10366_45 : _T_16792; // @[Mux.scala 46:16:@14576.4]
  assign _T_16795 = 6'h2d == _T_11317_58; // @[Mux.scala 46:19:@14577.4]
  assign _T_16796 = _T_16795 ? _T_10366_44 : _T_16794; // @[Mux.scala 46:16:@14578.4]
  assign _T_16797 = 6'h2c == _T_11317_58; // @[Mux.scala 46:19:@14579.4]
  assign _T_16798 = _T_16797 ? _T_10366_43 : _T_16796; // @[Mux.scala 46:16:@14580.4]
  assign _T_16799 = 6'h2b == _T_11317_58; // @[Mux.scala 46:19:@14581.4]
  assign _T_16800 = _T_16799 ? _T_10366_42 : _T_16798; // @[Mux.scala 46:16:@14582.4]
  assign _T_16801 = 6'h2a == _T_11317_58; // @[Mux.scala 46:19:@14583.4]
  assign _T_16802 = _T_16801 ? _T_10366_41 : _T_16800; // @[Mux.scala 46:16:@14584.4]
  assign _T_16803 = 6'h29 == _T_11317_58; // @[Mux.scala 46:19:@14585.4]
  assign _T_16804 = _T_16803 ? _T_10366_40 : _T_16802; // @[Mux.scala 46:16:@14586.4]
  assign _T_16805 = 6'h28 == _T_11317_58; // @[Mux.scala 46:19:@14587.4]
  assign _T_16806 = _T_16805 ? _T_10366_39 : _T_16804; // @[Mux.scala 46:16:@14588.4]
  assign _T_16807 = 6'h27 == _T_11317_58; // @[Mux.scala 46:19:@14589.4]
  assign _T_16808 = _T_16807 ? _T_10366_38 : _T_16806; // @[Mux.scala 46:16:@14590.4]
  assign _T_16809 = 6'h26 == _T_11317_58; // @[Mux.scala 46:19:@14591.4]
  assign _T_16810 = _T_16809 ? _T_10366_37 : _T_16808; // @[Mux.scala 46:16:@14592.4]
  assign _T_16811 = 6'h25 == _T_11317_58; // @[Mux.scala 46:19:@14593.4]
  assign _T_16812 = _T_16811 ? _T_10366_36 : _T_16810; // @[Mux.scala 46:16:@14594.4]
  assign _T_16813 = 6'h24 == _T_11317_58; // @[Mux.scala 46:19:@14595.4]
  assign _T_16814 = _T_16813 ? _T_10366_35 : _T_16812; // @[Mux.scala 46:16:@14596.4]
  assign _T_16815 = 6'h23 == _T_11317_58; // @[Mux.scala 46:19:@14597.4]
  assign _T_16816 = _T_16815 ? _T_10366_34 : _T_16814; // @[Mux.scala 46:16:@14598.4]
  assign _T_16817 = 6'h22 == _T_11317_58; // @[Mux.scala 46:19:@14599.4]
  assign _T_16818 = _T_16817 ? _T_10366_33 : _T_16816; // @[Mux.scala 46:16:@14600.4]
  assign _T_16819 = 6'h21 == _T_11317_58; // @[Mux.scala 46:19:@14601.4]
  assign _T_16820 = _T_16819 ? _T_10366_32 : _T_16818; // @[Mux.scala 46:16:@14602.4]
  assign _T_16821 = 6'h20 == _T_11317_58; // @[Mux.scala 46:19:@14603.4]
  assign _T_16822 = _T_16821 ? _T_10366_31 : _T_16820; // @[Mux.scala 46:16:@14604.4]
  assign _T_16823 = 6'h1f == _T_11317_58; // @[Mux.scala 46:19:@14605.4]
  assign _T_16824 = _T_16823 ? _T_10366_30 : _T_16822; // @[Mux.scala 46:16:@14606.4]
  assign _T_16825 = 6'h1e == _T_11317_58; // @[Mux.scala 46:19:@14607.4]
  assign _T_16826 = _T_16825 ? _T_10366_29 : _T_16824; // @[Mux.scala 46:16:@14608.4]
  assign _T_16827 = 6'h1d == _T_11317_58; // @[Mux.scala 46:19:@14609.4]
  assign _T_16828 = _T_16827 ? _T_10366_28 : _T_16826; // @[Mux.scala 46:16:@14610.4]
  assign _T_16829 = 6'h1c == _T_11317_58; // @[Mux.scala 46:19:@14611.4]
  assign _T_16830 = _T_16829 ? _T_10366_27 : _T_16828; // @[Mux.scala 46:16:@14612.4]
  assign _T_16831 = 6'h1b == _T_11317_58; // @[Mux.scala 46:19:@14613.4]
  assign _T_16832 = _T_16831 ? _T_10366_26 : _T_16830; // @[Mux.scala 46:16:@14614.4]
  assign _T_16833 = 6'h1a == _T_11317_58; // @[Mux.scala 46:19:@14615.4]
  assign _T_16834 = _T_16833 ? _T_10366_25 : _T_16832; // @[Mux.scala 46:16:@14616.4]
  assign _T_16835 = 6'h19 == _T_11317_58; // @[Mux.scala 46:19:@14617.4]
  assign _T_16836 = _T_16835 ? _T_10366_24 : _T_16834; // @[Mux.scala 46:16:@14618.4]
  assign _T_16837 = 6'h18 == _T_11317_58; // @[Mux.scala 46:19:@14619.4]
  assign _T_16838 = _T_16837 ? _T_10366_23 : _T_16836; // @[Mux.scala 46:16:@14620.4]
  assign _T_16839 = 6'h17 == _T_11317_58; // @[Mux.scala 46:19:@14621.4]
  assign _T_16840 = _T_16839 ? _T_10366_22 : _T_16838; // @[Mux.scala 46:16:@14622.4]
  assign _T_16841 = 6'h16 == _T_11317_58; // @[Mux.scala 46:19:@14623.4]
  assign _T_16842 = _T_16841 ? _T_10366_21 : _T_16840; // @[Mux.scala 46:16:@14624.4]
  assign _T_16843 = 6'h15 == _T_11317_58; // @[Mux.scala 46:19:@14625.4]
  assign _T_16844 = _T_16843 ? _T_10366_20 : _T_16842; // @[Mux.scala 46:16:@14626.4]
  assign _T_16845 = 6'h14 == _T_11317_58; // @[Mux.scala 46:19:@14627.4]
  assign _T_16846 = _T_16845 ? _T_10366_19 : _T_16844; // @[Mux.scala 46:16:@14628.4]
  assign _T_16847 = 6'h13 == _T_11317_58; // @[Mux.scala 46:19:@14629.4]
  assign _T_16848 = _T_16847 ? _T_10366_18 : _T_16846; // @[Mux.scala 46:16:@14630.4]
  assign _T_16849 = 6'h12 == _T_11317_58; // @[Mux.scala 46:19:@14631.4]
  assign _T_16850 = _T_16849 ? _T_10366_17 : _T_16848; // @[Mux.scala 46:16:@14632.4]
  assign _T_16851 = 6'h11 == _T_11317_58; // @[Mux.scala 46:19:@14633.4]
  assign _T_16852 = _T_16851 ? _T_10366_16 : _T_16850; // @[Mux.scala 46:16:@14634.4]
  assign _T_16853 = 6'h10 == _T_11317_58; // @[Mux.scala 46:19:@14635.4]
  assign _T_16854 = _T_16853 ? _T_10366_15 : _T_16852; // @[Mux.scala 46:16:@14636.4]
  assign _T_16855 = 6'hf == _T_11317_58; // @[Mux.scala 46:19:@14637.4]
  assign _T_16856 = _T_16855 ? _T_10366_14 : _T_16854; // @[Mux.scala 46:16:@14638.4]
  assign _T_16857 = 6'he == _T_11317_58; // @[Mux.scala 46:19:@14639.4]
  assign _T_16858 = _T_16857 ? _T_10366_13 : _T_16856; // @[Mux.scala 46:16:@14640.4]
  assign _T_16859 = 6'hd == _T_11317_58; // @[Mux.scala 46:19:@14641.4]
  assign _T_16860 = _T_16859 ? _T_10366_12 : _T_16858; // @[Mux.scala 46:16:@14642.4]
  assign _T_16861 = 6'hc == _T_11317_58; // @[Mux.scala 46:19:@14643.4]
  assign _T_16862 = _T_16861 ? _T_10366_11 : _T_16860; // @[Mux.scala 46:16:@14644.4]
  assign _T_16863 = 6'hb == _T_11317_58; // @[Mux.scala 46:19:@14645.4]
  assign _T_16864 = _T_16863 ? _T_10366_10 : _T_16862; // @[Mux.scala 46:16:@14646.4]
  assign _T_16865 = 6'ha == _T_11317_58; // @[Mux.scala 46:19:@14647.4]
  assign _T_16866 = _T_16865 ? _T_10366_9 : _T_16864; // @[Mux.scala 46:16:@14648.4]
  assign _T_16867 = 6'h9 == _T_11317_58; // @[Mux.scala 46:19:@14649.4]
  assign _T_16868 = _T_16867 ? _T_10366_8 : _T_16866; // @[Mux.scala 46:16:@14650.4]
  assign _T_16869 = 6'h8 == _T_11317_58; // @[Mux.scala 46:19:@14651.4]
  assign _T_16870 = _T_16869 ? _T_10366_7 : _T_16868; // @[Mux.scala 46:16:@14652.4]
  assign _T_16871 = 6'h7 == _T_11317_58; // @[Mux.scala 46:19:@14653.4]
  assign _T_16872 = _T_16871 ? _T_10366_6 : _T_16870; // @[Mux.scala 46:16:@14654.4]
  assign _T_16873 = 6'h6 == _T_11317_58; // @[Mux.scala 46:19:@14655.4]
  assign _T_16874 = _T_16873 ? _T_10366_5 : _T_16872; // @[Mux.scala 46:16:@14656.4]
  assign _T_16875 = 6'h5 == _T_11317_58; // @[Mux.scala 46:19:@14657.4]
  assign _T_16876 = _T_16875 ? _T_10366_4 : _T_16874; // @[Mux.scala 46:16:@14658.4]
  assign _T_16877 = 6'h4 == _T_11317_58; // @[Mux.scala 46:19:@14659.4]
  assign _T_16878 = _T_16877 ? _T_10366_3 : _T_16876; // @[Mux.scala 46:16:@14660.4]
  assign _T_16879 = 6'h3 == _T_11317_58; // @[Mux.scala 46:19:@14661.4]
  assign _T_16880 = _T_16879 ? _T_10366_2 : _T_16878; // @[Mux.scala 46:16:@14662.4]
  assign _T_16881 = 6'h2 == _T_11317_58; // @[Mux.scala 46:19:@14663.4]
  assign _T_16882 = _T_16881 ? _T_10366_1 : _T_16880; // @[Mux.scala 46:16:@14664.4]
  assign _T_16883 = 6'h1 == _T_11317_58; // @[Mux.scala 46:19:@14665.4]
  assign _T_16884 = _T_16883 ? _T_10366_0 : _T_16882; // @[Mux.scala 46:16:@14666.4]
  assign _T_16946 = 6'h3c == _T_11317_59; // @[Mux.scala 46:19:@14668.4]
  assign _T_16947 = _T_16946 ? _T_10366_59 : 8'h0; // @[Mux.scala 46:16:@14669.4]
  assign _T_16948 = 6'h3b == _T_11317_59; // @[Mux.scala 46:19:@14670.4]
  assign _T_16949 = _T_16948 ? _T_10366_58 : _T_16947; // @[Mux.scala 46:16:@14671.4]
  assign _T_16950 = 6'h3a == _T_11317_59; // @[Mux.scala 46:19:@14672.4]
  assign _T_16951 = _T_16950 ? _T_10366_57 : _T_16949; // @[Mux.scala 46:16:@14673.4]
  assign _T_16952 = 6'h39 == _T_11317_59; // @[Mux.scala 46:19:@14674.4]
  assign _T_16953 = _T_16952 ? _T_10366_56 : _T_16951; // @[Mux.scala 46:16:@14675.4]
  assign _T_16954 = 6'h38 == _T_11317_59; // @[Mux.scala 46:19:@14676.4]
  assign _T_16955 = _T_16954 ? _T_10366_55 : _T_16953; // @[Mux.scala 46:16:@14677.4]
  assign _T_16956 = 6'h37 == _T_11317_59; // @[Mux.scala 46:19:@14678.4]
  assign _T_16957 = _T_16956 ? _T_10366_54 : _T_16955; // @[Mux.scala 46:16:@14679.4]
  assign _T_16958 = 6'h36 == _T_11317_59; // @[Mux.scala 46:19:@14680.4]
  assign _T_16959 = _T_16958 ? _T_10366_53 : _T_16957; // @[Mux.scala 46:16:@14681.4]
  assign _T_16960 = 6'h35 == _T_11317_59; // @[Mux.scala 46:19:@14682.4]
  assign _T_16961 = _T_16960 ? _T_10366_52 : _T_16959; // @[Mux.scala 46:16:@14683.4]
  assign _T_16962 = 6'h34 == _T_11317_59; // @[Mux.scala 46:19:@14684.4]
  assign _T_16963 = _T_16962 ? _T_10366_51 : _T_16961; // @[Mux.scala 46:16:@14685.4]
  assign _T_16964 = 6'h33 == _T_11317_59; // @[Mux.scala 46:19:@14686.4]
  assign _T_16965 = _T_16964 ? _T_10366_50 : _T_16963; // @[Mux.scala 46:16:@14687.4]
  assign _T_16966 = 6'h32 == _T_11317_59; // @[Mux.scala 46:19:@14688.4]
  assign _T_16967 = _T_16966 ? _T_10366_49 : _T_16965; // @[Mux.scala 46:16:@14689.4]
  assign _T_16968 = 6'h31 == _T_11317_59; // @[Mux.scala 46:19:@14690.4]
  assign _T_16969 = _T_16968 ? _T_10366_48 : _T_16967; // @[Mux.scala 46:16:@14691.4]
  assign _T_16970 = 6'h30 == _T_11317_59; // @[Mux.scala 46:19:@14692.4]
  assign _T_16971 = _T_16970 ? _T_10366_47 : _T_16969; // @[Mux.scala 46:16:@14693.4]
  assign _T_16972 = 6'h2f == _T_11317_59; // @[Mux.scala 46:19:@14694.4]
  assign _T_16973 = _T_16972 ? _T_10366_46 : _T_16971; // @[Mux.scala 46:16:@14695.4]
  assign _T_16974 = 6'h2e == _T_11317_59; // @[Mux.scala 46:19:@14696.4]
  assign _T_16975 = _T_16974 ? _T_10366_45 : _T_16973; // @[Mux.scala 46:16:@14697.4]
  assign _T_16976 = 6'h2d == _T_11317_59; // @[Mux.scala 46:19:@14698.4]
  assign _T_16977 = _T_16976 ? _T_10366_44 : _T_16975; // @[Mux.scala 46:16:@14699.4]
  assign _T_16978 = 6'h2c == _T_11317_59; // @[Mux.scala 46:19:@14700.4]
  assign _T_16979 = _T_16978 ? _T_10366_43 : _T_16977; // @[Mux.scala 46:16:@14701.4]
  assign _T_16980 = 6'h2b == _T_11317_59; // @[Mux.scala 46:19:@14702.4]
  assign _T_16981 = _T_16980 ? _T_10366_42 : _T_16979; // @[Mux.scala 46:16:@14703.4]
  assign _T_16982 = 6'h2a == _T_11317_59; // @[Mux.scala 46:19:@14704.4]
  assign _T_16983 = _T_16982 ? _T_10366_41 : _T_16981; // @[Mux.scala 46:16:@14705.4]
  assign _T_16984 = 6'h29 == _T_11317_59; // @[Mux.scala 46:19:@14706.4]
  assign _T_16985 = _T_16984 ? _T_10366_40 : _T_16983; // @[Mux.scala 46:16:@14707.4]
  assign _T_16986 = 6'h28 == _T_11317_59; // @[Mux.scala 46:19:@14708.4]
  assign _T_16987 = _T_16986 ? _T_10366_39 : _T_16985; // @[Mux.scala 46:16:@14709.4]
  assign _T_16988 = 6'h27 == _T_11317_59; // @[Mux.scala 46:19:@14710.4]
  assign _T_16989 = _T_16988 ? _T_10366_38 : _T_16987; // @[Mux.scala 46:16:@14711.4]
  assign _T_16990 = 6'h26 == _T_11317_59; // @[Mux.scala 46:19:@14712.4]
  assign _T_16991 = _T_16990 ? _T_10366_37 : _T_16989; // @[Mux.scala 46:16:@14713.4]
  assign _T_16992 = 6'h25 == _T_11317_59; // @[Mux.scala 46:19:@14714.4]
  assign _T_16993 = _T_16992 ? _T_10366_36 : _T_16991; // @[Mux.scala 46:16:@14715.4]
  assign _T_16994 = 6'h24 == _T_11317_59; // @[Mux.scala 46:19:@14716.4]
  assign _T_16995 = _T_16994 ? _T_10366_35 : _T_16993; // @[Mux.scala 46:16:@14717.4]
  assign _T_16996 = 6'h23 == _T_11317_59; // @[Mux.scala 46:19:@14718.4]
  assign _T_16997 = _T_16996 ? _T_10366_34 : _T_16995; // @[Mux.scala 46:16:@14719.4]
  assign _T_16998 = 6'h22 == _T_11317_59; // @[Mux.scala 46:19:@14720.4]
  assign _T_16999 = _T_16998 ? _T_10366_33 : _T_16997; // @[Mux.scala 46:16:@14721.4]
  assign _T_17000 = 6'h21 == _T_11317_59; // @[Mux.scala 46:19:@14722.4]
  assign _T_17001 = _T_17000 ? _T_10366_32 : _T_16999; // @[Mux.scala 46:16:@14723.4]
  assign _T_17002 = 6'h20 == _T_11317_59; // @[Mux.scala 46:19:@14724.4]
  assign _T_17003 = _T_17002 ? _T_10366_31 : _T_17001; // @[Mux.scala 46:16:@14725.4]
  assign _T_17004 = 6'h1f == _T_11317_59; // @[Mux.scala 46:19:@14726.4]
  assign _T_17005 = _T_17004 ? _T_10366_30 : _T_17003; // @[Mux.scala 46:16:@14727.4]
  assign _T_17006 = 6'h1e == _T_11317_59; // @[Mux.scala 46:19:@14728.4]
  assign _T_17007 = _T_17006 ? _T_10366_29 : _T_17005; // @[Mux.scala 46:16:@14729.4]
  assign _T_17008 = 6'h1d == _T_11317_59; // @[Mux.scala 46:19:@14730.4]
  assign _T_17009 = _T_17008 ? _T_10366_28 : _T_17007; // @[Mux.scala 46:16:@14731.4]
  assign _T_17010 = 6'h1c == _T_11317_59; // @[Mux.scala 46:19:@14732.4]
  assign _T_17011 = _T_17010 ? _T_10366_27 : _T_17009; // @[Mux.scala 46:16:@14733.4]
  assign _T_17012 = 6'h1b == _T_11317_59; // @[Mux.scala 46:19:@14734.4]
  assign _T_17013 = _T_17012 ? _T_10366_26 : _T_17011; // @[Mux.scala 46:16:@14735.4]
  assign _T_17014 = 6'h1a == _T_11317_59; // @[Mux.scala 46:19:@14736.4]
  assign _T_17015 = _T_17014 ? _T_10366_25 : _T_17013; // @[Mux.scala 46:16:@14737.4]
  assign _T_17016 = 6'h19 == _T_11317_59; // @[Mux.scala 46:19:@14738.4]
  assign _T_17017 = _T_17016 ? _T_10366_24 : _T_17015; // @[Mux.scala 46:16:@14739.4]
  assign _T_17018 = 6'h18 == _T_11317_59; // @[Mux.scala 46:19:@14740.4]
  assign _T_17019 = _T_17018 ? _T_10366_23 : _T_17017; // @[Mux.scala 46:16:@14741.4]
  assign _T_17020 = 6'h17 == _T_11317_59; // @[Mux.scala 46:19:@14742.4]
  assign _T_17021 = _T_17020 ? _T_10366_22 : _T_17019; // @[Mux.scala 46:16:@14743.4]
  assign _T_17022 = 6'h16 == _T_11317_59; // @[Mux.scala 46:19:@14744.4]
  assign _T_17023 = _T_17022 ? _T_10366_21 : _T_17021; // @[Mux.scala 46:16:@14745.4]
  assign _T_17024 = 6'h15 == _T_11317_59; // @[Mux.scala 46:19:@14746.4]
  assign _T_17025 = _T_17024 ? _T_10366_20 : _T_17023; // @[Mux.scala 46:16:@14747.4]
  assign _T_17026 = 6'h14 == _T_11317_59; // @[Mux.scala 46:19:@14748.4]
  assign _T_17027 = _T_17026 ? _T_10366_19 : _T_17025; // @[Mux.scala 46:16:@14749.4]
  assign _T_17028 = 6'h13 == _T_11317_59; // @[Mux.scala 46:19:@14750.4]
  assign _T_17029 = _T_17028 ? _T_10366_18 : _T_17027; // @[Mux.scala 46:16:@14751.4]
  assign _T_17030 = 6'h12 == _T_11317_59; // @[Mux.scala 46:19:@14752.4]
  assign _T_17031 = _T_17030 ? _T_10366_17 : _T_17029; // @[Mux.scala 46:16:@14753.4]
  assign _T_17032 = 6'h11 == _T_11317_59; // @[Mux.scala 46:19:@14754.4]
  assign _T_17033 = _T_17032 ? _T_10366_16 : _T_17031; // @[Mux.scala 46:16:@14755.4]
  assign _T_17034 = 6'h10 == _T_11317_59; // @[Mux.scala 46:19:@14756.4]
  assign _T_17035 = _T_17034 ? _T_10366_15 : _T_17033; // @[Mux.scala 46:16:@14757.4]
  assign _T_17036 = 6'hf == _T_11317_59; // @[Mux.scala 46:19:@14758.4]
  assign _T_17037 = _T_17036 ? _T_10366_14 : _T_17035; // @[Mux.scala 46:16:@14759.4]
  assign _T_17038 = 6'he == _T_11317_59; // @[Mux.scala 46:19:@14760.4]
  assign _T_17039 = _T_17038 ? _T_10366_13 : _T_17037; // @[Mux.scala 46:16:@14761.4]
  assign _T_17040 = 6'hd == _T_11317_59; // @[Mux.scala 46:19:@14762.4]
  assign _T_17041 = _T_17040 ? _T_10366_12 : _T_17039; // @[Mux.scala 46:16:@14763.4]
  assign _T_17042 = 6'hc == _T_11317_59; // @[Mux.scala 46:19:@14764.4]
  assign _T_17043 = _T_17042 ? _T_10366_11 : _T_17041; // @[Mux.scala 46:16:@14765.4]
  assign _T_17044 = 6'hb == _T_11317_59; // @[Mux.scala 46:19:@14766.4]
  assign _T_17045 = _T_17044 ? _T_10366_10 : _T_17043; // @[Mux.scala 46:16:@14767.4]
  assign _T_17046 = 6'ha == _T_11317_59; // @[Mux.scala 46:19:@14768.4]
  assign _T_17047 = _T_17046 ? _T_10366_9 : _T_17045; // @[Mux.scala 46:16:@14769.4]
  assign _T_17048 = 6'h9 == _T_11317_59; // @[Mux.scala 46:19:@14770.4]
  assign _T_17049 = _T_17048 ? _T_10366_8 : _T_17047; // @[Mux.scala 46:16:@14771.4]
  assign _T_17050 = 6'h8 == _T_11317_59; // @[Mux.scala 46:19:@14772.4]
  assign _T_17051 = _T_17050 ? _T_10366_7 : _T_17049; // @[Mux.scala 46:16:@14773.4]
  assign _T_17052 = 6'h7 == _T_11317_59; // @[Mux.scala 46:19:@14774.4]
  assign _T_17053 = _T_17052 ? _T_10366_6 : _T_17051; // @[Mux.scala 46:16:@14775.4]
  assign _T_17054 = 6'h6 == _T_11317_59; // @[Mux.scala 46:19:@14776.4]
  assign _T_17055 = _T_17054 ? _T_10366_5 : _T_17053; // @[Mux.scala 46:16:@14777.4]
  assign _T_17056 = 6'h5 == _T_11317_59; // @[Mux.scala 46:19:@14778.4]
  assign _T_17057 = _T_17056 ? _T_10366_4 : _T_17055; // @[Mux.scala 46:16:@14779.4]
  assign _T_17058 = 6'h4 == _T_11317_59; // @[Mux.scala 46:19:@14780.4]
  assign _T_17059 = _T_17058 ? _T_10366_3 : _T_17057; // @[Mux.scala 46:16:@14781.4]
  assign _T_17060 = 6'h3 == _T_11317_59; // @[Mux.scala 46:19:@14782.4]
  assign _T_17061 = _T_17060 ? _T_10366_2 : _T_17059; // @[Mux.scala 46:16:@14783.4]
  assign _T_17062 = 6'h2 == _T_11317_59; // @[Mux.scala 46:19:@14784.4]
  assign _T_17063 = _T_17062 ? _T_10366_1 : _T_17061; // @[Mux.scala 46:16:@14785.4]
  assign _T_17064 = 6'h1 == _T_11317_59; // @[Mux.scala 46:19:@14786.4]
  assign _T_17065 = _T_17064 ? _T_10366_0 : _T_17063; // @[Mux.scala 46:16:@14787.4]
  assign _T_17128 = 6'h3d == _T_11317_60; // @[Mux.scala 46:19:@14789.4]
  assign _T_17129 = _T_17128 ? _T_10366_60 : 8'h0; // @[Mux.scala 46:16:@14790.4]
  assign _T_17130 = 6'h3c == _T_11317_60; // @[Mux.scala 46:19:@14791.4]
  assign _T_17131 = _T_17130 ? _T_10366_59 : _T_17129; // @[Mux.scala 46:16:@14792.4]
  assign _T_17132 = 6'h3b == _T_11317_60; // @[Mux.scala 46:19:@14793.4]
  assign _T_17133 = _T_17132 ? _T_10366_58 : _T_17131; // @[Mux.scala 46:16:@14794.4]
  assign _T_17134 = 6'h3a == _T_11317_60; // @[Mux.scala 46:19:@14795.4]
  assign _T_17135 = _T_17134 ? _T_10366_57 : _T_17133; // @[Mux.scala 46:16:@14796.4]
  assign _T_17136 = 6'h39 == _T_11317_60; // @[Mux.scala 46:19:@14797.4]
  assign _T_17137 = _T_17136 ? _T_10366_56 : _T_17135; // @[Mux.scala 46:16:@14798.4]
  assign _T_17138 = 6'h38 == _T_11317_60; // @[Mux.scala 46:19:@14799.4]
  assign _T_17139 = _T_17138 ? _T_10366_55 : _T_17137; // @[Mux.scala 46:16:@14800.4]
  assign _T_17140 = 6'h37 == _T_11317_60; // @[Mux.scala 46:19:@14801.4]
  assign _T_17141 = _T_17140 ? _T_10366_54 : _T_17139; // @[Mux.scala 46:16:@14802.4]
  assign _T_17142 = 6'h36 == _T_11317_60; // @[Mux.scala 46:19:@14803.4]
  assign _T_17143 = _T_17142 ? _T_10366_53 : _T_17141; // @[Mux.scala 46:16:@14804.4]
  assign _T_17144 = 6'h35 == _T_11317_60; // @[Mux.scala 46:19:@14805.4]
  assign _T_17145 = _T_17144 ? _T_10366_52 : _T_17143; // @[Mux.scala 46:16:@14806.4]
  assign _T_17146 = 6'h34 == _T_11317_60; // @[Mux.scala 46:19:@14807.4]
  assign _T_17147 = _T_17146 ? _T_10366_51 : _T_17145; // @[Mux.scala 46:16:@14808.4]
  assign _T_17148 = 6'h33 == _T_11317_60; // @[Mux.scala 46:19:@14809.4]
  assign _T_17149 = _T_17148 ? _T_10366_50 : _T_17147; // @[Mux.scala 46:16:@14810.4]
  assign _T_17150 = 6'h32 == _T_11317_60; // @[Mux.scala 46:19:@14811.4]
  assign _T_17151 = _T_17150 ? _T_10366_49 : _T_17149; // @[Mux.scala 46:16:@14812.4]
  assign _T_17152 = 6'h31 == _T_11317_60; // @[Mux.scala 46:19:@14813.4]
  assign _T_17153 = _T_17152 ? _T_10366_48 : _T_17151; // @[Mux.scala 46:16:@14814.4]
  assign _T_17154 = 6'h30 == _T_11317_60; // @[Mux.scala 46:19:@14815.4]
  assign _T_17155 = _T_17154 ? _T_10366_47 : _T_17153; // @[Mux.scala 46:16:@14816.4]
  assign _T_17156 = 6'h2f == _T_11317_60; // @[Mux.scala 46:19:@14817.4]
  assign _T_17157 = _T_17156 ? _T_10366_46 : _T_17155; // @[Mux.scala 46:16:@14818.4]
  assign _T_17158 = 6'h2e == _T_11317_60; // @[Mux.scala 46:19:@14819.4]
  assign _T_17159 = _T_17158 ? _T_10366_45 : _T_17157; // @[Mux.scala 46:16:@14820.4]
  assign _T_17160 = 6'h2d == _T_11317_60; // @[Mux.scala 46:19:@14821.4]
  assign _T_17161 = _T_17160 ? _T_10366_44 : _T_17159; // @[Mux.scala 46:16:@14822.4]
  assign _T_17162 = 6'h2c == _T_11317_60; // @[Mux.scala 46:19:@14823.4]
  assign _T_17163 = _T_17162 ? _T_10366_43 : _T_17161; // @[Mux.scala 46:16:@14824.4]
  assign _T_17164 = 6'h2b == _T_11317_60; // @[Mux.scala 46:19:@14825.4]
  assign _T_17165 = _T_17164 ? _T_10366_42 : _T_17163; // @[Mux.scala 46:16:@14826.4]
  assign _T_17166 = 6'h2a == _T_11317_60; // @[Mux.scala 46:19:@14827.4]
  assign _T_17167 = _T_17166 ? _T_10366_41 : _T_17165; // @[Mux.scala 46:16:@14828.4]
  assign _T_17168 = 6'h29 == _T_11317_60; // @[Mux.scala 46:19:@14829.4]
  assign _T_17169 = _T_17168 ? _T_10366_40 : _T_17167; // @[Mux.scala 46:16:@14830.4]
  assign _T_17170 = 6'h28 == _T_11317_60; // @[Mux.scala 46:19:@14831.4]
  assign _T_17171 = _T_17170 ? _T_10366_39 : _T_17169; // @[Mux.scala 46:16:@14832.4]
  assign _T_17172 = 6'h27 == _T_11317_60; // @[Mux.scala 46:19:@14833.4]
  assign _T_17173 = _T_17172 ? _T_10366_38 : _T_17171; // @[Mux.scala 46:16:@14834.4]
  assign _T_17174 = 6'h26 == _T_11317_60; // @[Mux.scala 46:19:@14835.4]
  assign _T_17175 = _T_17174 ? _T_10366_37 : _T_17173; // @[Mux.scala 46:16:@14836.4]
  assign _T_17176 = 6'h25 == _T_11317_60; // @[Mux.scala 46:19:@14837.4]
  assign _T_17177 = _T_17176 ? _T_10366_36 : _T_17175; // @[Mux.scala 46:16:@14838.4]
  assign _T_17178 = 6'h24 == _T_11317_60; // @[Mux.scala 46:19:@14839.4]
  assign _T_17179 = _T_17178 ? _T_10366_35 : _T_17177; // @[Mux.scala 46:16:@14840.4]
  assign _T_17180 = 6'h23 == _T_11317_60; // @[Mux.scala 46:19:@14841.4]
  assign _T_17181 = _T_17180 ? _T_10366_34 : _T_17179; // @[Mux.scala 46:16:@14842.4]
  assign _T_17182 = 6'h22 == _T_11317_60; // @[Mux.scala 46:19:@14843.4]
  assign _T_17183 = _T_17182 ? _T_10366_33 : _T_17181; // @[Mux.scala 46:16:@14844.4]
  assign _T_17184 = 6'h21 == _T_11317_60; // @[Mux.scala 46:19:@14845.4]
  assign _T_17185 = _T_17184 ? _T_10366_32 : _T_17183; // @[Mux.scala 46:16:@14846.4]
  assign _T_17186 = 6'h20 == _T_11317_60; // @[Mux.scala 46:19:@14847.4]
  assign _T_17187 = _T_17186 ? _T_10366_31 : _T_17185; // @[Mux.scala 46:16:@14848.4]
  assign _T_17188 = 6'h1f == _T_11317_60; // @[Mux.scala 46:19:@14849.4]
  assign _T_17189 = _T_17188 ? _T_10366_30 : _T_17187; // @[Mux.scala 46:16:@14850.4]
  assign _T_17190 = 6'h1e == _T_11317_60; // @[Mux.scala 46:19:@14851.4]
  assign _T_17191 = _T_17190 ? _T_10366_29 : _T_17189; // @[Mux.scala 46:16:@14852.4]
  assign _T_17192 = 6'h1d == _T_11317_60; // @[Mux.scala 46:19:@14853.4]
  assign _T_17193 = _T_17192 ? _T_10366_28 : _T_17191; // @[Mux.scala 46:16:@14854.4]
  assign _T_17194 = 6'h1c == _T_11317_60; // @[Mux.scala 46:19:@14855.4]
  assign _T_17195 = _T_17194 ? _T_10366_27 : _T_17193; // @[Mux.scala 46:16:@14856.4]
  assign _T_17196 = 6'h1b == _T_11317_60; // @[Mux.scala 46:19:@14857.4]
  assign _T_17197 = _T_17196 ? _T_10366_26 : _T_17195; // @[Mux.scala 46:16:@14858.4]
  assign _T_17198 = 6'h1a == _T_11317_60; // @[Mux.scala 46:19:@14859.4]
  assign _T_17199 = _T_17198 ? _T_10366_25 : _T_17197; // @[Mux.scala 46:16:@14860.4]
  assign _T_17200 = 6'h19 == _T_11317_60; // @[Mux.scala 46:19:@14861.4]
  assign _T_17201 = _T_17200 ? _T_10366_24 : _T_17199; // @[Mux.scala 46:16:@14862.4]
  assign _T_17202 = 6'h18 == _T_11317_60; // @[Mux.scala 46:19:@14863.4]
  assign _T_17203 = _T_17202 ? _T_10366_23 : _T_17201; // @[Mux.scala 46:16:@14864.4]
  assign _T_17204 = 6'h17 == _T_11317_60; // @[Mux.scala 46:19:@14865.4]
  assign _T_17205 = _T_17204 ? _T_10366_22 : _T_17203; // @[Mux.scala 46:16:@14866.4]
  assign _T_17206 = 6'h16 == _T_11317_60; // @[Mux.scala 46:19:@14867.4]
  assign _T_17207 = _T_17206 ? _T_10366_21 : _T_17205; // @[Mux.scala 46:16:@14868.4]
  assign _T_17208 = 6'h15 == _T_11317_60; // @[Mux.scala 46:19:@14869.4]
  assign _T_17209 = _T_17208 ? _T_10366_20 : _T_17207; // @[Mux.scala 46:16:@14870.4]
  assign _T_17210 = 6'h14 == _T_11317_60; // @[Mux.scala 46:19:@14871.4]
  assign _T_17211 = _T_17210 ? _T_10366_19 : _T_17209; // @[Mux.scala 46:16:@14872.4]
  assign _T_17212 = 6'h13 == _T_11317_60; // @[Mux.scala 46:19:@14873.4]
  assign _T_17213 = _T_17212 ? _T_10366_18 : _T_17211; // @[Mux.scala 46:16:@14874.4]
  assign _T_17214 = 6'h12 == _T_11317_60; // @[Mux.scala 46:19:@14875.4]
  assign _T_17215 = _T_17214 ? _T_10366_17 : _T_17213; // @[Mux.scala 46:16:@14876.4]
  assign _T_17216 = 6'h11 == _T_11317_60; // @[Mux.scala 46:19:@14877.4]
  assign _T_17217 = _T_17216 ? _T_10366_16 : _T_17215; // @[Mux.scala 46:16:@14878.4]
  assign _T_17218 = 6'h10 == _T_11317_60; // @[Mux.scala 46:19:@14879.4]
  assign _T_17219 = _T_17218 ? _T_10366_15 : _T_17217; // @[Mux.scala 46:16:@14880.4]
  assign _T_17220 = 6'hf == _T_11317_60; // @[Mux.scala 46:19:@14881.4]
  assign _T_17221 = _T_17220 ? _T_10366_14 : _T_17219; // @[Mux.scala 46:16:@14882.4]
  assign _T_17222 = 6'he == _T_11317_60; // @[Mux.scala 46:19:@14883.4]
  assign _T_17223 = _T_17222 ? _T_10366_13 : _T_17221; // @[Mux.scala 46:16:@14884.4]
  assign _T_17224 = 6'hd == _T_11317_60; // @[Mux.scala 46:19:@14885.4]
  assign _T_17225 = _T_17224 ? _T_10366_12 : _T_17223; // @[Mux.scala 46:16:@14886.4]
  assign _T_17226 = 6'hc == _T_11317_60; // @[Mux.scala 46:19:@14887.4]
  assign _T_17227 = _T_17226 ? _T_10366_11 : _T_17225; // @[Mux.scala 46:16:@14888.4]
  assign _T_17228 = 6'hb == _T_11317_60; // @[Mux.scala 46:19:@14889.4]
  assign _T_17229 = _T_17228 ? _T_10366_10 : _T_17227; // @[Mux.scala 46:16:@14890.4]
  assign _T_17230 = 6'ha == _T_11317_60; // @[Mux.scala 46:19:@14891.4]
  assign _T_17231 = _T_17230 ? _T_10366_9 : _T_17229; // @[Mux.scala 46:16:@14892.4]
  assign _T_17232 = 6'h9 == _T_11317_60; // @[Mux.scala 46:19:@14893.4]
  assign _T_17233 = _T_17232 ? _T_10366_8 : _T_17231; // @[Mux.scala 46:16:@14894.4]
  assign _T_17234 = 6'h8 == _T_11317_60; // @[Mux.scala 46:19:@14895.4]
  assign _T_17235 = _T_17234 ? _T_10366_7 : _T_17233; // @[Mux.scala 46:16:@14896.4]
  assign _T_17236 = 6'h7 == _T_11317_60; // @[Mux.scala 46:19:@14897.4]
  assign _T_17237 = _T_17236 ? _T_10366_6 : _T_17235; // @[Mux.scala 46:16:@14898.4]
  assign _T_17238 = 6'h6 == _T_11317_60; // @[Mux.scala 46:19:@14899.4]
  assign _T_17239 = _T_17238 ? _T_10366_5 : _T_17237; // @[Mux.scala 46:16:@14900.4]
  assign _T_17240 = 6'h5 == _T_11317_60; // @[Mux.scala 46:19:@14901.4]
  assign _T_17241 = _T_17240 ? _T_10366_4 : _T_17239; // @[Mux.scala 46:16:@14902.4]
  assign _T_17242 = 6'h4 == _T_11317_60; // @[Mux.scala 46:19:@14903.4]
  assign _T_17243 = _T_17242 ? _T_10366_3 : _T_17241; // @[Mux.scala 46:16:@14904.4]
  assign _T_17244 = 6'h3 == _T_11317_60; // @[Mux.scala 46:19:@14905.4]
  assign _T_17245 = _T_17244 ? _T_10366_2 : _T_17243; // @[Mux.scala 46:16:@14906.4]
  assign _T_17246 = 6'h2 == _T_11317_60; // @[Mux.scala 46:19:@14907.4]
  assign _T_17247 = _T_17246 ? _T_10366_1 : _T_17245; // @[Mux.scala 46:16:@14908.4]
  assign _T_17248 = 6'h1 == _T_11317_60; // @[Mux.scala 46:19:@14909.4]
  assign _T_17249 = _T_17248 ? _T_10366_0 : _T_17247; // @[Mux.scala 46:16:@14910.4]
  assign _T_17313 = 6'h3e == _T_11317_61; // @[Mux.scala 46:19:@14912.4]
  assign _T_17314 = _T_17313 ? _T_10366_61 : 8'h0; // @[Mux.scala 46:16:@14913.4]
  assign _T_17315 = 6'h3d == _T_11317_61; // @[Mux.scala 46:19:@14914.4]
  assign _T_17316 = _T_17315 ? _T_10366_60 : _T_17314; // @[Mux.scala 46:16:@14915.4]
  assign _T_17317 = 6'h3c == _T_11317_61; // @[Mux.scala 46:19:@14916.4]
  assign _T_17318 = _T_17317 ? _T_10366_59 : _T_17316; // @[Mux.scala 46:16:@14917.4]
  assign _T_17319 = 6'h3b == _T_11317_61; // @[Mux.scala 46:19:@14918.4]
  assign _T_17320 = _T_17319 ? _T_10366_58 : _T_17318; // @[Mux.scala 46:16:@14919.4]
  assign _T_17321 = 6'h3a == _T_11317_61; // @[Mux.scala 46:19:@14920.4]
  assign _T_17322 = _T_17321 ? _T_10366_57 : _T_17320; // @[Mux.scala 46:16:@14921.4]
  assign _T_17323 = 6'h39 == _T_11317_61; // @[Mux.scala 46:19:@14922.4]
  assign _T_17324 = _T_17323 ? _T_10366_56 : _T_17322; // @[Mux.scala 46:16:@14923.4]
  assign _T_17325 = 6'h38 == _T_11317_61; // @[Mux.scala 46:19:@14924.4]
  assign _T_17326 = _T_17325 ? _T_10366_55 : _T_17324; // @[Mux.scala 46:16:@14925.4]
  assign _T_17327 = 6'h37 == _T_11317_61; // @[Mux.scala 46:19:@14926.4]
  assign _T_17328 = _T_17327 ? _T_10366_54 : _T_17326; // @[Mux.scala 46:16:@14927.4]
  assign _T_17329 = 6'h36 == _T_11317_61; // @[Mux.scala 46:19:@14928.4]
  assign _T_17330 = _T_17329 ? _T_10366_53 : _T_17328; // @[Mux.scala 46:16:@14929.4]
  assign _T_17331 = 6'h35 == _T_11317_61; // @[Mux.scala 46:19:@14930.4]
  assign _T_17332 = _T_17331 ? _T_10366_52 : _T_17330; // @[Mux.scala 46:16:@14931.4]
  assign _T_17333 = 6'h34 == _T_11317_61; // @[Mux.scala 46:19:@14932.4]
  assign _T_17334 = _T_17333 ? _T_10366_51 : _T_17332; // @[Mux.scala 46:16:@14933.4]
  assign _T_17335 = 6'h33 == _T_11317_61; // @[Mux.scala 46:19:@14934.4]
  assign _T_17336 = _T_17335 ? _T_10366_50 : _T_17334; // @[Mux.scala 46:16:@14935.4]
  assign _T_17337 = 6'h32 == _T_11317_61; // @[Mux.scala 46:19:@14936.4]
  assign _T_17338 = _T_17337 ? _T_10366_49 : _T_17336; // @[Mux.scala 46:16:@14937.4]
  assign _T_17339 = 6'h31 == _T_11317_61; // @[Mux.scala 46:19:@14938.4]
  assign _T_17340 = _T_17339 ? _T_10366_48 : _T_17338; // @[Mux.scala 46:16:@14939.4]
  assign _T_17341 = 6'h30 == _T_11317_61; // @[Mux.scala 46:19:@14940.4]
  assign _T_17342 = _T_17341 ? _T_10366_47 : _T_17340; // @[Mux.scala 46:16:@14941.4]
  assign _T_17343 = 6'h2f == _T_11317_61; // @[Mux.scala 46:19:@14942.4]
  assign _T_17344 = _T_17343 ? _T_10366_46 : _T_17342; // @[Mux.scala 46:16:@14943.4]
  assign _T_17345 = 6'h2e == _T_11317_61; // @[Mux.scala 46:19:@14944.4]
  assign _T_17346 = _T_17345 ? _T_10366_45 : _T_17344; // @[Mux.scala 46:16:@14945.4]
  assign _T_17347 = 6'h2d == _T_11317_61; // @[Mux.scala 46:19:@14946.4]
  assign _T_17348 = _T_17347 ? _T_10366_44 : _T_17346; // @[Mux.scala 46:16:@14947.4]
  assign _T_17349 = 6'h2c == _T_11317_61; // @[Mux.scala 46:19:@14948.4]
  assign _T_17350 = _T_17349 ? _T_10366_43 : _T_17348; // @[Mux.scala 46:16:@14949.4]
  assign _T_17351 = 6'h2b == _T_11317_61; // @[Mux.scala 46:19:@14950.4]
  assign _T_17352 = _T_17351 ? _T_10366_42 : _T_17350; // @[Mux.scala 46:16:@14951.4]
  assign _T_17353 = 6'h2a == _T_11317_61; // @[Mux.scala 46:19:@14952.4]
  assign _T_17354 = _T_17353 ? _T_10366_41 : _T_17352; // @[Mux.scala 46:16:@14953.4]
  assign _T_17355 = 6'h29 == _T_11317_61; // @[Mux.scala 46:19:@14954.4]
  assign _T_17356 = _T_17355 ? _T_10366_40 : _T_17354; // @[Mux.scala 46:16:@14955.4]
  assign _T_17357 = 6'h28 == _T_11317_61; // @[Mux.scala 46:19:@14956.4]
  assign _T_17358 = _T_17357 ? _T_10366_39 : _T_17356; // @[Mux.scala 46:16:@14957.4]
  assign _T_17359 = 6'h27 == _T_11317_61; // @[Mux.scala 46:19:@14958.4]
  assign _T_17360 = _T_17359 ? _T_10366_38 : _T_17358; // @[Mux.scala 46:16:@14959.4]
  assign _T_17361 = 6'h26 == _T_11317_61; // @[Mux.scala 46:19:@14960.4]
  assign _T_17362 = _T_17361 ? _T_10366_37 : _T_17360; // @[Mux.scala 46:16:@14961.4]
  assign _T_17363 = 6'h25 == _T_11317_61; // @[Mux.scala 46:19:@14962.4]
  assign _T_17364 = _T_17363 ? _T_10366_36 : _T_17362; // @[Mux.scala 46:16:@14963.4]
  assign _T_17365 = 6'h24 == _T_11317_61; // @[Mux.scala 46:19:@14964.4]
  assign _T_17366 = _T_17365 ? _T_10366_35 : _T_17364; // @[Mux.scala 46:16:@14965.4]
  assign _T_17367 = 6'h23 == _T_11317_61; // @[Mux.scala 46:19:@14966.4]
  assign _T_17368 = _T_17367 ? _T_10366_34 : _T_17366; // @[Mux.scala 46:16:@14967.4]
  assign _T_17369 = 6'h22 == _T_11317_61; // @[Mux.scala 46:19:@14968.4]
  assign _T_17370 = _T_17369 ? _T_10366_33 : _T_17368; // @[Mux.scala 46:16:@14969.4]
  assign _T_17371 = 6'h21 == _T_11317_61; // @[Mux.scala 46:19:@14970.4]
  assign _T_17372 = _T_17371 ? _T_10366_32 : _T_17370; // @[Mux.scala 46:16:@14971.4]
  assign _T_17373 = 6'h20 == _T_11317_61; // @[Mux.scala 46:19:@14972.4]
  assign _T_17374 = _T_17373 ? _T_10366_31 : _T_17372; // @[Mux.scala 46:16:@14973.4]
  assign _T_17375 = 6'h1f == _T_11317_61; // @[Mux.scala 46:19:@14974.4]
  assign _T_17376 = _T_17375 ? _T_10366_30 : _T_17374; // @[Mux.scala 46:16:@14975.4]
  assign _T_17377 = 6'h1e == _T_11317_61; // @[Mux.scala 46:19:@14976.4]
  assign _T_17378 = _T_17377 ? _T_10366_29 : _T_17376; // @[Mux.scala 46:16:@14977.4]
  assign _T_17379 = 6'h1d == _T_11317_61; // @[Mux.scala 46:19:@14978.4]
  assign _T_17380 = _T_17379 ? _T_10366_28 : _T_17378; // @[Mux.scala 46:16:@14979.4]
  assign _T_17381 = 6'h1c == _T_11317_61; // @[Mux.scala 46:19:@14980.4]
  assign _T_17382 = _T_17381 ? _T_10366_27 : _T_17380; // @[Mux.scala 46:16:@14981.4]
  assign _T_17383 = 6'h1b == _T_11317_61; // @[Mux.scala 46:19:@14982.4]
  assign _T_17384 = _T_17383 ? _T_10366_26 : _T_17382; // @[Mux.scala 46:16:@14983.4]
  assign _T_17385 = 6'h1a == _T_11317_61; // @[Mux.scala 46:19:@14984.4]
  assign _T_17386 = _T_17385 ? _T_10366_25 : _T_17384; // @[Mux.scala 46:16:@14985.4]
  assign _T_17387 = 6'h19 == _T_11317_61; // @[Mux.scala 46:19:@14986.4]
  assign _T_17388 = _T_17387 ? _T_10366_24 : _T_17386; // @[Mux.scala 46:16:@14987.4]
  assign _T_17389 = 6'h18 == _T_11317_61; // @[Mux.scala 46:19:@14988.4]
  assign _T_17390 = _T_17389 ? _T_10366_23 : _T_17388; // @[Mux.scala 46:16:@14989.4]
  assign _T_17391 = 6'h17 == _T_11317_61; // @[Mux.scala 46:19:@14990.4]
  assign _T_17392 = _T_17391 ? _T_10366_22 : _T_17390; // @[Mux.scala 46:16:@14991.4]
  assign _T_17393 = 6'h16 == _T_11317_61; // @[Mux.scala 46:19:@14992.4]
  assign _T_17394 = _T_17393 ? _T_10366_21 : _T_17392; // @[Mux.scala 46:16:@14993.4]
  assign _T_17395 = 6'h15 == _T_11317_61; // @[Mux.scala 46:19:@14994.4]
  assign _T_17396 = _T_17395 ? _T_10366_20 : _T_17394; // @[Mux.scala 46:16:@14995.4]
  assign _T_17397 = 6'h14 == _T_11317_61; // @[Mux.scala 46:19:@14996.4]
  assign _T_17398 = _T_17397 ? _T_10366_19 : _T_17396; // @[Mux.scala 46:16:@14997.4]
  assign _T_17399 = 6'h13 == _T_11317_61; // @[Mux.scala 46:19:@14998.4]
  assign _T_17400 = _T_17399 ? _T_10366_18 : _T_17398; // @[Mux.scala 46:16:@14999.4]
  assign _T_17401 = 6'h12 == _T_11317_61; // @[Mux.scala 46:19:@15000.4]
  assign _T_17402 = _T_17401 ? _T_10366_17 : _T_17400; // @[Mux.scala 46:16:@15001.4]
  assign _T_17403 = 6'h11 == _T_11317_61; // @[Mux.scala 46:19:@15002.4]
  assign _T_17404 = _T_17403 ? _T_10366_16 : _T_17402; // @[Mux.scala 46:16:@15003.4]
  assign _T_17405 = 6'h10 == _T_11317_61; // @[Mux.scala 46:19:@15004.4]
  assign _T_17406 = _T_17405 ? _T_10366_15 : _T_17404; // @[Mux.scala 46:16:@15005.4]
  assign _T_17407 = 6'hf == _T_11317_61; // @[Mux.scala 46:19:@15006.4]
  assign _T_17408 = _T_17407 ? _T_10366_14 : _T_17406; // @[Mux.scala 46:16:@15007.4]
  assign _T_17409 = 6'he == _T_11317_61; // @[Mux.scala 46:19:@15008.4]
  assign _T_17410 = _T_17409 ? _T_10366_13 : _T_17408; // @[Mux.scala 46:16:@15009.4]
  assign _T_17411 = 6'hd == _T_11317_61; // @[Mux.scala 46:19:@15010.4]
  assign _T_17412 = _T_17411 ? _T_10366_12 : _T_17410; // @[Mux.scala 46:16:@15011.4]
  assign _T_17413 = 6'hc == _T_11317_61; // @[Mux.scala 46:19:@15012.4]
  assign _T_17414 = _T_17413 ? _T_10366_11 : _T_17412; // @[Mux.scala 46:16:@15013.4]
  assign _T_17415 = 6'hb == _T_11317_61; // @[Mux.scala 46:19:@15014.4]
  assign _T_17416 = _T_17415 ? _T_10366_10 : _T_17414; // @[Mux.scala 46:16:@15015.4]
  assign _T_17417 = 6'ha == _T_11317_61; // @[Mux.scala 46:19:@15016.4]
  assign _T_17418 = _T_17417 ? _T_10366_9 : _T_17416; // @[Mux.scala 46:16:@15017.4]
  assign _T_17419 = 6'h9 == _T_11317_61; // @[Mux.scala 46:19:@15018.4]
  assign _T_17420 = _T_17419 ? _T_10366_8 : _T_17418; // @[Mux.scala 46:16:@15019.4]
  assign _T_17421 = 6'h8 == _T_11317_61; // @[Mux.scala 46:19:@15020.4]
  assign _T_17422 = _T_17421 ? _T_10366_7 : _T_17420; // @[Mux.scala 46:16:@15021.4]
  assign _T_17423 = 6'h7 == _T_11317_61; // @[Mux.scala 46:19:@15022.4]
  assign _T_17424 = _T_17423 ? _T_10366_6 : _T_17422; // @[Mux.scala 46:16:@15023.4]
  assign _T_17425 = 6'h6 == _T_11317_61; // @[Mux.scala 46:19:@15024.4]
  assign _T_17426 = _T_17425 ? _T_10366_5 : _T_17424; // @[Mux.scala 46:16:@15025.4]
  assign _T_17427 = 6'h5 == _T_11317_61; // @[Mux.scala 46:19:@15026.4]
  assign _T_17428 = _T_17427 ? _T_10366_4 : _T_17426; // @[Mux.scala 46:16:@15027.4]
  assign _T_17429 = 6'h4 == _T_11317_61; // @[Mux.scala 46:19:@15028.4]
  assign _T_17430 = _T_17429 ? _T_10366_3 : _T_17428; // @[Mux.scala 46:16:@15029.4]
  assign _T_17431 = 6'h3 == _T_11317_61; // @[Mux.scala 46:19:@15030.4]
  assign _T_17432 = _T_17431 ? _T_10366_2 : _T_17430; // @[Mux.scala 46:16:@15031.4]
  assign _T_17433 = 6'h2 == _T_11317_61; // @[Mux.scala 46:19:@15032.4]
  assign _T_17434 = _T_17433 ? _T_10366_1 : _T_17432; // @[Mux.scala 46:16:@15033.4]
  assign _T_17435 = 6'h1 == _T_11317_61; // @[Mux.scala 46:19:@15034.4]
  assign _T_17436 = _T_17435 ? _T_10366_0 : _T_17434; // @[Mux.scala 46:16:@15035.4]
  assign _T_17501 = 6'h3f == _T_11317_62; // @[Mux.scala 46:19:@15037.4]
  assign _T_17502 = _T_17501 ? _T_10366_62 : 8'h0; // @[Mux.scala 46:16:@15038.4]
  assign _T_17503 = 6'h3e == _T_11317_62; // @[Mux.scala 46:19:@15039.4]
  assign _T_17504 = _T_17503 ? _T_10366_61 : _T_17502; // @[Mux.scala 46:16:@15040.4]
  assign _T_17505 = 6'h3d == _T_11317_62; // @[Mux.scala 46:19:@15041.4]
  assign _T_17506 = _T_17505 ? _T_10366_60 : _T_17504; // @[Mux.scala 46:16:@15042.4]
  assign _T_17507 = 6'h3c == _T_11317_62; // @[Mux.scala 46:19:@15043.4]
  assign _T_17508 = _T_17507 ? _T_10366_59 : _T_17506; // @[Mux.scala 46:16:@15044.4]
  assign _T_17509 = 6'h3b == _T_11317_62; // @[Mux.scala 46:19:@15045.4]
  assign _T_17510 = _T_17509 ? _T_10366_58 : _T_17508; // @[Mux.scala 46:16:@15046.4]
  assign _T_17511 = 6'h3a == _T_11317_62; // @[Mux.scala 46:19:@15047.4]
  assign _T_17512 = _T_17511 ? _T_10366_57 : _T_17510; // @[Mux.scala 46:16:@15048.4]
  assign _T_17513 = 6'h39 == _T_11317_62; // @[Mux.scala 46:19:@15049.4]
  assign _T_17514 = _T_17513 ? _T_10366_56 : _T_17512; // @[Mux.scala 46:16:@15050.4]
  assign _T_17515 = 6'h38 == _T_11317_62; // @[Mux.scala 46:19:@15051.4]
  assign _T_17516 = _T_17515 ? _T_10366_55 : _T_17514; // @[Mux.scala 46:16:@15052.4]
  assign _T_17517 = 6'h37 == _T_11317_62; // @[Mux.scala 46:19:@15053.4]
  assign _T_17518 = _T_17517 ? _T_10366_54 : _T_17516; // @[Mux.scala 46:16:@15054.4]
  assign _T_17519 = 6'h36 == _T_11317_62; // @[Mux.scala 46:19:@15055.4]
  assign _T_17520 = _T_17519 ? _T_10366_53 : _T_17518; // @[Mux.scala 46:16:@15056.4]
  assign _T_17521 = 6'h35 == _T_11317_62; // @[Mux.scala 46:19:@15057.4]
  assign _T_17522 = _T_17521 ? _T_10366_52 : _T_17520; // @[Mux.scala 46:16:@15058.4]
  assign _T_17523 = 6'h34 == _T_11317_62; // @[Mux.scala 46:19:@15059.4]
  assign _T_17524 = _T_17523 ? _T_10366_51 : _T_17522; // @[Mux.scala 46:16:@15060.4]
  assign _T_17525 = 6'h33 == _T_11317_62; // @[Mux.scala 46:19:@15061.4]
  assign _T_17526 = _T_17525 ? _T_10366_50 : _T_17524; // @[Mux.scala 46:16:@15062.4]
  assign _T_17527 = 6'h32 == _T_11317_62; // @[Mux.scala 46:19:@15063.4]
  assign _T_17528 = _T_17527 ? _T_10366_49 : _T_17526; // @[Mux.scala 46:16:@15064.4]
  assign _T_17529 = 6'h31 == _T_11317_62; // @[Mux.scala 46:19:@15065.4]
  assign _T_17530 = _T_17529 ? _T_10366_48 : _T_17528; // @[Mux.scala 46:16:@15066.4]
  assign _T_17531 = 6'h30 == _T_11317_62; // @[Mux.scala 46:19:@15067.4]
  assign _T_17532 = _T_17531 ? _T_10366_47 : _T_17530; // @[Mux.scala 46:16:@15068.4]
  assign _T_17533 = 6'h2f == _T_11317_62; // @[Mux.scala 46:19:@15069.4]
  assign _T_17534 = _T_17533 ? _T_10366_46 : _T_17532; // @[Mux.scala 46:16:@15070.4]
  assign _T_17535 = 6'h2e == _T_11317_62; // @[Mux.scala 46:19:@15071.4]
  assign _T_17536 = _T_17535 ? _T_10366_45 : _T_17534; // @[Mux.scala 46:16:@15072.4]
  assign _T_17537 = 6'h2d == _T_11317_62; // @[Mux.scala 46:19:@15073.4]
  assign _T_17538 = _T_17537 ? _T_10366_44 : _T_17536; // @[Mux.scala 46:16:@15074.4]
  assign _T_17539 = 6'h2c == _T_11317_62; // @[Mux.scala 46:19:@15075.4]
  assign _T_17540 = _T_17539 ? _T_10366_43 : _T_17538; // @[Mux.scala 46:16:@15076.4]
  assign _T_17541 = 6'h2b == _T_11317_62; // @[Mux.scala 46:19:@15077.4]
  assign _T_17542 = _T_17541 ? _T_10366_42 : _T_17540; // @[Mux.scala 46:16:@15078.4]
  assign _T_17543 = 6'h2a == _T_11317_62; // @[Mux.scala 46:19:@15079.4]
  assign _T_17544 = _T_17543 ? _T_10366_41 : _T_17542; // @[Mux.scala 46:16:@15080.4]
  assign _T_17545 = 6'h29 == _T_11317_62; // @[Mux.scala 46:19:@15081.4]
  assign _T_17546 = _T_17545 ? _T_10366_40 : _T_17544; // @[Mux.scala 46:16:@15082.4]
  assign _T_17547 = 6'h28 == _T_11317_62; // @[Mux.scala 46:19:@15083.4]
  assign _T_17548 = _T_17547 ? _T_10366_39 : _T_17546; // @[Mux.scala 46:16:@15084.4]
  assign _T_17549 = 6'h27 == _T_11317_62; // @[Mux.scala 46:19:@15085.4]
  assign _T_17550 = _T_17549 ? _T_10366_38 : _T_17548; // @[Mux.scala 46:16:@15086.4]
  assign _T_17551 = 6'h26 == _T_11317_62; // @[Mux.scala 46:19:@15087.4]
  assign _T_17552 = _T_17551 ? _T_10366_37 : _T_17550; // @[Mux.scala 46:16:@15088.4]
  assign _T_17553 = 6'h25 == _T_11317_62; // @[Mux.scala 46:19:@15089.4]
  assign _T_17554 = _T_17553 ? _T_10366_36 : _T_17552; // @[Mux.scala 46:16:@15090.4]
  assign _T_17555 = 6'h24 == _T_11317_62; // @[Mux.scala 46:19:@15091.4]
  assign _T_17556 = _T_17555 ? _T_10366_35 : _T_17554; // @[Mux.scala 46:16:@15092.4]
  assign _T_17557 = 6'h23 == _T_11317_62; // @[Mux.scala 46:19:@15093.4]
  assign _T_17558 = _T_17557 ? _T_10366_34 : _T_17556; // @[Mux.scala 46:16:@15094.4]
  assign _T_17559 = 6'h22 == _T_11317_62; // @[Mux.scala 46:19:@15095.4]
  assign _T_17560 = _T_17559 ? _T_10366_33 : _T_17558; // @[Mux.scala 46:16:@15096.4]
  assign _T_17561 = 6'h21 == _T_11317_62; // @[Mux.scala 46:19:@15097.4]
  assign _T_17562 = _T_17561 ? _T_10366_32 : _T_17560; // @[Mux.scala 46:16:@15098.4]
  assign _T_17563 = 6'h20 == _T_11317_62; // @[Mux.scala 46:19:@15099.4]
  assign _T_17564 = _T_17563 ? _T_10366_31 : _T_17562; // @[Mux.scala 46:16:@15100.4]
  assign _T_17565 = 6'h1f == _T_11317_62; // @[Mux.scala 46:19:@15101.4]
  assign _T_17566 = _T_17565 ? _T_10366_30 : _T_17564; // @[Mux.scala 46:16:@15102.4]
  assign _T_17567 = 6'h1e == _T_11317_62; // @[Mux.scala 46:19:@15103.4]
  assign _T_17568 = _T_17567 ? _T_10366_29 : _T_17566; // @[Mux.scala 46:16:@15104.4]
  assign _T_17569 = 6'h1d == _T_11317_62; // @[Mux.scala 46:19:@15105.4]
  assign _T_17570 = _T_17569 ? _T_10366_28 : _T_17568; // @[Mux.scala 46:16:@15106.4]
  assign _T_17571 = 6'h1c == _T_11317_62; // @[Mux.scala 46:19:@15107.4]
  assign _T_17572 = _T_17571 ? _T_10366_27 : _T_17570; // @[Mux.scala 46:16:@15108.4]
  assign _T_17573 = 6'h1b == _T_11317_62; // @[Mux.scala 46:19:@15109.4]
  assign _T_17574 = _T_17573 ? _T_10366_26 : _T_17572; // @[Mux.scala 46:16:@15110.4]
  assign _T_17575 = 6'h1a == _T_11317_62; // @[Mux.scala 46:19:@15111.4]
  assign _T_17576 = _T_17575 ? _T_10366_25 : _T_17574; // @[Mux.scala 46:16:@15112.4]
  assign _T_17577 = 6'h19 == _T_11317_62; // @[Mux.scala 46:19:@15113.4]
  assign _T_17578 = _T_17577 ? _T_10366_24 : _T_17576; // @[Mux.scala 46:16:@15114.4]
  assign _T_17579 = 6'h18 == _T_11317_62; // @[Mux.scala 46:19:@15115.4]
  assign _T_17580 = _T_17579 ? _T_10366_23 : _T_17578; // @[Mux.scala 46:16:@15116.4]
  assign _T_17581 = 6'h17 == _T_11317_62; // @[Mux.scala 46:19:@15117.4]
  assign _T_17582 = _T_17581 ? _T_10366_22 : _T_17580; // @[Mux.scala 46:16:@15118.4]
  assign _T_17583 = 6'h16 == _T_11317_62; // @[Mux.scala 46:19:@15119.4]
  assign _T_17584 = _T_17583 ? _T_10366_21 : _T_17582; // @[Mux.scala 46:16:@15120.4]
  assign _T_17585 = 6'h15 == _T_11317_62; // @[Mux.scala 46:19:@15121.4]
  assign _T_17586 = _T_17585 ? _T_10366_20 : _T_17584; // @[Mux.scala 46:16:@15122.4]
  assign _T_17587 = 6'h14 == _T_11317_62; // @[Mux.scala 46:19:@15123.4]
  assign _T_17588 = _T_17587 ? _T_10366_19 : _T_17586; // @[Mux.scala 46:16:@15124.4]
  assign _T_17589 = 6'h13 == _T_11317_62; // @[Mux.scala 46:19:@15125.4]
  assign _T_17590 = _T_17589 ? _T_10366_18 : _T_17588; // @[Mux.scala 46:16:@15126.4]
  assign _T_17591 = 6'h12 == _T_11317_62; // @[Mux.scala 46:19:@15127.4]
  assign _T_17592 = _T_17591 ? _T_10366_17 : _T_17590; // @[Mux.scala 46:16:@15128.4]
  assign _T_17593 = 6'h11 == _T_11317_62; // @[Mux.scala 46:19:@15129.4]
  assign _T_17594 = _T_17593 ? _T_10366_16 : _T_17592; // @[Mux.scala 46:16:@15130.4]
  assign _T_17595 = 6'h10 == _T_11317_62; // @[Mux.scala 46:19:@15131.4]
  assign _T_17596 = _T_17595 ? _T_10366_15 : _T_17594; // @[Mux.scala 46:16:@15132.4]
  assign _T_17597 = 6'hf == _T_11317_62; // @[Mux.scala 46:19:@15133.4]
  assign _T_17598 = _T_17597 ? _T_10366_14 : _T_17596; // @[Mux.scala 46:16:@15134.4]
  assign _T_17599 = 6'he == _T_11317_62; // @[Mux.scala 46:19:@15135.4]
  assign _T_17600 = _T_17599 ? _T_10366_13 : _T_17598; // @[Mux.scala 46:16:@15136.4]
  assign _T_17601 = 6'hd == _T_11317_62; // @[Mux.scala 46:19:@15137.4]
  assign _T_17602 = _T_17601 ? _T_10366_12 : _T_17600; // @[Mux.scala 46:16:@15138.4]
  assign _T_17603 = 6'hc == _T_11317_62; // @[Mux.scala 46:19:@15139.4]
  assign _T_17604 = _T_17603 ? _T_10366_11 : _T_17602; // @[Mux.scala 46:16:@15140.4]
  assign _T_17605 = 6'hb == _T_11317_62; // @[Mux.scala 46:19:@15141.4]
  assign _T_17606 = _T_17605 ? _T_10366_10 : _T_17604; // @[Mux.scala 46:16:@15142.4]
  assign _T_17607 = 6'ha == _T_11317_62; // @[Mux.scala 46:19:@15143.4]
  assign _T_17608 = _T_17607 ? _T_10366_9 : _T_17606; // @[Mux.scala 46:16:@15144.4]
  assign _T_17609 = 6'h9 == _T_11317_62; // @[Mux.scala 46:19:@15145.4]
  assign _T_17610 = _T_17609 ? _T_10366_8 : _T_17608; // @[Mux.scala 46:16:@15146.4]
  assign _T_17611 = 6'h8 == _T_11317_62; // @[Mux.scala 46:19:@15147.4]
  assign _T_17612 = _T_17611 ? _T_10366_7 : _T_17610; // @[Mux.scala 46:16:@15148.4]
  assign _T_17613 = 6'h7 == _T_11317_62; // @[Mux.scala 46:19:@15149.4]
  assign _T_17614 = _T_17613 ? _T_10366_6 : _T_17612; // @[Mux.scala 46:16:@15150.4]
  assign _T_17615 = 6'h6 == _T_11317_62; // @[Mux.scala 46:19:@15151.4]
  assign _T_17616 = _T_17615 ? _T_10366_5 : _T_17614; // @[Mux.scala 46:16:@15152.4]
  assign _T_17617 = 6'h5 == _T_11317_62; // @[Mux.scala 46:19:@15153.4]
  assign _T_17618 = _T_17617 ? _T_10366_4 : _T_17616; // @[Mux.scala 46:16:@15154.4]
  assign _T_17619 = 6'h4 == _T_11317_62; // @[Mux.scala 46:19:@15155.4]
  assign _T_17620 = _T_17619 ? _T_10366_3 : _T_17618; // @[Mux.scala 46:16:@15156.4]
  assign _T_17621 = 6'h3 == _T_11317_62; // @[Mux.scala 46:19:@15157.4]
  assign _T_17622 = _T_17621 ? _T_10366_2 : _T_17620; // @[Mux.scala 46:16:@15158.4]
  assign _T_17623 = 6'h2 == _T_11317_62; // @[Mux.scala 46:19:@15159.4]
  assign _T_17624 = _T_17623 ? _T_10366_1 : _T_17622; // @[Mux.scala 46:16:@15160.4]
  assign _T_17625 = 6'h1 == _T_11317_62; // @[Mux.scala 46:19:@15161.4]
  assign _T_17626 = _T_17625 ? _T_10366_0 : _T_17624; // @[Mux.scala 46:16:@15162.4]
  assign _T_17692 = 7'h40 == _T_11317_63; // @[Mux.scala 46:19:@15164.4]
  assign _T_17693 = _T_17692 ? _T_10366_63 : 8'h0; // @[Mux.scala 46:16:@15165.4]
  assign _T_17694 = 7'h3f == _T_11317_63; // @[Mux.scala 46:19:@15166.4]
  assign _T_17695 = _T_17694 ? _T_10366_62 : _T_17693; // @[Mux.scala 46:16:@15167.4]
  assign _T_17696 = 7'h3e == _T_11317_63; // @[Mux.scala 46:19:@15168.4]
  assign _T_17697 = _T_17696 ? _T_10366_61 : _T_17695; // @[Mux.scala 46:16:@15169.4]
  assign _T_17698 = 7'h3d == _T_11317_63; // @[Mux.scala 46:19:@15170.4]
  assign _T_17699 = _T_17698 ? _T_10366_60 : _T_17697; // @[Mux.scala 46:16:@15171.4]
  assign _T_17700 = 7'h3c == _T_11317_63; // @[Mux.scala 46:19:@15172.4]
  assign _T_17701 = _T_17700 ? _T_10366_59 : _T_17699; // @[Mux.scala 46:16:@15173.4]
  assign _T_17702 = 7'h3b == _T_11317_63; // @[Mux.scala 46:19:@15174.4]
  assign _T_17703 = _T_17702 ? _T_10366_58 : _T_17701; // @[Mux.scala 46:16:@15175.4]
  assign _T_17704 = 7'h3a == _T_11317_63; // @[Mux.scala 46:19:@15176.4]
  assign _T_17705 = _T_17704 ? _T_10366_57 : _T_17703; // @[Mux.scala 46:16:@15177.4]
  assign _T_17706 = 7'h39 == _T_11317_63; // @[Mux.scala 46:19:@15178.4]
  assign _T_17707 = _T_17706 ? _T_10366_56 : _T_17705; // @[Mux.scala 46:16:@15179.4]
  assign _T_17708 = 7'h38 == _T_11317_63; // @[Mux.scala 46:19:@15180.4]
  assign _T_17709 = _T_17708 ? _T_10366_55 : _T_17707; // @[Mux.scala 46:16:@15181.4]
  assign _T_17710 = 7'h37 == _T_11317_63; // @[Mux.scala 46:19:@15182.4]
  assign _T_17711 = _T_17710 ? _T_10366_54 : _T_17709; // @[Mux.scala 46:16:@15183.4]
  assign _T_17712 = 7'h36 == _T_11317_63; // @[Mux.scala 46:19:@15184.4]
  assign _T_17713 = _T_17712 ? _T_10366_53 : _T_17711; // @[Mux.scala 46:16:@15185.4]
  assign _T_17714 = 7'h35 == _T_11317_63; // @[Mux.scala 46:19:@15186.4]
  assign _T_17715 = _T_17714 ? _T_10366_52 : _T_17713; // @[Mux.scala 46:16:@15187.4]
  assign _T_17716 = 7'h34 == _T_11317_63; // @[Mux.scala 46:19:@15188.4]
  assign _T_17717 = _T_17716 ? _T_10366_51 : _T_17715; // @[Mux.scala 46:16:@15189.4]
  assign _T_17718 = 7'h33 == _T_11317_63; // @[Mux.scala 46:19:@15190.4]
  assign _T_17719 = _T_17718 ? _T_10366_50 : _T_17717; // @[Mux.scala 46:16:@15191.4]
  assign _T_17720 = 7'h32 == _T_11317_63; // @[Mux.scala 46:19:@15192.4]
  assign _T_17721 = _T_17720 ? _T_10366_49 : _T_17719; // @[Mux.scala 46:16:@15193.4]
  assign _T_17722 = 7'h31 == _T_11317_63; // @[Mux.scala 46:19:@15194.4]
  assign _T_17723 = _T_17722 ? _T_10366_48 : _T_17721; // @[Mux.scala 46:16:@15195.4]
  assign _T_17724 = 7'h30 == _T_11317_63; // @[Mux.scala 46:19:@15196.4]
  assign _T_17725 = _T_17724 ? _T_10366_47 : _T_17723; // @[Mux.scala 46:16:@15197.4]
  assign _T_17726 = 7'h2f == _T_11317_63; // @[Mux.scala 46:19:@15198.4]
  assign _T_17727 = _T_17726 ? _T_10366_46 : _T_17725; // @[Mux.scala 46:16:@15199.4]
  assign _T_17728 = 7'h2e == _T_11317_63; // @[Mux.scala 46:19:@15200.4]
  assign _T_17729 = _T_17728 ? _T_10366_45 : _T_17727; // @[Mux.scala 46:16:@15201.4]
  assign _T_17730 = 7'h2d == _T_11317_63; // @[Mux.scala 46:19:@15202.4]
  assign _T_17731 = _T_17730 ? _T_10366_44 : _T_17729; // @[Mux.scala 46:16:@15203.4]
  assign _T_17732 = 7'h2c == _T_11317_63; // @[Mux.scala 46:19:@15204.4]
  assign _T_17733 = _T_17732 ? _T_10366_43 : _T_17731; // @[Mux.scala 46:16:@15205.4]
  assign _T_17734 = 7'h2b == _T_11317_63; // @[Mux.scala 46:19:@15206.4]
  assign _T_17735 = _T_17734 ? _T_10366_42 : _T_17733; // @[Mux.scala 46:16:@15207.4]
  assign _T_17736 = 7'h2a == _T_11317_63; // @[Mux.scala 46:19:@15208.4]
  assign _T_17737 = _T_17736 ? _T_10366_41 : _T_17735; // @[Mux.scala 46:16:@15209.4]
  assign _T_17738 = 7'h29 == _T_11317_63; // @[Mux.scala 46:19:@15210.4]
  assign _T_17739 = _T_17738 ? _T_10366_40 : _T_17737; // @[Mux.scala 46:16:@15211.4]
  assign _T_17740 = 7'h28 == _T_11317_63; // @[Mux.scala 46:19:@15212.4]
  assign _T_17741 = _T_17740 ? _T_10366_39 : _T_17739; // @[Mux.scala 46:16:@15213.4]
  assign _T_17742 = 7'h27 == _T_11317_63; // @[Mux.scala 46:19:@15214.4]
  assign _T_17743 = _T_17742 ? _T_10366_38 : _T_17741; // @[Mux.scala 46:16:@15215.4]
  assign _T_17744 = 7'h26 == _T_11317_63; // @[Mux.scala 46:19:@15216.4]
  assign _T_17745 = _T_17744 ? _T_10366_37 : _T_17743; // @[Mux.scala 46:16:@15217.4]
  assign _T_17746 = 7'h25 == _T_11317_63; // @[Mux.scala 46:19:@15218.4]
  assign _T_17747 = _T_17746 ? _T_10366_36 : _T_17745; // @[Mux.scala 46:16:@15219.4]
  assign _T_17748 = 7'h24 == _T_11317_63; // @[Mux.scala 46:19:@15220.4]
  assign _T_17749 = _T_17748 ? _T_10366_35 : _T_17747; // @[Mux.scala 46:16:@15221.4]
  assign _T_17750 = 7'h23 == _T_11317_63; // @[Mux.scala 46:19:@15222.4]
  assign _T_17751 = _T_17750 ? _T_10366_34 : _T_17749; // @[Mux.scala 46:16:@15223.4]
  assign _T_17752 = 7'h22 == _T_11317_63; // @[Mux.scala 46:19:@15224.4]
  assign _T_17753 = _T_17752 ? _T_10366_33 : _T_17751; // @[Mux.scala 46:16:@15225.4]
  assign _T_17754 = 7'h21 == _T_11317_63; // @[Mux.scala 46:19:@15226.4]
  assign _T_17755 = _T_17754 ? _T_10366_32 : _T_17753; // @[Mux.scala 46:16:@15227.4]
  assign _T_17756 = 7'h20 == _T_11317_63; // @[Mux.scala 46:19:@15228.4]
  assign _T_17757 = _T_17756 ? _T_10366_31 : _T_17755; // @[Mux.scala 46:16:@15229.4]
  assign _T_17758 = 7'h1f == _T_11317_63; // @[Mux.scala 46:19:@15230.4]
  assign _T_17759 = _T_17758 ? _T_10366_30 : _T_17757; // @[Mux.scala 46:16:@15231.4]
  assign _T_17760 = 7'h1e == _T_11317_63; // @[Mux.scala 46:19:@15232.4]
  assign _T_17761 = _T_17760 ? _T_10366_29 : _T_17759; // @[Mux.scala 46:16:@15233.4]
  assign _T_17762 = 7'h1d == _T_11317_63; // @[Mux.scala 46:19:@15234.4]
  assign _T_17763 = _T_17762 ? _T_10366_28 : _T_17761; // @[Mux.scala 46:16:@15235.4]
  assign _T_17764 = 7'h1c == _T_11317_63; // @[Mux.scala 46:19:@15236.4]
  assign _T_17765 = _T_17764 ? _T_10366_27 : _T_17763; // @[Mux.scala 46:16:@15237.4]
  assign _T_17766 = 7'h1b == _T_11317_63; // @[Mux.scala 46:19:@15238.4]
  assign _T_17767 = _T_17766 ? _T_10366_26 : _T_17765; // @[Mux.scala 46:16:@15239.4]
  assign _T_17768 = 7'h1a == _T_11317_63; // @[Mux.scala 46:19:@15240.4]
  assign _T_17769 = _T_17768 ? _T_10366_25 : _T_17767; // @[Mux.scala 46:16:@15241.4]
  assign _T_17770 = 7'h19 == _T_11317_63; // @[Mux.scala 46:19:@15242.4]
  assign _T_17771 = _T_17770 ? _T_10366_24 : _T_17769; // @[Mux.scala 46:16:@15243.4]
  assign _T_17772 = 7'h18 == _T_11317_63; // @[Mux.scala 46:19:@15244.4]
  assign _T_17773 = _T_17772 ? _T_10366_23 : _T_17771; // @[Mux.scala 46:16:@15245.4]
  assign _T_17774 = 7'h17 == _T_11317_63; // @[Mux.scala 46:19:@15246.4]
  assign _T_17775 = _T_17774 ? _T_10366_22 : _T_17773; // @[Mux.scala 46:16:@15247.4]
  assign _T_17776 = 7'h16 == _T_11317_63; // @[Mux.scala 46:19:@15248.4]
  assign _T_17777 = _T_17776 ? _T_10366_21 : _T_17775; // @[Mux.scala 46:16:@15249.4]
  assign _T_17778 = 7'h15 == _T_11317_63; // @[Mux.scala 46:19:@15250.4]
  assign _T_17779 = _T_17778 ? _T_10366_20 : _T_17777; // @[Mux.scala 46:16:@15251.4]
  assign _T_17780 = 7'h14 == _T_11317_63; // @[Mux.scala 46:19:@15252.4]
  assign _T_17781 = _T_17780 ? _T_10366_19 : _T_17779; // @[Mux.scala 46:16:@15253.4]
  assign _T_17782 = 7'h13 == _T_11317_63; // @[Mux.scala 46:19:@15254.4]
  assign _T_17783 = _T_17782 ? _T_10366_18 : _T_17781; // @[Mux.scala 46:16:@15255.4]
  assign _T_17784 = 7'h12 == _T_11317_63; // @[Mux.scala 46:19:@15256.4]
  assign _T_17785 = _T_17784 ? _T_10366_17 : _T_17783; // @[Mux.scala 46:16:@15257.4]
  assign _T_17786 = 7'h11 == _T_11317_63; // @[Mux.scala 46:19:@15258.4]
  assign _T_17787 = _T_17786 ? _T_10366_16 : _T_17785; // @[Mux.scala 46:16:@15259.4]
  assign _T_17788 = 7'h10 == _T_11317_63; // @[Mux.scala 46:19:@15260.4]
  assign _T_17789 = _T_17788 ? _T_10366_15 : _T_17787; // @[Mux.scala 46:16:@15261.4]
  assign _T_17790 = 7'hf == _T_11317_63; // @[Mux.scala 46:19:@15262.4]
  assign _T_17791 = _T_17790 ? _T_10366_14 : _T_17789; // @[Mux.scala 46:16:@15263.4]
  assign _T_17792 = 7'he == _T_11317_63; // @[Mux.scala 46:19:@15264.4]
  assign _T_17793 = _T_17792 ? _T_10366_13 : _T_17791; // @[Mux.scala 46:16:@15265.4]
  assign _T_17794 = 7'hd == _T_11317_63; // @[Mux.scala 46:19:@15266.4]
  assign _T_17795 = _T_17794 ? _T_10366_12 : _T_17793; // @[Mux.scala 46:16:@15267.4]
  assign _T_17796 = 7'hc == _T_11317_63; // @[Mux.scala 46:19:@15268.4]
  assign _T_17797 = _T_17796 ? _T_10366_11 : _T_17795; // @[Mux.scala 46:16:@15269.4]
  assign _T_17798 = 7'hb == _T_11317_63; // @[Mux.scala 46:19:@15270.4]
  assign _T_17799 = _T_17798 ? _T_10366_10 : _T_17797; // @[Mux.scala 46:16:@15271.4]
  assign _T_17800 = 7'ha == _T_11317_63; // @[Mux.scala 46:19:@15272.4]
  assign _T_17801 = _T_17800 ? _T_10366_9 : _T_17799; // @[Mux.scala 46:16:@15273.4]
  assign _T_17802 = 7'h9 == _T_11317_63; // @[Mux.scala 46:19:@15274.4]
  assign _T_17803 = _T_17802 ? _T_10366_8 : _T_17801; // @[Mux.scala 46:16:@15275.4]
  assign _T_17804 = 7'h8 == _T_11317_63; // @[Mux.scala 46:19:@15276.4]
  assign _T_17805 = _T_17804 ? _T_10366_7 : _T_17803; // @[Mux.scala 46:16:@15277.4]
  assign _T_17806 = 7'h7 == _T_11317_63; // @[Mux.scala 46:19:@15278.4]
  assign _T_17807 = _T_17806 ? _T_10366_6 : _T_17805; // @[Mux.scala 46:16:@15279.4]
  assign _T_17808 = 7'h6 == _T_11317_63; // @[Mux.scala 46:19:@15280.4]
  assign _T_17809 = _T_17808 ? _T_10366_5 : _T_17807; // @[Mux.scala 46:16:@15281.4]
  assign _T_17810 = 7'h5 == _T_11317_63; // @[Mux.scala 46:19:@15282.4]
  assign _T_17811 = _T_17810 ? _T_10366_4 : _T_17809; // @[Mux.scala 46:16:@15283.4]
  assign _T_17812 = 7'h4 == _T_11317_63; // @[Mux.scala 46:19:@15284.4]
  assign _T_17813 = _T_17812 ? _T_10366_3 : _T_17811; // @[Mux.scala 46:16:@15285.4]
  assign _T_17814 = 7'h3 == _T_11317_63; // @[Mux.scala 46:19:@15286.4]
  assign _T_17815 = _T_17814 ? _T_10366_2 : _T_17813; // @[Mux.scala 46:16:@15287.4]
  assign _T_17816 = 7'h2 == _T_11317_63; // @[Mux.scala 46:19:@15288.4]
  assign _T_17817 = _T_17816 ? _T_10366_1 : _T_17815; // @[Mux.scala 46:16:@15289.4]
  assign _T_17818 = 7'h1 == _T_11317_63; // @[Mux.scala 46:19:@15290.4]
  assign _T_17819 = _T_17818 ? _T_10366_0 : _T_17817; // @[Mux.scala 46:16:@15291.4]
  assign _GEN_224 = _T_10362 ? _T_10641_0 : _T_17961_0; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_225 = _T_10362 ? _T_10641_1 : _T_17961_1; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_226 = _T_10362 ? _T_10641_2 : _T_17961_2; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_227 = _T_10362 ? _T_10641_3 : _T_17961_3; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_228 = _T_10362 ? _T_10641_4 : _T_17961_4; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_229 = _T_10362 ? _T_10641_5 : _T_17961_5; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_230 = _T_10362 ? _T_10641_6 : _T_17961_6; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_231 = _T_10362 ? _T_10641_7 : _T_17961_7; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_232 = _T_10362 ? _T_10641_8 : _T_17961_8; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_233 = _T_10362 ? _T_10641_9 : _T_17961_9; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_234 = _T_10362 ? _T_10641_10 : _T_17961_10; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_235 = _T_10362 ? _T_10641_11 : _T_17961_11; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_236 = _T_10362 ? _T_10641_12 : _T_17961_12; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_237 = _T_10362 ? _T_10641_13 : _T_17961_13; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_238 = _T_10362 ? _T_10641_14 : _T_17961_14; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_239 = _T_10362 ? _T_10641_15 : _T_17961_15; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_240 = _T_10362 ? _T_10641_16 : _T_17961_16; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_241 = _T_10362 ? _T_10641_17 : _T_17961_17; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_242 = _T_10362 ? _T_10641_18 : _T_17961_18; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_243 = _T_10362 ? _T_10641_19 : _T_17961_19; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_244 = _T_10362 ? _T_10641_20 : _T_17961_20; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_245 = _T_10362 ? _T_10641_21 : _T_17961_21; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_246 = _T_10362 ? _T_10641_22 : _T_17961_22; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_247 = _T_10362 ? _T_10641_23 : _T_17961_23; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_248 = _T_10362 ? _T_10641_24 : _T_17961_24; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_249 = _T_10362 ? _T_10641_25 : _T_17961_25; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_250 = _T_10362 ? _T_10641_26 : _T_17961_26; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_251 = _T_10362 ? _T_10641_27 : _T_17961_27; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_252 = _T_10362 ? _T_10641_28 : _T_17961_28; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_253 = _T_10362 ? _T_10641_29 : _T_17961_29; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_254 = _T_10362 ? _T_10641_30 : _T_17961_30; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_255 = _T_10362 ? _T_10641_31 : _T_17961_31; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@15330.4]
  assign _GEN_256 = _T_10436_0 ? _T_11519 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15365.6]
  assign _GEN_258 = _T_10436_1 ? _T_11526 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15373.6]
  assign _GEN_260 = _T_10436_2 ? _T_11536 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15381.6]
  assign _GEN_262 = _T_10436_3 ? _T_11549 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15389.6]
  assign _GEN_264 = _T_10436_4 ? _T_11565 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15397.6]
  assign _GEN_266 = _T_10436_5 ? _T_11584 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15405.6]
  assign _GEN_268 = _T_10436_6 ? _T_11606 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15413.6]
  assign _GEN_270 = _T_10436_7 ? _T_11631 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15421.6]
  assign _GEN_272 = _T_10436_8 ? _T_11659 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15429.6]
  assign _GEN_274 = _T_10436_9 ? _T_11690 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15437.6]
  assign _GEN_276 = _T_10436_10 ? _T_11724 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15445.6]
  assign _GEN_278 = _T_10436_11 ? _T_11761 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15453.6]
  assign _GEN_280 = _T_10436_12 ? _T_11801 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15461.6]
  assign _GEN_282 = _T_10436_13 ? _T_11844 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15469.6]
  assign _GEN_284 = _T_10436_14 ? _T_11890 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15477.6]
  assign _GEN_286 = _T_10436_15 ? _T_11939 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15485.6]
  assign _GEN_288 = _T_10436_16 ? _T_11991 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15493.6]
  assign _GEN_290 = _T_10436_17 ? _T_12046 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15501.6]
  assign _GEN_292 = _T_10436_18 ? _T_12104 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15509.6]
  assign _GEN_294 = _T_10436_19 ? _T_12165 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15517.6]
  assign _GEN_296 = _T_10436_20 ? _T_12229 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15525.6]
  assign _GEN_298 = _T_10436_21 ? _T_12296 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15533.6]
  assign _GEN_300 = _T_10436_22 ? _T_12366 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15541.6]
  assign _GEN_302 = _T_10436_23 ? _T_12439 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15549.6]
  assign _GEN_304 = _T_10436_24 ? _T_12515 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15557.6]
  assign _GEN_306 = _T_10436_25 ? _T_12594 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15565.6]
  assign _GEN_308 = _T_10436_26 ? _T_12676 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15573.6]
  assign _GEN_310 = _T_10436_27 ? _T_12761 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15581.6]
  assign _GEN_312 = _T_10436_28 ? _T_12849 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15589.6]
  assign _GEN_314 = _T_10436_29 ? _T_12940 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15597.6]
  assign _GEN_316 = _T_10436_30 ? _T_13034 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15605.6]
  assign _GEN_318 = _T_10436_31 ? _T_13131 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15613.6]
  assign _GEN_320 = _T_10436_32 ? _T_13231 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15621.6]
  assign _GEN_322 = _T_10436_33 ? _T_13334 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15629.6]
  assign _GEN_324 = _T_10436_34 ? _T_13440 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15637.6]
  assign _GEN_326 = _T_10436_35 ? _T_13549 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15645.6]
  assign _GEN_328 = _T_10436_36 ? _T_13661 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15653.6]
  assign _GEN_330 = _T_10436_37 ? _T_13776 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15661.6]
  assign _GEN_332 = _T_10436_38 ? _T_13894 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15669.6]
  assign _GEN_334 = _T_10436_39 ? _T_14015 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15677.6]
  assign _GEN_336 = _T_10436_40 ? _T_14139 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15685.6]
  assign _GEN_338 = _T_10436_41 ? _T_14266 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15693.6]
  assign _GEN_340 = _T_10436_42 ? _T_14396 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15701.6]
  assign _GEN_342 = _T_10436_43 ? _T_14529 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15709.6]
  assign _GEN_344 = _T_10436_44 ? _T_14665 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15717.6]
  assign _GEN_346 = _T_10436_45 ? _T_14804 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15725.6]
  assign _GEN_348 = _T_10436_46 ? _T_14946 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15733.6]
  assign _GEN_350 = _T_10436_47 ? _T_15091 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15741.6]
  assign _GEN_352 = _T_10436_48 ? _T_15239 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15749.6]
  assign _GEN_354 = _T_10436_49 ? _T_15390 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15757.6]
  assign _GEN_356 = _T_10436_50 ? _T_15544 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15765.6]
  assign _GEN_358 = _T_10436_51 ? _T_15701 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15773.6]
  assign _GEN_360 = _T_10436_52 ? _T_15861 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15781.6]
  assign _GEN_362 = _T_10436_53 ? _T_16024 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15789.6]
  assign _GEN_364 = _T_10436_54 ? _T_16190 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15797.6]
  assign _GEN_366 = _T_10436_55 ? _T_16359 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15805.6]
  assign _GEN_368 = _T_10436_56 ? _T_16531 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15813.6]
  assign _GEN_370 = _T_10436_57 ? _T_16706 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15821.6]
  assign _GEN_372 = _T_10436_58 ? _T_16884 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15829.6]
  assign _GEN_374 = _T_10436_59 ? _T_17065 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15837.6]
  assign _GEN_376 = _T_10436_60 ? _T_17249 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15845.6]
  assign _GEN_378 = _T_10436_61 ? _T_17436 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15853.6]
  assign _GEN_380 = _T_10436_62 ? _T_17626 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15861.6]
  assign _GEN_382 = _T_10436_63 ? _T_17819 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@15869.6]
  assign _T_18267 = _T_11519 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15877.4]
  assign _T_18269 = _T_11526 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15879.4]
  assign _T_18271 = _T_11536 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15881.4]
  assign _T_18273 = _T_11549 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15883.4]
  assign _T_18275 = _T_11565 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15885.4]
  assign _T_18277 = _T_11584 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15887.4]
  assign _T_18279 = _T_11606 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15889.4]
  assign _T_18281 = _T_11631 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15891.4]
  assign _T_18283 = _T_11659 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15893.4]
  assign _T_18285 = _T_11690 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15895.4]
  assign _T_18287 = _T_11724 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15897.4]
  assign _T_18289 = _T_11761 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15899.4]
  assign _T_18291 = _T_11801 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15901.4]
  assign _T_18293 = _T_11844 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15903.4]
  assign _T_18295 = _T_11890 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15905.4]
  assign _T_18297 = _T_11939 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15907.4]
  assign _T_18299 = _T_11991 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15909.4]
  assign _T_18301 = _T_12046 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15911.4]
  assign _T_18303 = _T_12104 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15913.4]
  assign _T_18305 = _T_12165 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15915.4]
  assign _T_18307 = _T_12229 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15917.4]
  assign _T_18309 = _T_12296 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15919.4]
  assign _T_18311 = _T_12366 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15921.4]
  assign _T_18313 = _T_12439 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15923.4]
  assign _T_18315 = _T_12515 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15925.4]
  assign _T_18317 = _T_12594 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15927.4]
  assign _T_18319 = _T_12676 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15929.4]
  assign _T_18321 = _T_12761 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15931.4]
  assign _T_18323 = _T_12849 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15933.4]
  assign _T_18325 = _T_12940 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15935.4]
  assign _T_18327 = _T_13034 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15937.4]
  assign _T_18329 = _T_13131 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15939.4]
  assign _T_18331 = _T_13231 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15941.4]
  assign _T_18333 = _T_13334 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15943.4]
  assign _T_18335 = _T_13440 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15945.4]
  assign _T_18337 = _T_13549 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15947.4]
  assign _T_18339 = _T_13661 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15949.4]
  assign _T_18341 = _T_13776 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15951.4]
  assign _T_18343 = _T_13894 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15953.4]
  assign _T_18345 = _T_14015 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15955.4]
  assign _T_18347 = _T_14139 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15957.4]
  assign _T_18349 = _T_14266 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15959.4]
  assign _T_18351 = _T_14396 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15961.4]
  assign _T_18353 = _T_14529 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15963.4]
  assign _T_18355 = _T_14665 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15965.4]
  assign _T_18357 = _T_14804 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15967.4]
  assign _T_18359 = _T_14946 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15969.4]
  assign _T_18361 = _T_15091 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15971.4]
  assign _T_18363 = _T_15239 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15973.4]
  assign _T_18365 = _T_15390 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15975.4]
  assign _T_18367 = _T_15544 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15977.4]
  assign _T_18369 = _T_15701 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15979.4]
  assign _T_18371 = _T_15861 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15981.4]
  assign _T_18373 = _T_16024 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15983.4]
  assign _T_18375 = _T_16190 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15985.4]
  assign _T_18377 = _T_16359 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15987.4]
  assign _T_18379 = _T_16531 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15989.4]
  assign _T_18381 = _T_16706 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15991.4]
  assign _T_18383 = _T_16884 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15993.4]
  assign _T_18385 = _T_17065 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15995.4]
  assign _T_18387 = _T_17249 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15997.4]
  assign _T_18389 = _T_17436 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@15999.4]
  assign _T_18391 = _T_17626 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@16001.4]
  assign _T_18393 = _T_17819 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@16003.4]
  assign _GEN_448 = _T_17822 ? _T_17961_0 : _T_18605_0; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_449 = _T_17822 ? _T_17961_1 : _T_18605_1; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_450 = _T_17822 ? _T_17961_2 : _T_18605_2; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_451 = _T_17822 ? _T_17961_3 : _T_18605_3; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_452 = _T_17822 ? _T_17961_4 : _T_18605_4; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_453 = _T_17822 ? _T_17961_5 : _T_18605_5; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_454 = _T_17822 ? _T_17961_6 : _T_18605_6; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_455 = _T_17822 ? _T_17961_7 : _T_18605_7; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_456 = _T_17822 ? _T_17961_8 : _T_18605_8; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_457 = _T_17822 ? _T_17961_9 : _T_18605_9; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_458 = _T_17822 ? _T_17961_10 : _T_18605_10; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_459 = _T_17822 ? _T_17961_11 : _T_18605_11; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_460 = _T_17822 ? _T_17961_12 : _T_18605_12; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_461 = _T_17822 ? _T_17961_13 : _T_18605_13; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_462 = _T_17822 ? _T_17961_14 : _T_18605_14; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_463 = _T_17822 ? _T_17961_15 : _T_18605_15; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_464 = _T_17822 ? _T_17961_16 : _T_18605_16; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_465 = _T_17822 ? _T_17961_17 : _T_18605_17; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_466 = _T_17822 ? _T_17961_18 : _T_18605_18; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_467 = _T_17822 ? _T_17961_19 : _T_18605_19; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_468 = _T_17822 ? _T_17961_20 : _T_18605_20; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_469 = _T_17822 ? _T_17961_21 : _T_18605_21; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_470 = _T_17822 ? _T_17961_22 : _T_18605_22; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_471 = _T_17822 ? _T_17961_23 : _T_18605_23; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_472 = _T_17822 ? _T_17961_24 : _T_18605_24; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_473 = _T_17822 ? _T_17961_25 : _T_18605_25; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_474 = _T_17822 ? _T_17961_26 : _T_18605_26; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_475 = _T_17822 ? _T_17961_27 : _T_18605_27; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_476 = _T_17822 ? _T_17961_28 : _T_18605_28; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_477 = _T_17822 ? _T_17961_29 : _T_18605_29; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_478 = _T_17822 ? _T_17961_30 : _T_18605_30; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign _GEN_479 = _T_17822 ? _T_17961_31 : _T_18605_31; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@16043.4]
  assign io_output_valid = _T_18396; // @[NV_NVDLA_CSC_WL_dec.scala 135:21:@16205.4]
  assign io_output_bits_mask_0 = _T_18400_0; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16206.4]
  assign io_output_bits_mask_1 = _T_18400_1; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16207.4]
  assign io_output_bits_mask_2 = _T_18400_2; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16208.4]
  assign io_output_bits_mask_3 = _T_18400_3; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16209.4]
  assign io_output_bits_mask_4 = _T_18400_4; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16210.4]
  assign io_output_bits_mask_5 = _T_18400_5; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16211.4]
  assign io_output_bits_mask_6 = _T_18400_6; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16212.4]
  assign io_output_bits_mask_7 = _T_18400_7; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16213.4]
  assign io_output_bits_mask_8 = _T_18400_8; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16214.4]
  assign io_output_bits_mask_9 = _T_18400_9; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16215.4]
  assign io_output_bits_mask_10 = _T_18400_10; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16216.4]
  assign io_output_bits_mask_11 = _T_18400_11; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16217.4]
  assign io_output_bits_mask_12 = _T_18400_12; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16218.4]
  assign io_output_bits_mask_13 = _T_18400_13; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16219.4]
  assign io_output_bits_mask_14 = _T_18400_14; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16220.4]
  assign io_output_bits_mask_15 = _T_18400_15; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16221.4]
  assign io_output_bits_mask_16 = _T_18400_16; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16222.4]
  assign io_output_bits_mask_17 = _T_18400_17; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16223.4]
  assign io_output_bits_mask_18 = _T_18400_18; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16224.4]
  assign io_output_bits_mask_19 = _T_18400_19; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16225.4]
  assign io_output_bits_mask_20 = _T_18400_20; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16226.4]
  assign io_output_bits_mask_21 = _T_18400_21; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16227.4]
  assign io_output_bits_mask_22 = _T_18400_22; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16228.4]
  assign io_output_bits_mask_23 = _T_18400_23; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16229.4]
  assign io_output_bits_mask_24 = _T_18400_24; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16230.4]
  assign io_output_bits_mask_25 = _T_18400_25; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16231.4]
  assign io_output_bits_mask_26 = _T_18400_26; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16232.4]
  assign io_output_bits_mask_27 = _T_18400_27; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16233.4]
  assign io_output_bits_mask_28 = _T_18400_28; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16234.4]
  assign io_output_bits_mask_29 = _T_18400_29; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16235.4]
  assign io_output_bits_mask_30 = _T_18400_30; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16236.4]
  assign io_output_bits_mask_31 = _T_18400_31; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16237.4]
  assign io_output_bits_mask_32 = _T_18400_32; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16238.4]
  assign io_output_bits_mask_33 = _T_18400_33; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16239.4]
  assign io_output_bits_mask_34 = _T_18400_34; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16240.4]
  assign io_output_bits_mask_35 = _T_18400_35; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16241.4]
  assign io_output_bits_mask_36 = _T_18400_36; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16242.4]
  assign io_output_bits_mask_37 = _T_18400_37; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16243.4]
  assign io_output_bits_mask_38 = _T_18400_38; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16244.4]
  assign io_output_bits_mask_39 = _T_18400_39; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16245.4]
  assign io_output_bits_mask_40 = _T_18400_40; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16246.4]
  assign io_output_bits_mask_41 = _T_18400_41; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16247.4]
  assign io_output_bits_mask_42 = _T_18400_42; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16248.4]
  assign io_output_bits_mask_43 = _T_18400_43; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16249.4]
  assign io_output_bits_mask_44 = _T_18400_44; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16250.4]
  assign io_output_bits_mask_45 = _T_18400_45; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16251.4]
  assign io_output_bits_mask_46 = _T_18400_46; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16252.4]
  assign io_output_bits_mask_47 = _T_18400_47; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16253.4]
  assign io_output_bits_mask_48 = _T_18400_48; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16254.4]
  assign io_output_bits_mask_49 = _T_18400_49; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16255.4]
  assign io_output_bits_mask_50 = _T_18400_50; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16256.4]
  assign io_output_bits_mask_51 = _T_18400_51; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16257.4]
  assign io_output_bits_mask_52 = _T_18400_52; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16258.4]
  assign io_output_bits_mask_53 = _T_18400_53; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16259.4]
  assign io_output_bits_mask_54 = _T_18400_54; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16260.4]
  assign io_output_bits_mask_55 = _T_18400_55; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16261.4]
  assign io_output_bits_mask_56 = _T_18400_56; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16262.4]
  assign io_output_bits_mask_57 = _T_18400_57; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16263.4]
  assign io_output_bits_mask_58 = _T_18400_58; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16264.4]
  assign io_output_bits_mask_59 = _T_18400_59; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16265.4]
  assign io_output_bits_mask_60 = _T_18400_60; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16266.4]
  assign io_output_bits_mask_61 = _T_18400_61; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16267.4]
  assign io_output_bits_mask_62 = _T_18400_62; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16268.4]
  assign io_output_bits_mask_63 = _T_18400_63; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@16269.4]
  assign io_output_bits_data_0 = _T_18709_0; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16302.4]
  assign io_output_bits_data_1 = _T_18709_1; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16303.4]
  assign io_output_bits_data_2 = _T_18709_2; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16304.4]
  assign io_output_bits_data_3 = _T_18709_3; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16305.4]
  assign io_output_bits_data_4 = _T_18709_4; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16306.4]
  assign io_output_bits_data_5 = _T_18709_5; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16307.4]
  assign io_output_bits_data_6 = _T_18709_6; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16308.4]
  assign io_output_bits_data_7 = _T_18709_7; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16309.4]
  assign io_output_bits_data_8 = _T_18709_8; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16310.4]
  assign io_output_bits_data_9 = _T_18709_9; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16311.4]
  assign io_output_bits_data_10 = _T_18709_10; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16312.4]
  assign io_output_bits_data_11 = _T_18709_11; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16313.4]
  assign io_output_bits_data_12 = _T_18709_12; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16314.4]
  assign io_output_bits_data_13 = _T_18709_13; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16315.4]
  assign io_output_bits_data_14 = _T_18709_14; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16316.4]
  assign io_output_bits_data_15 = _T_18709_15; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16317.4]
  assign io_output_bits_data_16 = _T_18709_16; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16318.4]
  assign io_output_bits_data_17 = _T_18709_17; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16319.4]
  assign io_output_bits_data_18 = _T_18709_18; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16320.4]
  assign io_output_bits_data_19 = _T_18709_19; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16321.4]
  assign io_output_bits_data_20 = _T_18709_20; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16322.4]
  assign io_output_bits_data_21 = _T_18709_21; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16323.4]
  assign io_output_bits_data_22 = _T_18709_22; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16324.4]
  assign io_output_bits_data_23 = _T_18709_23; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16325.4]
  assign io_output_bits_data_24 = _T_18709_24; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16326.4]
  assign io_output_bits_data_25 = _T_18709_25; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16327.4]
  assign io_output_bits_data_26 = _T_18709_26; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16328.4]
  assign io_output_bits_data_27 = _T_18709_27; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16329.4]
  assign io_output_bits_data_28 = _T_18709_28; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16330.4]
  assign io_output_bits_data_29 = _T_18709_29; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16331.4]
  assign io_output_bits_data_30 = _T_18709_30; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16332.4]
  assign io_output_bits_data_31 = _T_18709_31; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16333.4]
  assign io_output_bits_data_32 = _T_18709_32; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16334.4]
  assign io_output_bits_data_33 = _T_18709_33; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16335.4]
  assign io_output_bits_data_34 = _T_18709_34; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16336.4]
  assign io_output_bits_data_35 = _T_18709_35; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16337.4]
  assign io_output_bits_data_36 = _T_18709_36; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16338.4]
  assign io_output_bits_data_37 = _T_18709_37; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16339.4]
  assign io_output_bits_data_38 = _T_18709_38; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16340.4]
  assign io_output_bits_data_39 = _T_18709_39; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16341.4]
  assign io_output_bits_data_40 = _T_18709_40; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16342.4]
  assign io_output_bits_data_41 = _T_18709_41; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16343.4]
  assign io_output_bits_data_42 = _T_18709_42; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16344.4]
  assign io_output_bits_data_43 = _T_18709_43; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16345.4]
  assign io_output_bits_data_44 = _T_18709_44; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16346.4]
  assign io_output_bits_data_45 = _T_18709_45; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16347.4]
  assign io_output_bits_data_46 = _T_18709_46; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16348.4]
  assign io_output_bits_data_47 = _T_18709_47; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16349.4]
  assign io_output_bits_data_48 = _T_18709_48; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16350.4]
  assign io_output_bits_data_49 = _T_18709_49; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16351.4]
  assign io_output_bits_data_50 = _T_18709_50; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16352.4]
  assign io_output_bits_data_51 = _T_18709_51; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16353.4]
  assign io_output_bits_data_52 = _T_18709_52; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16354.4]
  assign io_output_bits_data_53 = _T_18709_53; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16355.4]
  assign io_output_bits_data_54 = _T_18709_54; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16356.4]
  assign io_output_bits_data_55 = _T_18709_55; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16357.4]
  assign io_output_bits_data_56 = _T_18709_56; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16358.4]
  assign io_output_bits_data_57 = _T_18709_57; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16359.4]
  assign io_output_bits_data_58 = _T_18709_58; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16360.4]
  assign io_output_bits_data_59 = _T_18709_59; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16361.4]
  assign io_output_bits_data_60 = _T_18709_60; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16362.4]
  assign io_output_bits_data_61 = _T_18709_61; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16363.4]
  assign io_output_bits_data_62 = _T_18709_62; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16364.4]
  assign io_output_bits_data_63 = _T_18709_63; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@16365.4]
  assign io_output_bits_sel_0 = _T_18605_0; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16270.4]
  assign io_output_bits_sel_1 = _T_18605_1; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16271.4]
  assign io_output_bits_sel_2 = _T_18605_2; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16272.4]
  assign io_output_bits_sel_3 = _T_18605_3; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16273.4]
  assign io_output_bits_sel_4 = _T_18605_4; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16274.4]
  assign io_output_bits_sel_5 = _T_18605_5; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16275.4]
  assign io_output_bits_sel_6 = _T_18605_6; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16276.4]
  assign io_output_bits_sel_7 = _T_18605_7; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16277.4]
  assign io_output_bits_sel_8 = _T_18605_8; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16278.4]
  assign io_output_bits_sel_9 = _T_18605_9; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16279.4]
  assign io_output_bits_sel_10 = _T_18605_10; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16280.4]
  assign io_output_bits_sel_11 = _T_18605_11; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16281.4]
  assign io_output_bits_sel_12 = _T_18605_12; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16282.4]
  assign io_output_bits_sel_13 = _T_18605_13; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16283.4]
  assign io_output_bits_sel_14 = _T_18605_14; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16284.4]
  assign io_output_bits_sel_15 = _T_18605_15; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16285.4]
  assign io_output_bits_sel_16 = _T_18605_16; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16286.4]
  assign io_output_bits_sel_17 = _T_18605_17; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16287.4]
  assign io_output_bits_sel_18 = _T_18605_18; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16288.4]
  assign io_output_bits_sel_19 = _T_18605_19; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16289.4]
  assign io_output_bits_sel_20 = _T_18605_20; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16290.4]
  assign io_output_bits_sel_21 = _T_18605_21; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16291.4]
  assign io_output_bits_sel_22 = _T_18605_22; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16292.4]
  assign io_output_bits_sel_23 = _T_18605_23; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16293.4]
  assign io_output_bits_sel_24 = _T_18605_24; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16294.4]
  assign io_output_bits_sel_25 = _T_18605_25; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16295.4]
  assign io_output_bits_sel_26 = _T_18605_26; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16296.4]
  assign io_output_bits_sel_27 = _T_18605_27; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16297.4]
  assign io_output_bits_sel_28 = _T_18605_28; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16298.4]
  assign io_output_bits_sel_29 = _T_18605_29; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16299.4]
  assign io_output_bits_sel_30 = _T_18605_30; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16300.4]
  assign io_output_bits_sel_31 = _T_18605_31; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@16301.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_10366_0 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_10366_1 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_10366_2 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_10366_3 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_10366_4 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_10366_5 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_10366_6 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_10366_7 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_10366_8 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_10366_9 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_10366_10 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_10366_11 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_10366_12 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_10366_13 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_10366_14 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_10366_15 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_10366_16 = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_10366_17 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_10366_18 = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_10366_19 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_10366_20 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_10366_21 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_10366_22 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_10366_23 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_10366_24 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_10366_25 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_10366_26 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_10366_27 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_10366_28 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_10366_29 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_10366_30 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_10366_31 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_10366_32 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_10366_33 = _RAND_34[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_10366_34 = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_10366_35 = _RAND_36[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_10366_36 = _RAND_37[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_10366_37 = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_10366_38 = _RAND_39[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_10366_39 = _RAND_40[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_10366_40 = _RAND_41[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_10366_41 = _RAND_42[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_10366_42 = _RAND_43[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_10366_43 = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_10366_44 = _RAND_45[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_10366_45 = _RAND_46[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_10366_46 = _RAND_47[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_10366_47 = _RAND_48[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_10366_48 = _RAND_49[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_10366_49 = _RAND_50[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_10366_50 = _RAND_51[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_10366_51 = _RAND_52[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_10366_52 = _RAND_53[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_10366_53 = _RAND_54[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_10366_54 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_10366_55 = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_10366_56 = _RAND_57[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_10366_57 = _RAND_58[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_10366_58 = _RAND_59[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_10366_59 = _RAND_60[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_10366_60 = _RAND_61[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_10366_61 = _RAND_62[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_10366_62 = _RAND_63[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_10366_63 = _RAND_64[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_10436_0 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_10436_1 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_10436_2 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_10436_3 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_10436_4 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_10436_5 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_10436_6 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_10436_7 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_10436_8 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_10436_9 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_10436_10 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_10436_11 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_10436_12 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_10436_13 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_10436_14 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_10436_15 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_10436_16 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_10436_17 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_10436_18 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_10436_19 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_10436_20 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_10436_21 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_10436_22 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_10436_23 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_10436_24 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_10436_25 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_10436_26 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_10436_27 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_10436_28 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_10436_29 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_10436_30 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_10436_31 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_10436_32 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_10436_33 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_10436_34 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_10436_35 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_10436_36 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_10436_37 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_10436_38 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_10436_39 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_10436_40 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_10436_41 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_10436_42 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_10436_43 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_10436_44 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_10436_45 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_10436_46 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_10436_47 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_10436_48 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_10436_49 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_10436_50 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_10436_51 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_10436_52 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_10436_53 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_10436_54 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_10436_55 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_10436_56 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_10436_57 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_10436_58 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_10436_59 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_10436_60 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_10436_61 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_10436_62 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_10436_63 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_10641_0 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_10641_1 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_10641_2 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_10641_3 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_10641_4 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_10641_5 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_10641_6 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_10641_7 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_10641_8 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_10641_9 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_10641_10 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_10641_11 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_10641_12 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_10641_13 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_10641_14 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_10641_15 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_10641_16 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_10641_17 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_10641_18 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_10641_19 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_10641_20 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_10641_21 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_10641_22 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_10641_23 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_10641_24 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_10641_25 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_10641_26 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_10641_27 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_10641_28 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_10641_29 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_10641_30 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_10641_31 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_11317_63 = _RAND_161[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_11317_62 = _RAND_162[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_11317_61 = _RAND_163[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_11317_60 = _RAND_164[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_11317_59 = _RAND_165[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_11317_58 = _RAND_166[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_11317_57 = _RAND_167[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_11317_56 = _RAND_168[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_11317_55 = _RAND_169[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_11317_54 = _RAND_170[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_11317_53 = _RAND_171[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_11317_52 = _RAND_172[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_11317_51 = _RAND_173[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_11317_50 = _RAND_174[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_11317_49 = _RAND_175[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_11317_48 = _RAND_176[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_11317_47 = _RAND_177[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_11317_46 = _RAND_178[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_11317_45 = _RAND_179[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_11317_44 = _RAND_180[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_11317_43 = _RAND_181[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_11317_42 = _RAND_182[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_11317_41 = _RAND_183[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_11317_40 = _RAND_184[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_11317_39 = _RAND_185[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_11317_38 = _RAND_186[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_11317_37 = _RAND_187[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_11317_36 = _RAND_188[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_11317_35 = _RAND_189[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_11317_34 = _RAND_190[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_11317_33 = _RAND_191[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_11317_32 = _RAND_192[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_11317_31 = _RAND_193[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_11317_30 = _RAND_194[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_11317_29 = _RAND_195[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_11317_28 = _RAND_196[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_11317_27 = _RAND_197[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_11317_26 = _RAND_198[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_11317_25 = _RAND_199[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_11317_24 = _RAND_200[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_11317_23 = _RAND_201[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_11317_22 = _RAND_202[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_11317_21 = _RAND_203[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_11317_20 = _RAND_204[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_11317_19 = _RAND_205[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_11317_18 = _RAND_206[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_11317_17 = _RAND_207[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_11317_16 = _RAND_208[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_11317_15 = _RAND_209[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_11317_14 = _RAND_210[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_11317_13 = _RAND_211[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_11317_12 = _RAND_212[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_11317_11 = _RAND_213[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_11317_10 = _RAND_214[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_11317_9 = _RAND_215[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_11317_8 = _RAND_216[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_11317_7 = _RAND_217[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_11317_6 = _RAND_218[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_11317_5 = _RAND_219[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_11317_4 = _RAND_220[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_11317_3 = _RAND_221[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_11317_2 = _RAND_222[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_11317_1 = _RAND_223[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_11317_0 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_17822 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_17961_0 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_17961_1 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_17961_2 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_17961_3 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_17961_4 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_17961_5 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_17961_6 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_17961_7 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_17961_8 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_17961_9 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_17961_10 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_17961_11 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_17961_12 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_17961_13 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_17961_14 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_17961_15 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_17961_16 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_17961_17 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_17961_18 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_17961_19 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_17961_20 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_17961_21 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_17961_22 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_17961_23 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_17961_24 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_17961_25 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_17961_26 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_17961_27 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_17961_28 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_17961_29 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_17961_30 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_17961_31 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_18065_0 = _RAND_258[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_18065_1 = _RAND_259[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_18065_2 = _RAND_260[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_18065_3 = _RAND_261[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_18065_4 = _RAND_262[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_18065_5 = _RAND_263[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_18065_6 = _RAND_264[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_18065_7 = _RAND_265[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_18065_8 = _RAND_266[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_18065_9 = _RAND_267[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_18065_10 = _RAND_268[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_18065_11 = _RAND_269[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_18065_12 = _RAND_270[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_18065_13 = _RAND_271[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_18065_14 = _RAND_272[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_18065_15 = _RAND_273[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_18065_16 = _RAND_274[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_18065_17 = _RAND_275[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_18065_18 = _RAND_276[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_18065_19 = _RAND_277[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_18065_20 = _RAND_278[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_18065_21 = _RAND_279[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_18065_22 = _RAND_280[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_18065_23 = _RAND_281[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_18065_24 = _RAND_282[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_18065_25 = _RAND_283[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_18065_26 = _RAND_284[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_18065_27 = _RAND_285[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_18065_28 = _RAND_286[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_18065_29 = _RAND_287[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_18065_30 = _RAND_288[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_18065_31 = _RAND_289[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_18065_32 = _RAND_290[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_18065_33 = _RAND_291[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_18065_34 = _RAND_292[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_18065_35 = _RAND_293[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_18065_36 = _RAND_294[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_18065_37 = _RAND_295[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_18065_38 = _RAND_296[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_18065_39 = _RAND_297[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_18065_40 = _RAND_298[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_18065_41 = _RAND_299[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_18065_42 = _RAND_300[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_18065_43 = _RAND_301[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_18065_44 = _RAND_302[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_18065_45 = _RAND_303[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_18065_46 = _RAND_304[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_18065_47 = _RAND_305[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_18065_48 = _RAND_306[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_18065_49 = _RAND_307[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_18065_50 = _RAND_308[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_18065_51 = _RAND_309[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_18065_52 = _RAND_310[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_18065_53 = _RAND_311[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_18065_54 = _RAND_312[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_18065_55 = _RAND_313[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_18065_56 = _RAND_314[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_18065_57 = _RAND_315[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_18065_58 = _RAND_316[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_18065_59 = _RAND_317[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_18065_60 = _RAND_318[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_18065_61 = _RAND_319[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_18065_62 = _RAND_320[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_18065_63 = _RAND_321[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_18396 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_18400_0 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_18400_1 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_18400_2 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_18400_3 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_18400_4 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_18400_5 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_18400_6 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_18400_7 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_18400_8 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_18400_9 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_18400_10 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_18400_11 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_18400_12 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_18400_13 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_18400_14 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_18400_15 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_18400_16 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_18400_17 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_18400_18 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_18400_19 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_18400_20 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_18400_21 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_18400_22 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_18400_23 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_18400_24 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_18400_25 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_18400_26 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_18400_27 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_18400_28 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_18400_29 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_18400_30 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_18400_31 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_18400_32 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_18400_33 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_18400_34 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_18400_35 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_18400_36 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_18400_37 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_18400_38 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_18400_39 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_18400_40 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_18400_41 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_18400_42 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_18400_43 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_18400_44 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_18400_45 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_18400_46 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_18400_47 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_18400_48 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_18400_49 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_18400_50 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_18400_51 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_18400_52 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_18400_53 = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_18400_54 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_18400_55 = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_18400_56 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_18400_57 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_18400_58 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_18400_59 = _RAND_382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_18400_60 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_18400_61 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_18400_62 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_18400_63 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_18605_0 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_18605_1 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_18605_2 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_18605_3 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_18605_4 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_18605_5 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_18605_6 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_18605_7 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_18605_8 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_18605_9 = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_18605_10 = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_18605_11 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_18605_12 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_18605_13 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_18605_14 = _RAND_401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_18605_15 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_18605_16 = _RAND_403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_18605_17 = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_18605_18 = _RAND_405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_18605_19 = _RAND_406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_18605_20 = _RAND_407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_18605_21 = _RAND_408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_18605_22 = _RAND_409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_18605_23 = _RAND_410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_18605_24 = _RAND_411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_18605_25 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_18605_26 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_18605_27 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_18605_28 = _RAND_415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_18605_29 = _RAND_416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_18605_30 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_18605_31 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_18709_0 = _RAND_419[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_18709_1 = _RAND_420[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_18709_2 = _RAND_421[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_18709_3 = _RAND_422[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_18709_4 = _RAND_423[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_18709_5 = _RAND_424[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_18709_6 = _RAND_425[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_18709_7 = _RAND_426[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_18709_8 = _RAND_427[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_18709_9 = _RAND_428[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_18709_10 = _RAND_429[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_18709_11 = _RAND_430[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_18709_12 = _RAND_431[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_18709_13 = _RAND_432[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_18709_14 = _RAND_433[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_18709_15 = _RAND_434[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_18709_16 = _RAND_435[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_18709_17 = _RAND_436[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_18709_18 = _RAND_437[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_18709_19 = _RAND_438[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_18709_20 = _RAND_439[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_18709_21 = _RAND_440[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_18709_22 = _RAND_441[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_18709_23 = _RAND_442[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_18709_24 = _RAND_443[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_18709_25 = _RAND_444[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_18709_26 = _RAND_445[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_18709_27 = _RAND_446[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_18709_28 = _RAND_447[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_18709_29 = _RAND_448[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_18709_30 = _RAND_449[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_18709_31 = _RAND_450[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_18709_32 = _RAND_451[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_18709_33 = _RAND_452[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_18709_34 = _RAND_453[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_18709_35 = _RAND_454[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_18709_36 = _RAND_455[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_18709_37 = _RAND_456[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_18709_38 = _RAND_457[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_18709_39 = _RAND_458[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_18709_40 = _RAND_459[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_18709_41 = _RAND_460[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_18709_42 = _RAND_461[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_18709_43 = _RAND_462[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_18709_44 = _RAND_463[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_18709_45 = _RAND_464[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_18709_46 = _RAND_465[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_18709_47 = _RAND_466[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_18709_48 = _RAND_467[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_18709_49 = _RAND_468[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_18709_50 = _RAND_469[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_18709_51 = _RAND_470[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_18709_52 = _RAND_471[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_18709_53 = _RAND_472[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_18709_54 = _RAND_473[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_18709_55 = _RAND_474[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_18709_56 = _RAND_475[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_18709_57 = _RAND_476[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_18709_58 = _RAND_477[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_18709_59 = _RAND_478[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_18709_60 = _RAND_479[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_18709_61 = _RAND_480[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_18709_62 = _RAND_481[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_18709_63 = _RAND_482[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_10362 <= 1'h0;
    end else begin
      _T_10362 <= io_input_valid;
    end
    if (io_input_valid) begin
      _T_10366_0 <= io_input_bits_data_0;
    end
    if (io_input_valid) begin
      _T_10366_1 <= io_input_bits_data_1;
    end
    if (io_input_valid) begin
      _T_10366_2 <= io_input_bits_data_2;
    end
    if (io_input_valid) begin
      _T_10366_3 <= io_input_bits_data_3;
    end
    if (io_input_valid) begin
      _T_10366_4 <= io_input_bits_data_4;
    end
    if (io_input_valid) begin
      _T_10366_5 <= io_input_bits_data_5;
    end
    if (io_input_valid) begin
      _T_10366_6 <= io_input_bits_data_6;
    end
    if (io_input_valid) begin
      _T_10366_7 <= io_input_bits_data_7;
    end
    if (io_input_valid) begin
      _T_10366_8 <= io_input_bits_data_8;
    end
    if (io_input_valid) begin
      _T_10366_9 <= io_input_bits_data_9;
    end
    if (io_input_valid) begin
      _T_10366_10 <= io_input_bits_data_10;
    end
    if (io_input_valid) begin
      _T_10366_11 <= io_input_bits_data_11;
    end
    if (io_input_valid) begin
      _T_10366_12 <= io_input_bits_data_12;
    end
    if (io_input_valid) begin
      _T_10366_13 <= io_input_bits_data_13;
    end
    if (io_input_valid) begin
      _T_10366_14 <= io_input_bits_data_14;
    end
    if (io_input_valid) begin
      _T_10366_15 <= io_input_bits_data_15;
    end
    if (io_input_valid) begin
      _T_10366_16 <= io_input_bits_data_16;
    end
    if (io_input_valid) begin
      _T_10366_17 <= io_input_bits_data_17;
    end
    if (io_input_valid) begin
      _T_10366_18 <= io_input_bits_data_18;
    end
    if (io_input_valid) begin
      _T_10366_19 <= io_input_bits_data_19;
    end
    if (io_input_valid) begin
      _T_10366_20 <= io_input_bits_data_20;
    end
    if (io_input_valid) begin
      _T_10366_21 <= io_input_bits_data_21;
    end
    if (io_input_valid) begin
      _T_10366_22 <= io_input_bits_data_22;
    end
    if (io_input_valid) begin
      _T_10366_23 <= io_input_bits_data_23;
    end
    if (io_input_valid) begin
      _T_10366_24 <= io_input_bits_data_24;
    end
    if (io_input_valid) begin
      _T_10366_25 <= io_input_bits_data_25;
    end
    if (io_input_valid) begin
      _T_10366_26 <= io_input_bits_data_26;
    end
    if (io_input_valid) begin
      _T_10366_27 <= io_input_bits_data_27;
    end
    if (io_input_valid) begin
      _T_10366_28 <= io_input_bits_data_28;
    end
    if (io_input_valid) begin
      _T_10366_29 <= io_input_bits_data_29;
    end
    if (io_input_valid) begin
      _T_10366_30 <= io_input_bits_data_30;
    end
    if (io_input_valid) begin
      _T_10366_31 <= io_input_bits_data_31;
    end
    if (io_input_valid) begin
      _T_10366_32 <= io_input_bits_data_32;
    end
    if (io_input_valid) begin
      _T_10366_33 <= io_input_bits_data_33;
    end
    if (io_input_valid) begin
      _T_10366_34 <= io_input_bits_data_34;
    end
    if (io_input_valid) begin
      _T_10366_35 <= io_input_bits_data_35;
    end
    if (io_input_valid) begin
      _T_10366_36 <= io_input_bits_data_36;
    end
    if (io_input_valid) begin
      _T_10366_37 <= io_input_bits_data_37;
    end
    if (io_input_valid) begin
      _T_10366_38 <= io_input_bits_data_38;
    end
    if (io_input_valid) begin
      _T_10366_39 <= io_input_bits_data_39;
    end
    if (io_input_valid) begin
      _T_10366_40 <= io_input_bits_data_40;
    end
    if (io_input_valid) begin
      _T_10366_41 <= io_input_bits_data_41;
    end
    if (io_input_valid) begin
      _T_10366_42 <= io_input_bits_data_42;
    end
    if (io_input_valid) begin
      _T_10366_43 <= io_input_bits_data_43;
    end
    if (io_input_valid) begin
      _T_10366_44 <= io_input_bits_data_44;
    end
    if (io_input_valid) begin
      _T_10366_45 <= io_input_bits_data_45;
    end
    if (io_input_valid) begin
      _T_10366_46 <= io_input_bits_data_46;
    end
    if (io_input_valid) begin
      _T_10366_47 <= io_input_bits_data_47;
    end
    if (io_input_valid) begin
      _T_10366_48 <= io_input_bits_data_48;
    end
    if (io_input_valid) begin
      _T_10366_49 <= io_input_bits_data_49;
    end
    if (io_input_valid) begin
      _T_10366_50 <= io_input_bits_data_50;
    end
    if (io_input_valid) begin
      _T_10366_51 <= io_input_bits_data_51;
    end
    if (io_input_valid) begin
      _T_10366_52 <= io_input_bits_data_52;
    end
    if (io_input_valid) begin
      _T_10366_53 <= io_input_bits_data_53;
    end
    if (io_input_valid) begin
      _T_10366_54 <= io_input_bits_data_54;
    end
    if (io_input_valid) begin
      _T_10366_55 <= io_input_bits_data_55;
    end
    if (io_input_valid) begin
      _T_10366_56 <= io_input_bits_data_56;
    end
    if (io_input_valid) begin
      _T_10366_57 <= io_input_bits_data_57;
    end
    if (io_input_valid) begin
      _T_10366_58 <= io_input_bits_data_58;
    end
    if (io_input_valid) begin
      _T_10366_59 <= io_input_bits_data_59;
    end
    if (io_input_valid) begin
      _T_10366_60 <= io_input_bits_data_60;
    end
    if (io_input_valid) begin
      _T_10366_61 <= io_input_bits_data_61;
    end
    if (io_input_valid) begin
      _T_10366_62 <= io_input_bits_data_62;
    end
    if (io_input_valid) begin
      _T_10366_63 <= io_input_bits_data_63;
    end
    if (io_input_valid) begin
      _T_10436_0 <= io_input_bits_mask_0;
    end
    if (io_input_valid) begin
      _T_10436_1 <= io_input_bits_mask_1;
    end
    if (io_input_valid) begin
      _T_10436_2 <= io_input_bits_mask_2;
    end
    if (io_input_valid) begin
      _T_10436_3 <= io_input_bits_mask_3;
    end
    if (io_input_valid) begin
      _T_10436_4 <= io_input_bits_mask_4;
    end
    if (io_input_valid) begin
      _T_10436_5 <= io_input_bits_mask_5;
    end
    if (io_input_valid) begin
      _T_10436_6 <= io_input_bits_mask_6;
    end
    if (io_input_valid) begin
      _T_10436_7 <= io_input_bits_mask_7;
    end
    if (io_input_valid) begin
      _T_10436_8 <= io_input_bits_mask_8;
    end
    if (io_input_valid) begin
      _T_10436_9 <= io_input_bits_mask_9;
    end
    if (io_input_valid) begin
      _T_10436_10 <= io_input_bits_mask_10;
    end
    if (io_input_valid) begin
      _T_10436_11 <= io_input_bits_mask_11;
    end
    if (io_input_valid) begin
      _T_10436_12 <= io_input_bits_mask_12;
    end
    if (io_input_valid) begin
      _T_10436_13 <= io_input_bits_mask_13;
    end
    if (io_input_valid) begin
      _T_10436_14 <= io_input_bits_mask_14;
    end
    if (io_input_valid) begin
      _T_10436_15 <= io_input_bits_mask_15;
    end
    if (io_input_valid) begin
      _T_10436_16 <= io_input_bits_mask_16;
    end
    if (io_input_valid) begin
      _T_10436_17 <= io_input_bits_mask_17;
    end
    if (io_input_valid) begin
      _T_10436_18 <= io_input_bits_mask_18;
    end
    if (io_input_valid) begin
      _T_10436_19 <= io_input_bits_mask_19;
    end
    if (io_input_valid) begin
      _T_10436_20 <= io_input_bits_mask_20;
    end
    if (io_input_valid) begin
      _T_10436_21 <= io_input_bits_mask_21;
    end
    if (io_input_valid) begin
      _T_10436_22 <= io_input_bits_mask_22;
    end
    if (io_input_valid) begin
      _T_10436_23 <= io_input_bits_mask_23;
    end
    if (io_input_valid) begin
      _T_10436_24 <= io_input_bits_mask_24;
    end
    if (io_input_valid) begin
      _T_10436_25 <= io_input_bits_mask_25;
    end
    if (io_input_valid) begin
      _T_10436_26 <= io_input_bits_mask_26;
    end
    if (io_input_valid) begin
      _T_10436_27 <= io_input_bits_mask_27;
    end
    if (io_input_valid) begin
      _T_10436_28 <= io_input_bits_mask_28;
    end
    if (io_input_valid) begin
      _T_10436_29 <= io_input_bits_mask_29;
    end
    if (io_input_valid) begin
      _T_10436_30 <= io_input_bits_mask_30;
    end
    if (io_input_valid) begin
      _T_10436_31 <= io_input_bits_mask_31;
    end
    if (io_input_valid) begin
      _T_10436_32 <= io_input_bits_mask_32;
    end
    if (io_input_valid) begin
      _T_10436_33 <= io_input_bits_mask_33;
    end
    if (io_input_valid) begin
      _T_10436_34 <= io_input_bits_mask_34;
    end
    if (io_input_valid) begin
      _T_10436_35 <= io_input_bits_mask_35;
    end
    if (io_input_valid) begin
      _T_10436_36 <= io_input_bits_mask_36;
    end
    if (io_input_valid) begin
      _T_10436_37 <= io_input_bits_mask_37;
    end
    if (io_input_valid) begin
      _T_10436_38 <= io_input_bits_mask_38;
    end
    if (io_input_valid) begin
      _T_10436_39 <= io_input_bits_mask_39;
    end
    if (io_input_valid) begin
      _T_10436_40 <= io_input_bits_mask_40;
    end
    if (io_input_valid) begin
      _T_10436_41 <= io_input_bits_mask_41;
    end
    if (io_input_valid) begin
      _T_10436_42 <= io_input_bits_mask_42;
    end
    if (io_input_valid) begin
      _T_10436_43 <= io_input_bits_mask_43;
    end
    if (io_input_valid) begin
      _T_10436_44 <= io_input_bits_mask_44;
    end
    if (io_input_valid) begin
      _T_10436_45 <= io_input_bits_mask_45;
    end
    if (io_input_valid) begin
      _T_10436_46 <= io_input_bits_mask_46;
    end
    if (io_input_valid) begin
      _T_10436_47 <= io_input_bits_mask_47;
    end
    if (io_input_valid) begin
      _T_10436_48 <= io_input_bits_mask_48;
    end
    if (io_input_valid) begin
      _T_10436_49 <= io_input_bits_mask_49;
    end
    if (io_input_valid) begin
      _T_10436_50 <= io_input_bits_mask_50;
    end
    if (io_input_valid) begin
      _T_10436_51 <= io_input_bits_mask_51;
    end
    if (io_input_valid) begin
      _T_10436_52 <= io_input_bits_mask_52;
    end
    if (io_input_valid) begin
      _T_10436_53 <= io_input_bits_mask_53;
    end
    if (io_input_valid) begin
      _T_10436_54 <= io_input_bits_mask_54;
    end
    if (io_input_valid) begin
      _T_10436_55 <= io_input_bits_mask_55;
    end
    if (io_input_valid) begin
      _T_10436_56 <= io_input_bits_mask_56;
    end
    if (io_input_valid) begin
      _T_10436_57 <= io_input_bits_mask_57;
    end
    if (io_input_valid) begin
      _T_10436_58 <= io_input_bits_mask_58;
    end
    if (io_input_valid) begin
      _T_10436_59 <= io_input_bits_mask_59;
    end
    if (io_input_valid) begin
      _T_10436_60 <= io_input_bits_mask_60;
    end
    if (io_input_valid) begin
      _T_10436_61 <= io_input_bits_mask_61;
    end
    if (io_input_valid) begin
      _T_10436_62 <= io_input_bits_mask_62;
    end
    if (io_input_valid) begin
      _T_10436_63 <= io_input_bits_mask_63;
    end
    if (reset) begin
      _T_10641_0 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_0 <= io_input_bits_sel_0;
      end
    end
    if (reset) begin
      _T_10641_1 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_1 <= io_input_bits_sel_1;
      end
    end
    if (reset) begin
      _T_10641_2 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_2 <= io_input_bits_sel_2;
      end
    end
    if (reset) begin
      _T_10641_3 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_3 <= io_input_bits_sel_3;
      end
    end
    if (reset) begin
      _T_10641_4 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_4 <= io_input_bits_sel_4;
      end
    end
    if (reset) begin
      _T_10641_5 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_5 <= io_input_bits_sel_5;
      end
    end
    if (reset) begin
      _T_10641_6 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_6 <= io_input_bits_sel_6;
      end
    end
    if (reset) begin
      _T_10641_7 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_7 <= io_input_bits_sel_7;
      end
    end
    if (reset) begin
      _T_10641_8 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_8 <= io_input_bits_sel_8;
      end
    end
    if (reset) begin
      _T_10641_9 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_9 <= io_input_bits_sel_9;
      end
    end
    if (reset) begin
      _T_10641_10 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_10 <= io_input_bits_sel_10;
      end
    end
    if (reset) begin
      _T_10641_11 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_11 <= io_input_bits_sel_11;
      end
    end
    if (reset) begin
      _T_10641_12 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_12 <= io_input_bits_sel_12;
      end
    end
    if (reset) begin
      _T_10641_13 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_13 <= io_input_bits_sel_13;
      end
    end
    if (reset) begin
      _T_10641_14 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_14 <= io_input_bits_sel_14;
      end
    end
    if (reset) begin
      _T_10641_15 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_15 <= io_input_bits_sel_15;
      end
    end
    if (reset) begin
      _T_10641_16 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_16 <= io_input_bits_sel_16;
      end
    end
    if (reset) begin
      _T_10641_17 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_17 <= io_input_bits_sel_17;
      end
    end
    if (reset) begin
      _T_10641_18 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_18 <= io_input_bits_sel_18;
      end
    end
    if (reset) begin
      _T_10641_19 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_19 <= io_input_bits_sel_19;
      end
    end
    if (reset) begin
      _T_10641_20 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_20 <= io_input_bits_sel_20;
      end
    end
    if (reset) begin
      _T_10641_21 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_21 <= io_input_bits_sel_21;
      end
    end
    if (reset) begin
      _T_10641_22 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_22 <= io_input_bits_sel_22;
      end
    end
    if (reset) begin
      _T_10641_23 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_23 <= io_input_bits_sel_23;
      end
    end
    if (reset) begin
      _T_10641_24 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_24 <= io_input_bits_sel_24;
      end
    end
    if (reset) begin
      _T_10641_25 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_25 <= io_input_bits_sel_25;
      end
    end
    if (reset) begin
      _T_10641_26 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_26 <= io_input_bits_sel_26;
      end
    end
    if (reset) begin
      _T_10641_27 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_27 <= io_input_bits_sel_27;
      end
    end
    if (reset) begin
      _T_10641_28 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_28 <= io_input_bits_sel_28;
      end
    end
    if (reset) begin
      _T_10641_29 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_29 <= io_input_bits_sel_29;
      end
    end
    if (reset) begin
      _T_10641_30 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_30 <= io_input_bits_sel_30;
      end
    end
    if (reset) begin
      _T_10641_31 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_31 <= io_input_bits_sel_31;
      end
    end
    if (reset) begin
      _T_11317_63 <= 7'h0;
    end else begin
      if (_T_11431) begin
        _T_11317_63 <= _T_10359;
      end
    end
    if (reset) begin
      _T_11317_62 <= 6'h0;
    end else begin
      if (_T_11431) begin
        _T_11317_62 <= _T_2167_62;
      end
    end
    if (reset) begin
      _T_11317_61 <= 6'h0;
    end else begin
      if (_T_11431) begin
        _T_11317_61 <= _T_2167_61;
      end
    end
    if (reset) begin
      _T_11317_60 <= 6'h0;
    end else begin
      if (_T_11431) begin
        _T_11317_60 <= _T_2167_60;
      end
    end
    if (reset) begin
      _T_11317_59 <= 6'h0;
    end else begin
      if (_T_11431) begin
        _T_11317_59 <= _T_2167_59;
      end
    end
    if (reset) begin
      _T_11317_58 <= 6'h0;
    end else begin
      if (_T_11431) begin
        _T_11317_58 <= _T_2167_58;
      end
    end
    if (reset) begin
      _T_11317_57 <= 6'h0;
    end else begin
      if (_T_11431) begin
        _T_11317_57 <= _T_2167_57;
      end
    end
    if (reset) begin
      _T_11317_56 <= 6'h0;
    end else begin
      if (_T_11431) begin
        _T_11317_56 <= _T_2167_56;
      end
    end
    if (reset) begin
      _T_11317_55 <= 6'h0;
    end else begin
      if (_T_11415) begin
        _T_11317_55 <= _T_2167_55;
      end
    end
    if (reset) begin
      _T_11317_54 <= 6'h0;
    end else begin
      if (_T_11415) begin
        _T_11317_54 <= _T_2167_54;
      end
    end
    if (reset) begin
      _T_11317_53 <= 6'h0;
    end else begin
      if (_T_11415) begin
        _T_11317_53 <= _T_2167_53;
      end
    end
    if (reset) begin
      _T_11317_52 <= 6'h0;
    end else begin
      if (_T_11415) begin
        _T_11317_52 <= _T_2167_52;
      end
    end
    if (reset) begin
      _T_11317_51 <= 6'h0;
    end else begin
      if (_T_11415) begin
        _T_11317_51 <= _T_2167_51;
      end
    end
    if (reset) begin
      _T_11317_50 <= 6'h0;
    end else begin
      if (_T_11415) begin
        _T_11317_50 <= _T_2167_50;
      end
    end
    if (reset) begin
      _T_11317_49 <= 6'h0;
    end else begin
      if (_T_11415) begin
        _T_11317_49 <= _T_2167_49;
      end
    end
    if (reset) begin
      _T_11317_48 <= 6'h0;
    end else begin
      if (_T_11415) begin
        _T_11317_48 <= _T_2167_48;
      end
    end
    if (reset) begin
      _T_11317_47 <= 6'h0;
    end else begin
      if (_T_11399) begin
        _T_11317_47 <= _T_2167_47;
      end
    end
    if (reset) begin
      _T_11317_46 <= 6'h0;
    end else begin
      if (_T_11399) begin
        _T_11317_46 <= _T_2167_46;
      end
    end
    if (reset) begin
      _T_11317_45 <= 6'h0;
    end else begin
      if (_T_11399) begin
        _T_11317_45 <= _T_2167_45;
      end
    end
    if (reset) begin
      _T_11317_44 <= 6'h0;
    end else begin
      if (_T_11399) begin
        _T_11317_44 <= _T_2167_44;
      end
    end
    if (reset) begin
      _T_11317_43 <= 6'h0;
    end else begin
      if (_T_11399) begin
        _T_11317_43 <= _T_2167_43;
      end
    end
    if (reset) begin
      _T_11317_42 <= 6'h0;
    end else begin
      if (_T_11399) begin
        _T_11317_42 <= _T_2167_42;
      end
    end
    if (reset) begin
      _T_11317_41 <= 6'h0;
    end else begin
      if (_T_11399) begin
        _T_11317_41 <= _T_2167_41;
      end
    end
    if (reset) begin
      _T_11317_40 <= 6'h0;
    end else begin
      if (_T_11399) begin
        _T_11317_40 <= _T_2167_40;
      end
    end
    if (reset) begin
      _T_11317_39 <= 6'h0;
    end else begin
      if (_T_11383) begin
        _T_11317_39 <= _T_2167_39;
      end
    end
    if (reset) begin
      _T_11317_38 <= 6'h0;
    end else begin
      if (_T_11383) begin
        _T_11317_38 <= _T_2167_38;
      end
    end
    if (reset) begin
      _T_11317_37 <= 6'h0;
    end else begin
      if (_T_11383) begin
        _T_11317_37 <= _T_2167_37;
      end
    end
    if (reset) begin
      _T_11317_36 <= 6'h0;
    end else begin
      if (_T_11383) begin
        _T_11317_36 <= _T_2167_36;
      end
    end
    if (reset) begin
      _T_11317_35 <= 6'h0;
    end else begin
      if (_T_11383) begin
        _T_11317_35 <= _T_2167_35;
      end
    end
    if (reset) begin
      _T_11317_34 <= 6'h0;
    end else begin
      if (_T_11383) begin
        _T_11317_34 <= _T_2167_34;
      end
    end
    if (reset) begin
      _T_11317_33 <= 6'h0;
    end else begin
      if (_T_11383) begin
        _T_11317_33 <= _T_2167_33;
      end
    end
    if (reset) begin
      _T_11317_32 <= 6'h0;
    end else begin
      if (_T_11383) begin
        _T_11317_32 <= _T_2167_32;
      end
    end
    if (reset) begin
      _T_11317_31 <= 6'h0;
    end else begin
      if (_T_11367) begin
        _T_11317_31 <= _T_5239;
      end
    end
    if (reset) begin
      _T_11317_30 <= 5'h0;
    end else begin
      if (_T_11367) begin
        _T_11317_30 <= _T_2167_30;
      end
    end
    if (reset) begin
      _T_11317_29 <= 5'h0;
    end else begin
      if (_T_11367) begin
        _T_11317_29 <= _T_2167_29;
      end
    end
    if (reset) begin
      _T_11317_28 <= 5'h0;
    end else begin
      if (_T_11367) begin
        _T_11317_28 <= _T_2167_28;
      end
    end
    if (reset) begin
      _T_11317_27 <= 5'h0;
    end else begin
      if (_T_11367) begin
        _T_11317_27 <= _T_2167_27;
      end
    end
    if (reset) begin
      _T_11317_26 <= 5'h0;
    end else begin
      if (_T_11367) begin
        _T_11317_26 <= _T_2167_26;
      end
    end
    if (reset) begin
      _T_11317_25 <= 5'h0;
    end else begin
      if (_T_11367) begin
        _T_11317_25 <= _T_2167_25;
      end
    end
    if (reset) begin
      _T_11317_24 <= 5'h0;
    end else begin
      if (_T_11367) begin
        _T_11317_24 <= _T_2167_24;
      end
    end
    if (reset) begin
      _T_11317_23 <= 5'h0;
    end else begin
      if (_T_11351) begin
        _T_11317_23 <= _T_2167_23;
      end
    end
    if (reset) begin
      _T_11317_22 <= 5'h0;
    end else begin
      if (_T_11351) begin
        _T_11317_22 <= _T_2167_22;
      end
    end
    if (reset) begin
      _T_11317_21 <= 5'h0;
    end else begin
      if (_T_11351) begin
        _T_11317_21 <= _T_2167_21;
      end
    end
    if (reset) begin
      _T_11317_20 <= 5'h0;
    end else begin
      if (_T_11351) begin
        _T_11317_20 <= _T_2167_20;
      end
    end
    if (reset) begin
      _T_11317_19 <= 5'h0;
    end else begin
      if (_T_11351) begin
        _T_11317_19 <= _T_2167_19;
      end
    end
    if (reset) begin
      _T_11317_18 <= 5'h0;
    end else begin
      if (_T_11351) begin
        _T_11317_18 <= _T_2167_18;
      end
    end
    if (reset) begin
      _T_11317_17 <= 5'h0;
    end else begin
      if (_T_11351) begin
        _T_11317_17 <= _T_2167_17;
      end
    end
    if (reset) begin
      _T_11317_16 <= 5'h0;
    end else begin
      if (_T_11351) begin
        _T_11317_16 <= _T_2167_16;
      end
    end
    if (reset) begin
      _T_11317_15 <= 5'h0;
    end else begin
      if (_T_11335) begin
        _T_11317_15 <= _T_3447;
      end
    end
    if (reset) begin
      _T_11317_14 <= 4'h0;
    end else begin
      if (_T_11335) begin
        _T_11317_14 <= _T_2167_14;
      end
    end
    if (reset) begin
      _T_11317_13 <= 4'h0;
    end else begin
      if (_T_11335) begin
        _T_11317_13 <= _T_2167_13;
      end
    end
    if (reset) begin
      _T_11317_12 <= 4'h0;
    end else begin
      if (_T_11335) begin
        _T_11317_12 <= _T_2167_12;
      end
    end
    if (reset) begin
      _T_11317_11 <= 4'h0;
    end else begin
      if (_T_11335) begin
        _T_11317_11 <= _T_2167_11;
      end
    end
    if (reset) begin
      _T_11317_10 <= 4'h0;
    end else begin
      if (_T_11335) begin
        _T_11317_10 <= _T_2167_10;
      end
    end
    if (reset) begin
      _T_11317_9 <= 4'h0;
    end else begin
      if (_T_11335) begin
        _T_11317_9 <= _T_2167_9;
      end
    end
    if (reset) begin
      _T_11317_8 <= 4'h0;
    end else begin
      if (_T_11335) begin
        _T_11317_8 <= _T_2167_8;
      end
    end
    if (reset) begin
      _T_11317_7 <= 4'h0;
    end else begin
      if (_T_11319) begin
        _T_11317_7 <= _T_2743;
      end
    end
    if (reset) begin
      _T_11317_6 <= 3'h0;
    end else begin
      if (_T_11319) begin
        _T_11317_6 <= _T_2167_6;
      end
    end
    if (reset) begin
      _T_11317_5 <= 3'h0;
    end else begin
      if (_T_11319) begin
        _T_11317_5 <= _T_2167_5;
      end
    end
    if (reset) begin
      _T_11317_4 <= 3'h0;
    end else begin
      if (_T_11319) begin
        _T_11317_4 <= _T_2167_4;
      end
    end
    if (reset) begin
      _T_11317_3 <= 3'h0;
    end else begin
      if (_T_11319) begin
        _T_11317_3 <= _T_2439;
      end
    end
    if (reset) begin
      _T_11317_2 <= 2'h0;
    end else begin
      if (_T_11319) begin
        _T_11317_2 <= _T_2167_2;
      end
    end
    if (reset) begin
      _T_11317_1 <= 2'h0;
    end else begin
      if (_T_11319) begin
        _T_11317_1 <= _T_2299;
      end
    end
    if (reset) begin
      _T_11317_0 <= 1'h0;
    end else begin
      if (_T_11319) begin
        _T_11317_0 <= _T_2231;
      end
    end
    if (reset) begin
      _T_17822 <= 1'h0;
    end else begin
      _T_17822 <= _T_10362;
    end
    if (reset) begin
      _T_17961_0 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_0 <= _T_10641_0;
      end
    end
    if (reset) begin
      _T_17961_1 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_1 <= _T_10641_1;
      end
    end
    if (reset) begin
      _T_17961_2 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_2 <= _T_10641_2;
      end
    end
    if (reset) begin
      _T_17961_3 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_3 <= _T_10641_3;
      end
    end
    if (reset) begin
      _T_17961_4 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_4 <= _T_10641_4;
      end
    end
    if (reset) begin
      _T_17961_5 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_5 <= _T_10641_5;
      end
    end
    if (reset) begin
      _T_17961_6 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_6 <= _T_10641_6;
      end
    end
    if (reset) begin
      _T_17961_7 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_7 <= _T_10641_7;
      end
    end
    if (reset) begin
      _T_17961_8 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_8 <= _T_10641_8;
      end
    end
    if (reset) begin
      _T_17961_9 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_9 <= _T_10641_9;
      end
    end
    if (reset) begin
      _T_17961_10 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_10 <= _T_10641_10;
      end
    end
    if (reset) begin
      _T_17961_11 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_11 <= _T_10641_11;
      end
    end
    if (reset) begin
      _T_17961_12 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_12 <= _T_10641_12;
      end
    end
    if (reset) begin
      _T_17961_13 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_13 <= _T_10641_13;
      end
    end
    if (reset) begin
      _T_17961_14 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_14 <= _T_10641_14;
      end
    end
    if (reset) begin
      _T_17961_15 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_15 <= _T_10641_15;
      end
    end
    if (reset) begin
      _T_17961_16 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_16 <= _T_10641_16;
      end
    end
    if (reset) begin
      _T_17961_17 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_17 <= _T_10641_17;
      end
    end
    if (reset) begin
      _T_17961_18 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_18 <= _T_10641_18;
      end
    end
    if (reset) begin
      _T_17961_19 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_19 <= _T_10641_19;
      end
    end
    if (reset) begin
      _T_17961_20 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_20 <= _T_10641_20;
      end
    end
    if (reset) begin
      _T_17961_21 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_21 <= _T_10641_21;
      end
    end
    if (reset) begin
      _T_17961_22 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_22 <= _T_10641_22;
      end
    end
    if (reset) begin
      _T_17961_23 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_23 <= _T_10641_23;
      end
    end
    if (reset) begin
      _T_17961_24 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_24 <= _T_10641_24;
      end
    end
    if (reset) begin
      _T_17961_25 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_25 <= _T_10641_25;
      end
    end
    if (reset) begin
      _T_17961_26 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_26 <= _T_10641_26;
      end
    end
    if (reset) begin
      _T_17961_27 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_27 <= _T_10641_27;
      end
    end
    if (reset) begin
      _T_17961_28 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_28 <= _T_10641_28;
      end
    end
    if (reset) begin
      _T_17961_29 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_29 <= _T_10641_29;
      end
    end
    if (reset) begin
      _T_17961_30 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_30 <= _T_10641_30;
      end
    end
    if (reset) begin
      _T_17961_31 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_31 <= _T_10641_31;
      end
    end
    if (_T_10362) begin
      if (_T_10436_0) begin
        if (_T_11317_0) begin
          _T_18065_0 <= _T_10366_0;
        end else begin
          _T_18065_0 <= 8'h0;
        end
      end else begin
        _T_18065_0 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_1) begin
        if (_T_11525) begin
          _T_18065_1 <= _T_10366_0;
        end else begin
          if (_T_11523) begin
            _T_18065_1 <= _T_10366_1;
          end else begin
            _T_18065_1 <= 8'h0;
          end
        end
      end else begin
        _T_18065_1 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_2) begin
        if (_T_11535) begin
          _T_18065_2 <= _T_10366_0;
        end else begin
          if (_T_11533) begin
            _T_18065_2 <= _T_10366_1;
          end else begin
            if (_T_11531) begin
              _T_18065_2 <= _T_10366_2;
            end else begin
              _T_18065_2 <= 8'h0;
            end
          end
        end
      end else begin
        _T_18065_2 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_3) begin
        if (_T_11548) begin
          _T_18065_3 <= _T_10366_0;
        end else begin
          if (_T_11546) begin
            _T_18065_3 <= _T_10366_1;
          end else begin
            if (_T_11544) begin
              _T_18065_3 <= _T_10366_2;
            end else begin
              if (_T_11542) begin
                _T_18065_3 <= _T_10366_3;
              end else begin
                _T_18065_3 <= 8'h0;
              end
            end
          end
        end
      end else begin
        _T_18065_3 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_4) begin
        if (_T_11564) begin
          _T_18065_4 <= _T_10366_0;
        end else begin
          if (_T_11562) begin
            _T_18065_4 <= _T_10366_1;
          end else begin
            if (_T_11560) begin
              _T_18065_4 <= _T_10366_2;
            end else begin
              if (_T_11558) begin
                _T_18065_4 <= _T_10366_3;
              end else begin
                if (_T_11556) begin
                  _T_18065_4 <= _T_10366_4;
                end else begin
                  _T_18065_4 <= 8'h0;
                end
              end
            end
          end
        end
      end else begin
        _T_18065_4 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_5) begin
        if (_T_11583) begin
          _T_18065_5 <= _T_10366_0;
        end else begin
          if (_T_11581) begin
            _T_18065_5 <= _T_10366_1;
          end else begin
            if (_T_11579) begin
              _T_18065_5 <= _T_10366_2;
            end else begin
              if (_T_11577) begin
                _T_18065_5 <= _T_10366_3;
              end else begin
                if (_T_11575) begin
                  _T_18065_5 <= _T_10366_4;
                end else begin
                  if (_T_11573) begin
                    _T_18065_5 <= _T_10366_5;
                  end else begin
                    _T_18065_5 <= 8'h0;
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_5 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_6) begin
        if (_T_11605) begin
          _T_18065_6 <= _T_10366_0;
        end else begin
          if (_T_11603) begin
            _T_18065_6 <= _T_10366_1;
          end else begin
            if (_T_11601) begin
              _T_18065_6 <= _T_10366_2;
            end else begin
              if (_T_11599) begin
                _T_18065_6 <= _T_10366_3;
              end else begin
                if (_T_11597) begin
                  _T_18065_6 <= _T_10366_4;
                end else begin
                  if (_T_11595) begin
                    _T_18065_6 <= _T_10366_5;
                  end else begin
                    if (_T_11593) begin
                      _T_18065_6 <= _T_10366_6;
                    end else begin
                      _T_18065_6 <= 8'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_6 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_7) begin
        if (_T_11630) begin
          _T_18065_7 <= _T_10366_0;
        end else begin
          if (_T_11628) begin
            _T_18065_7 <= _T_10366_1;
          end else begin
            if (_T_11626) begin
              _T_18065_7 <= _T_10366_2;
            end else begin
              if (_T_11624) begin
                _T_18065_7 <= _T_10366_3;
              end else begin
                if (_T_11622) begin
                  _T_18065_7 <= _T_10366_4;
                end else begin
                  if (_T_11620) begin
                    _T_18065_7 <= _T_10366_5;
                  end else begin
                    if (_T_11618) begin
                      _T_18065_7 <= _T_10366_6;
                    end else begin
                      if (_T_11616) begin
                        _T_18065_7 <= _T_10366_7;
                      end else begin
                        _T_18065_7 <= 8'h0;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_7 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_8) begin
        if (_T_11658) begin
          _T_18065_8 <= _T_10366_0;
        end else begin
          if (_T_11656) begin
            _T_18065_8 <= _T_10366_1;
          end else begin
            if (_T_11654) begin
              _T_18065_8 <= _T_10366_2;
            end else begin
              if (_T_11652) begin
                _T_18065_8 <= _T_10366_3;
              end else begin
                if (_T_11650) begin
                  _T_18065_8 <= _T_10366_4;
                end else begin
                  if (_T_11648) begin
                    _T_18065_8 <= _T_10366_5;
                  end else begin
                    if (_T_11646) begin
                      _T_18065_8 <= _T_10366_6;
                    end else begin
                      if (_T_11644) begin
                        _T_18065_8 <= _T_10366_7;
                      end else begin
                        if (_T_11642) begin
                          _T_18065_8 <= _T_10366_8;
                        end else begin
                          _T_18065_8 <= 8'h0;
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_8 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_9) begin
        if (_T_11689) begin
          _T_18065_9 <= _T_10366_0;
        end else begin
          if (_T_11687) begin
            _T_18065_9 <= _T_10366_1;
          end else begin
            if (_T_11685) begin
              _T_18065_9 <= _T_10366_2;
            end else begin
              if (_T_11683) begin
                _T_18065_9 <= _T_10366_3;
              end else begin
                if (_T_11681) begin
                  _T_18065_9 <= _T_10366_4;
                end else begin
                  if (_T_11679) begin
                    _T_18065_9 <= _T_10366_5;
                  end else begin
                    if (_T_11677) begin
                      _T_18065_9 <= _T_10366_6;
                    end else begin
                      if (_T_11675) begin
                        _T_18065_9 <= _T_10366_7;
                      end else begin
                        if (_T_11673) begin
                          _T_18065_9 <= _T_10366_8;
                        end else begin
                          if (_T_11671) begin
                            _T_18065_9 <= _T_10366_9;
                          end else begin
                            _T_18065_9 <= 8'h0;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_9 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_10) begin
        if (_T_11723) begin
          _T_18065_10 <= _T_10366_0;
        end else begin
          if (_T_11721) begin
            _T_18065_10 <= _T_10366_1;
          end else begin
            if (_T_11719) begin
              _T_18065_10 <= _T_10366_2;
            end else begin
              if (_T_11717) begin
                _T_18065_10 <= _T_10366_3;
              end else begin
                if (_T_11715) begin
                  _T_18065_10 <= _T_10366_4;
                end else begin
                  if (_T_11713) begin
                    _T_18065_10 <= _T_10366_5;
                  end else begin
                    if (_T_11711) begin
                      _T_18065_10 <= _T_10366_6;
                    end else begin
                      if (_T_11709) begin
                        _T_18065_10 <= _T_10366_7;
                      end else begin
                        if (_T_11707) begin
                          _T_18065_10 <= _T_10366_8;
                        end else begin
                          if (_T_11705) begin
                            _T_18065_10 <= _T_10366_9;
                          end else begin
                            if (_T_11703) begin
                              _T_18065_10 <= _T_10366_10;
                            end else begin
                              _T_18065_10 <= 8'h0;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_10 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_11) begin
        if (_T_11760) begin
          _T_18065_11 <= _T_10366_0;
        end else begin
          if (_T_11758) begin
            _T_18065_11 <= _T_10366_1;
          end else begin
            if (_T_11756) begin
              _T_18065_11 <= _T_10366_2;
            end else begin
              if (_T_11754) begin
                _T_18065_11 <= _T_10366_3;
              end else begin
                if (_T_11752) begin
                  _T_18065_11 <= _T_10366_4;
                end else begin
                  if (_T_11750) begin
                    _T_18065_11 <= _T_10366_5;
                  end else begin
                    if (_T_11748) begin
                      _T_18065_11 <= _T_10366_6;
                    end else begin
                      if (_T_11746) begin
                        _T_18065_11 <= _T_10366_7;
                      end else begin
                        if (_T_11744) begin
                          _T_18065_11 <= _T_10366_8;
                        end else begin
                          if (_T_11742) begin
                            _T_18065_11 <= _T_10366_9;
                          end else begin
                            if (_T_11740) begin
                              _T_18065_11 <= _T_10366_10;
                            end else begin
                              if (_T_11738) begin
                                _T_18065_11 <= _T_10366_11;
                              end else begin
                                _T_18065_11 <= 8'h0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_11 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_12) begin
        if (_T_11800) begin
          _T_18065_12 <= _T_10366_0;
        end else begin
          if (_T_11798) begin
            _T_18065_12 <= _T_10366_1;
          end else begin
            if (_T_11796) begin
              _T_18065_12 <= _T_10366_2;
            end else begin
              if (_T_11794) begin
                _T_18065_12 <= _T_10366_3;
              end else begin
                if (_T_11792) begin
                  _T_18065_12 <= _T_10366_4;
                end else begin
                  if (_T_11790) begin
                    _T_18065_12 <= _T_10366_5;
                  end else begin
                    if (_T_11788) begin
                      _T_18065_12 <= _T_10366_6;
                    end else begin
                      if (_T_11786) begin
                        _T_18065_12 <= _T_10366_7;
                      end else begin
                        if (_T_11784) begin
                          _T_18065_12 <= _T_10366_8;
                        end else begin
                          if (_T_11782) begin
                            _T_18065_12 <= _T_10366_9;
                          end else begin
                            if (_T_11780) begin
                              _T_18065_12 <= _T_10366_10;
                            end else begin
                              if (_T_11778) begin
                                _T_18065_12 <= _T_10366_11;
                              end else begin
                                if (_T_11776) begin
                                  _T_18065_12 <= _T_10366_12;
                                end else begin
                                  _T_18065_12 <= 8'h0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_12 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_13) begin
        if (_T_11843) begin
          _T_18065_13 <= _T_10366_0;
        end else begin
          if (_T_11841) begin
            _T_18065_13 <= _T_10366_1;
          end else begin
            if (_T_11839) begin
              _T_18065_13 <= _T_10366_2;
            end else begin
              if (_T_11837) begin
                _T_18065_13 <= _T_10366_3;
              end else begin
                if (_T_11835) begin
                  _T_18065_13 <= _T_10366_4;
                end else begin
                  if (_T_11833) begin
                    _T_18065_13 <= _T_10366_5;
                  end else begin
                    if (_T_11831) begin
                      _T_18065_13 <= _T_10366_6;
                    end else begin
                      if (_T_11829) begin
                        _T_18065_13 <= _T_10366_7;
                      end else begin
                        if (_T_11827) begin
                          _T_18065_13 <= _T_10366_8;
                        end else begin
                          if (_T_11825) begin
                            _T_18065_13 <= _T_10366_9;
                          end else begin
                            if (_T_11823) begin
                              _T_18065_13 <= _T_10366_10;
                            end else begin
                              if (_T_11821) begin
                                _T_18065_13 <= _T_10366_11;
                              end else begin
                                if (_T_11819) begin
                                  _T_18065_13 <= _T_10366_12;
                                end else begin
                                  if (_T_11817) begin
                                    _T_18065_13 <= _T_10366_13;
                                  end else begin
                                    _T_18065_13 <= 8'h0;
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_13 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_14) begin
        if (_T_11889) begin
          _T_18065_14 <= _T_10366_0;
        end else begin
          if (_T_11887) begin
            _T_18065_14 <= _T_10366_1;
          end else begin
            if (_T_11885) begin
              _T_18065_14 <= _T_10366_2;
            end else begin
              if (_T_11883) begin
                _T_18065_14 <= _T_10366_3;
              end else begin
                if (_T_11881) begin
                  _T_18065_14 <= _T_10366_4;
                end else begin
                  if (_T_11879) begin
                    _T_18065_14 <= _T_10366_5;
                  end else begin
                    if (_T_11877) begin
                      _T_18065_14 <= _T_10366_6;
                    end else begin
                      if (_T_11875) begin
                        _T_18065_14 <= _T_10366_7;
                      end else begin
                        if (_T_11873) begin
                          _T_18065_14 <= _T_10366_8;
                        end else begin
                          if (_T_11871) begin
                            _T_18065_14 <= _T_10366_9;
                          end else begin
                            if (_T_11869) begin
                              _T_18065_14 <= _T_10366_10;
                            end else begin
                              if (_T_11867) begin
                                _T_18065_14 <= _T_10366_11;
                              end else begin
                                if (_T_11865) begin
                                  _T_18065_14 <= _T_10366_12;
                                end else begin
                                  if (_T_11863) begin
                                    _T_18065_14 <= _T_10366_13;
                                  end else begin
                                    if (_T_11861) begin
                                      _T_18065_14 <= _T_10366_14;
                                    end else begin
                                      _T_18065_14 <= 8'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_14 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_15) begin
        if (_T_11938) begin
          _T_18065_15 <= _T_10366_0;
        end else begin
          if (_T_11936) begin
            _T_18065_15 <= _T_10366_1;
          end else begin
            if (_T_11934) begin
              _T_18065_15 <= _T_10366_2;
            end else begin
              if (_T_11932) begin
                _T_18065_15 <= _T_10366_3;
              end else begin
                if (_T_11930) begin
                  _T_18065_15 <= _T_10366_4;
                end else begin
                  if (_T_11928) begin
                    _T_18065_15 <= _T_10366_5;
                  end else begin
                    if (_T_11926) begin
                      _T_18065_15 <= _T_10366_6;
                    end else begin
                      if (_T_11924) begin
                        _T_18065_15 <= _T_10366_7;
                      end else begin
                        if (_T_11922) begin
                          _T_18065_15 <= _T_10366_8;
                        end else begin
                          if (_T_11920) begin
                            _T_18065_15 <= _T_10366_9;
                          end else begin
                            if (_T_11918) begin
                              _T_18065_15 <= _T_10366_10;
                            end else begin
                              if (_T_11916) begin
                                _T_18065_15 <= _T_10366_11;
                              end else begin
                                if (_T_11914) begin
                                  _T_18065_15 <= _T_10366_12;
                                end else begin
                                  if (_T_11912) begin
                                    _T_18065_15 <= _T_10366_13;
                                  end else begin
                                    if (_T_11910) begin
                                      _T_18065_15 <= _T_10366_14;
                                    end else begin
                                      if (_T_11908) begin
                                        _T_18065_15 <= _T_10366_15;
                                      end else begin
                                        _T_18065_15 <= 8'h0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_15 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_16) begin
        if (_T_11990) begin
          _T_18065_16 <= _T_10366_0;
        end else begin
          if (_T_11988) begin
            _T_18065_16 <= _T_10366_1;
          end else begin
            if (_T_11986) begin
              _T_18065_16 <= _T_10366_2;
            end else begin
              if (_T_11984) begin
                _T_18065_16 <= _T_10366_3;
              end else begin
                if (_T_11982) begin
                  _T_18065_16 <= _T_10366_4;
                end else begin
                  if (_T_11980) begin
                    _T_18065_16 <= _T_10366_5;
                  end else begin
                    if (_T_11978) begin
                      _T_18065_16 <= _T_10366_6;
                    end else begin
                      if (_T_11976) begin
                        _T_18065_16 <= _T_10366_7;
                      end else begin
                        if (_T_11974) begin
                          _T_18065_16 <= _T_10366_8;
                        end else begin
                          if (_T_11972) begin
                            _T_18065_16 <= _T_10366_9;
                          end else begin
                            if (_T_11970) begin
                              _T_18065_16 <= _T_10366_10;
                            end else begin
                              if (_T_11968) begin
                                _T_18065_16 <= _T_10366_11;
                              end else begin
                                if (_T_11966) begin
                                  _T_18065_16 <= _T_10366_12;
                                end else begin
                                  if (_T_11964) begin
                                    _T_18065_16 <= _T_10366_13;
                                  end else begin
                                    if (_T_11962) begin
                                      _T_18065_16 <= _T_10366_14;
                                    end else begin
                                      if (_T_11960) begin
                                        _T_18065_16 <= _T_10366_15;
                                      end else begin
                                        if (_T_11958) begin
                                          _T_18065_16 <= _T_10366_16;
                                        end else begin
                                          _T_18065_16 <= 8'h0;
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_16 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_17) begin
        if (_T_12045) begin
          _T_18065_17 <= _T_10366_0;
        end else begin
          if (_T_12043) begin
            _T_18065_17 <= _T_10366_1;
          end else begin
            if (_T_12041) begin
              _T_18065_17 <= _T_10366_2;
            end else begin
              if (_T_12039) begin
                _T_18065_17 <= _T_10366_3;
              end else begin
                if (_T_12037) begin
                  _T_18065_17 <= _T_10366_4;
                end else begin
                  if (_T_12035) begin
                    _T_18065_17 <= _T_10366_5;
                  end else begin
                    if (_T_12033) begin
                      _T_18065_17 <= _T_10366_6;
                    end else begin
                      if (_T_12031) begin
                        _T_18065_17 <= _T_10366_7;
                      end else begin
                        if (_T_12029) begin
                          _T_18065_17 <= _T_10366_8;
                        end else begin
                          if (_T_12027) begin
                            _T_18065_17 <= _T_10366_9;
                          end else begin
                            if (_T_12025) begin
                              _T_18065_17 <= _T_10366_10;
                            end else begin
                              if (_T_12023) begin
                                _T_18065_17 <= _T_10366_11;
                              end else begin
                                if (_T_12021) begin
                                  _T_18065_17 <= _T_10366_12;
                                end else begin
                                  if (_T_12019) begin
                                    _T_18065_17 <= _T_10366_13;
                                  end else begin
                                    if (_T_12017) begin
                                      _T_18065_17 <= _T_10366_14;
                                    end else begin
                                      if (_T_12015) begin
                                        _T_18065_17 <= _T_10366_15;
                                      end else begin
                                        if (_T_12013) begin
                                          _T_18065_17 <= _T_10366_16;
                                        end else begin
                                          if (_T_12011) begin
                                            _T_18065_17 <= _T_10366_17;
                                          end else begin
                                            _T_18065_17 <= 8'h0;
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_17 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_18) begin
        if (_T_12103) begin
          _T_18065_18 <= _T_10366_0;
        end else begin
          if (_T_12101) begin
            _T_18065_18 <= _T_10366_1;
          end else begin
            if (_T_12099) begin
              _T_18065_18 <= _T_10366_2;
            end else begin
              if (_T_12097) begin
                _T_18065_18 <= _T_10366_3;
              end else begin
                if (_T_12095) begin
                  _T_18065_18 <= _T_10366_4;
                end else begin
                  if (_T_12093) begin
                    _T_18065_18 <= _T_10366_5;
                  end else begin
                    if (_T_12091) begin
                      _T_18065_18 <= _T_10366_6;
                    end else begin
                      if (_T_12089) begin
                        _T_18065_18 <= _T_10366_7;
                      end else begin
                        if (_T_12087) begin
                          _T_18065_18 <= _T_10366_8;
                        end else begin
                          if (_T_12085) begin
                            _T_18065_18 <= _T_10366_9;
                          end else begin
                            if (_T_12083) begin
                              _T_18065_18 <= _T_10366_10;
                            end else begin
                              if (_T_12081) begin
                                _T_18065_18 <= _T_10366_11;
                              end else begin
                                if (_T_12079) begin
                                  _T_18065_18 <= _T_10366_12;
                                end else begin
                                  if (_T_12077) begin
                                    _T_18065_18 <= _T_10366_13;
                                  end else begin
                                    if (_T_12075) begin
                                      _T_18065_18 <= _T_10366_14;
                                    end else begin
                                      if (_T_12073) begin
                                        _T_18065_18 <= _T_10366_15;
                                      end else begin
                                        if (_T_12071) begin
                                          _T_18065_18 <= _T_10366_16;
                                        end else begin
                                          if (_T_12069) begin
                                            _T_18065_18 <= _T_10366_17;
                                          end else begin
                                            if (_T_12067) begin
                                              _T_18065_18 <= _T_10366_18;
                                            end else begin
                                              _T_18065_18 <= 8'h0;
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_18 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_19) begin
        if (_T_12164) begin
          _T_18065_19 <= _T_10366_0;
        end else begin
          if (_T_12162) begin
            _T_18065_19 <= _T_10366_1;
          end else begin
            if (_T_12160) begin
              _T_18065_19 <= _T_10366_2;
            end else begin
              if (_T_12158) begin
                _T_18065_19 <= _T_10366_3;
              end else begin
                if (_T_12156) begin
                  _T_18065_19 <= _T_10366_4;
                end else begin
                  if (_T_12154) begin
                    _T_18065_19 <= _T_10366_5;
                  end else begin
                    if (_T_12152) begin
                      _T_18065_19 <= _T_10366_6;
                    end else begin
                      if (_T_12150) begin
                        _T_18065_19 <= _T_10366_7;
                      end else begin
                        if (_T_12148) begin
                          _T_18065_19 <= _T_10366_8;
                        end else begin
                          if (_T_12146) begin
                            _T_18065_19 <= _T_10366_9;
                          end else begin
                            if (_T_12144) begin
                              _T_18065_19 <= _T_10366_10;
                            end else begin
                              if (_T_12142) begin
                                _T_18065_19 <= _T_10366_11;
                              end else begin
                                if (_T_12140) begin
                                  _T_18065_19 <= _T_10366_12;
                                end else begin
                                  if (_T_12138) begin
                                    _T_18065_19 <= _T_10366_13;
                                  end else begin
                                    if (_T_12136) begin
                                      _T_18065_19 <= _T_10366_14;
                                    end else begin
                                      if (_T_12134) begin
                                        _T_18065_19 <= _T_10366_15;
                                      end else begin
                                        if (_T_12132) begin
                                          _T_18065_19 <= _T_10366_16;
                                        end else begin
                                          if (_T_12130) begin
                                            _T_18065_19 <= _T_10366_17;
                                          end else begin
                                            if (_T_12128) begin
                                              _T_18065_19 <= _T_10366_18;
                                            end else begin
                                              if (_T_12126) begin
                                                _T_18065_19 <= _T_10366_19;
                                              end else begin
                                                _T_18065_19 <= 8'h0;
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_19 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_20) begin
        if (_T_12228) begin
          _T_18065_20 <= _T_10366_0;
        end else begin
          if (_T_12226) begin
            _T_18065_20 <= _T_10366_1;
          end else begin
            if (_T_12224) begin
              _T_18065_20 <= _T_10366_2;
            end else begin
              if (_T_12222) begin
                _T_18065_20 <= _T_10366_3;
              end else begin
                if (_T_12220) begin
                  _T_18065_20 <= _T_10366_4;
                end else begin
                  if (_T_12218) begin
                    _T_18065_20 <= _T_10366_5;
                  end else begin
                    if (_T_12216) begin
                      _T_18065_20 <= _T_10366_6;
                    end else begin
                      if (_T_12214) begin
                        _T_18065_20 <= _T_10366_7;
                      end else begin
                        if (_T_12212) begin
                          _T_18065_20 <= _T_10366_8;
                        end else begin
                          if (_T_12210) begin
                            _T_18065_20 <= _T_10366_9;
                          end else begin
                            if (_T_12208) begin
                              _T_18065_20 <= _T_10366_10;
                            end else begin
                              if (_T_12206) begin
                                _T_18065_20 <= _T_10366_11;
                              end else begin
                                if (_T_12204) begin
                                  _T_18065_20 <= _T_10366_12;
                                end else begin
                                  if (_T_12202) begin
                                    _T_18065_20 <= _T_10366_13;
                                  end else begin
                                    if (_T_12200) begin
                                      _T_18065_20 <= _T_10366_14;
                                    end else begin
                                      if (_T_12198) begin
                                        _T_18065_20 <= _T_10366_15;
                                      end else begin
                                        if (_T_12196) begin
                                          _T_18065_20 <= _T_10366_16;
                                        end else begin
                                          if (_T_12194) begin
                                            _T_18065_20 <= _T_10366_17;
                                          end else begin
                                            if (_T_12192) begin
                                              _T_18065_20 <= _T_10366_18;
                                            end else begin
                                              if (_T_12190) begin
                                                _T_18065_20 <= _T_10366_19;
                                              end else begin
                                                if (_T_12188) begin
                                                  _T_18065_20 <= _T_10366_20;
                                                end else begin
                                                  _T_18065_20 <= 8'h0;
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_20 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_21) begin
        if (_T_12295) begin
          _T_18065_21 <= _T_10366_0;
        end else begin
          if (_T_12293) begin
            _T_18065_21 <= _T_10366_1;
          end else begin
            if (_T_12291) begin
              _T_18065_21 <= _T_10366_2;
            end else begin
              if (_T_12289) begin
                _T_18065_21 <= _T_10366_3;
              end else begin
                if (_T_12287) begin
                  _T_18065_21 <= _T_10366_4;
                end else begin
                  if (_T_12285) begin
                    _T_18065_21 <= _T_10366_5;
                  end else begin
                    if (_T_12283) begin
                      _T_18065_21 <= _T_10366_6;
                    end else begin
                      if (_T_12281) begin
                        _T_18065_21 <= _T_10366_7;
                      end else begin
                        if (_T_12279) begin
                          _T_18065_21 <= _T_10366_8;
                        end else begin
                          if (_T_12277) begin
                            _T_18065_21 <= _T_10366_9;
                          end else begin
                            if (_T_12275) begin
                              _T_18065_21 <= _T_10366_10;
                            end else begin
                              if (_T_12273) begin
                                _T_18065_21 <= _T_10366_11;
                              end else begin
                                if (_T_12271) begin
                                  _T_18065_21 <= _T_10366_12;
                                end else begin
                                  if (_T_12269) begin
                                    _T_18065_21 <= _T_10366_13;
                                  end else begin
                                    if (_T_12267) begin
                                      _T_18065_21 <= _T_10366_14;
                                    end else begin
                                      if (_T_12265) begin
                                        _T_18065_21 <= _T_10366_15;
                                      end else begin
                                        if (_T_12263) begin
                                          _T_18065_21 <= _T_10366_16;
                                        end else begin
                                          if (_T_12261) begin
                                            _T_18065_21 <= _T_10366_17;
                                          end else begin
                                            if (_T_12259) begin
                                              _T_18065_21 <= _T_10366_18;
                                            end else begin
                                              if (_T_12257) begin
                                                _T_18065_21 <= _T_10366_19;
                                              end else begin
                                                if (_T_12255) begin
                                                  _T_18065_21 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12253) begin
                                                    _T_18065_21 <= _T_10366_21;
                                                  end else begin
                                                    _T_18065_21 <= 8'h0;
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_21 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_22) begin
        if (_T_12365) begin
          _T_18065_22 <= _T_10366_0;
        end else begin
          if (_T_12363) begin
            _T_18065_22 <= _T_10366_1;
          end else begin
            if (_T_12361) begin
              _T_18065_22 <= _T_10366_2;
            end else begin
              if (_T_12359) begin
                _T_18065_22 <= _T_10366_3;
              end else begin
                if (_T_12357) begin
                  _T_18065_22 <= _T_10366_4;
                end else begin
                  if (_T_12355) begin
                    _T_18065_22 <= _T_10366_5;
                  end else begin
                    if (_T_12353) begin
                      _T_18065_22 <= _T_10366_6;
                    end else begin
                      if (_T_12351) begin
                        _T_18065_22 <= _T_10366_7;
                      end else begin
                        if (_T_12349) begin
                          _T_18065_22 <= _T_10366_8;
                        end else begin
                          if (_T_12347) begin
                            _T_18065_22 <= _T_10366_9;
                          end else begin
                            if (_T_12345) begin
                              _T_18065_22 <= _T_10366_10;
                            end else begin
                              if (_T_12343) begin
                                _T_18065_22 <= _T_10366_11;
                              end else begin
                                if (_T_12341) begin
                                  _T_18065_22 <= _T_10366_12;
                                end else begin
                                  if (_T_12339) begin
                                    _T_18065_22 <= _T_10366_13;
                                  end else begin
                                    if (_T_12337) begin
                                      _T_18065_22 <= _T_10366_14;
                                    end else begin
                                      if (_T_12335) begin
                                        _T_18065_22 <= _T_10366_15;
                                      end else begin
                                        if (_T_12333) begin
                                          _T_18065_22 <= _T_10366_16;
                                        end else begin
                                          if (_T_12331) begin
                                            _T_18065_22 <= _T_10366_17;
                                          end else begin
                                            if (_T_12329) begin
                                              _T_18065_22 <= _T_10366_18;
                                            end else begin
                                              if (_T_12327) begin
                                                _T_18065_22 <= _T_10366_19;
                                              end else begin
                                                if (_T_12325) begin
                                                  _T_18065_22 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12323) begin
                                                    _T_18065_22 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12321) begin
                                                      _T_18065_22 <= _T_10366_22;
                                                    end else begin
                                                      _T_18065_22 <= 8'h0;
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_22 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_23) begin
        if (_T_12438) begin
          _T_18065_23 <= _T_10366_0;
        end else begin
          if (_T_12436) begin
            _T_18065_23 <= _T_10366_1;
          end else begin
            if (_T_12434) begin
              _T_18065_23 <= _T_10366_2;
            end else begin
              if (_T_12432) begin
                _T_18065_23 <= _T_10366_3;
              end else begin
                if (_T_12430) begin
                  _T_18065_23 <= _T_10366_4;
                end else begin
                  if (_T_12428) begin
                    _T_18065_23 <= _T_10366_5;
                  end else begin
                    if (_T_12426) begin
                      _T_18065_23 <= _T_10366_6;
                    end else begin
                      if (_T_12424) begin
                        _T_18065_23 <= _T_10366_7;
                      end else begin
                        if (_T_12422) begin
                          _T_18065_23 <= _T_10366_8;
                        end else begin
                          if (_T_12420) begin
                            _T_18065_23 <= _T_10366_9;
                          end else begin
                            if (_T_12418) begin
                              _T_18065_23 <= _T_10366_10;
                            end else begin
                              if (_T_12416) begin
                                _T_18065_23 <= _T_10366_11;
                              end else begin
                                if (_T_12414) begin
                                  _T_18065_23 <= _T_10366_12;
                                end else begin
                                  if (_T_12412) begin
                                    _T_18065_23 <= _T_10366_13;
                                  end else begin
                                    if (_T_12410) begin
                                      _T_18065_23 <= _T_10366_14;
                                    end else begin
                                      if (_T_12408) begin
                                        _T_18065_23 <= _T_10366_15;
                                      end else begin
                                        if (_T_12406) begin
                                          _T_18065_23 <= _T_10366_16;
                                        end else begin
                                          if (_T_12404) begin
                                            _T_18065_23 <= _T_10366_17;
                                          end else begin
                                            if (_T_12402) begin
                                              _T_18065_23 <= _T_10366_18;
                                            end else begin
                                              if (_T_12400) begin
                                                _T_18065_23 <= _T_10366_19;
                                              end else begin
                                                if (_T_12398) begin
                                                  _T_18065_23 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12396) begin
                                                    _T_18065_23 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12394) begin
                                                      _T_18065_23 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_12392) begin
                                                        _T_18065_23 <= _T_10366_23;
                                                      end else begin
                                                        _T_18065_23 <= 8'h0;
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_23 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_24) begin
        if (_T_12514) begin
          _T_18065_24 <= _T_10366_0;
        end else begin
          if (_T_12512) begin
            _T_18065_24 <= _T_10366_1;
          end else begin
            if (_T_12510) begin
              _T_18065_24 <= _T_10366_2;
            end else begin
              if (_T_12508) begin
                _T_18065_24 <= _T_10366_3;
              end else begin
                if (_T_12506) begin
                  _T_18065_24 <= _T_10366_4;
                end else begin
                  if (_T_12504) begin
                    _T_18065_24 <= _T_10366_5;
                  end else begin
                    if (_T_12502) begin
                      _T_18065_24 <= _T_10366_6;
                    end else begin
                      if (_T_12500) begin
                        _T_18065_24 <= _T_10366_7;
                      end else begin
                        if (_T_12498) begin
                          _T_18065_24 <= _T_10366_8;
                        end else begin
                          if (_T_12496) begin
                            _T_18065_24 <= _T_10366_9;
                          end else begin
                            if (_T_12494) begin
                              _T_18065_24 <= _T_10366_10;
                            end else begin
                              if (_T_12492) begin
                                _T_18065_24 <= _T_10366_11;
                              end else begin
                                if (_T_12490) begin
                                  _T_18065_24 <= _T_10366_12;
                                end else begin
                                  if (_T_12488) begin
                                    _T_18065_24 <= _T_10366_13;
                                  end else begin
                                    if (_T_12486) begin
                                      _T_18065_24 <= _T_10366_14;
                                    end else begin
                                      if (_T_12484) begin
                                        _T_18065_24 <= _T_10366_15;
                                      end else begin
                                        if (_T_12482) begin
                                          _T_18065_24 <= _T_10366_16;
                                        end else begin
                                          if (_T_12480) begin
                                            _T_18065_24 <= _T_10366_17;
                                          end else begin
                                            if (_T_12478) begin
                                              _T_18065_24 <= _T_10366_18;
                                            end else begin
                                              if (_T_12476) begin
                                                _T_18065_24 <= _T_10366_19;
                                              end else begin
                                                if (_T_12474) begin
                                                  _T_18065_24 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12472) begin
                                                    _T_18065_24 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12470) begin
                                                      _T_18065_24 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_12468) begin
                                                        _T_18065_24 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_12466) begin
                                                          _T_18065_24 <= _T_10366_24;
                                                        end else begin
                                                          _T_18065_24 <= 8'h0;
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_24 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_25) begin
        if (_T_12593) begin
          _T_18065_25 <= _T_10366_0;
        end else begin
          if (_T_12591) begin
            _T_18065_25 <= _T_10366_1;
          end else begin
            if (_T_12589) begin
              _T_18065_25 <= _T_10366_2;
            end else begin
              if (_T_12587) begin
                _T_18065_25 <= _T_10366_3;
              end else begin
                if (_T_12585) begin
                  _T_18065_25 <= _T_10366_4;
                end else begin
                  if (_T_12583) begin
                    _T_18065_25 <= _T_10366_5;
                  end else begin
                    if (_T_12581) begin
                      _T_18065_25 <= _T_10366_6;
                    end else begin
                      if (_T_12579) begin
                        _T_18065_25 <= _T_10366_7;
                      end else begin
                        if (_T_12577) begin
                          _T_18065_25 <= _T_10366_8;
                        end else begin
                          if (_T_12575) begin
                            _T_18065_25 <= _T_10366_9;
                          end else begin
                            if (_T_12573) begin
                              _T_18065_25 <= _T_10366_10;
                            end else begin
                              if (_T_12571) begin
                                _T_18065_25 <= _T_10366_11;
                              end else begin
                                if (_T_12569) begin
                                  _T_18065_25 <= _T_10366_12;
                                end else begin
                                  if (_T_12567) begin
                                    _T_18065_25 <= _T_10366_13;
                                  end else begin
                                    if (_T_12565) begin
                                      _T_18065_25 <= _T_10366_14;
                                    end else begin
                                      if (_T_12563) begin
                                        _T_18065_25 <= _T_10366_15;
                                      end else begin
                                        if (_T_12561) begin
                                          _T_18065_25 <= _T_10366_16;
                                        end else begin
                                          if (_T_12559) begin
                                            _T_18065_25 <= _T_10366_17;
                                          end else begin
                                            if (_T_12557) begin
                                              _T_18065_25 <= _T_10366_18;
                                            end else begin
                                              if (_T_12555) begin
                                                _T_18065_25 <= _T_10366_19;
                                              end else begin
                                                if (_T_12553) begin
                                                  _T_18065_25 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12551) begin
                                                    _T_18065_25 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12549) begin
                                                      _T_18065_25 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_12547) begin
                                                        _T_18065_25 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_12545) begin
                                                          _T_18065_25 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_12543) begin
                                                            _T_18065_25 <= _T_10366_25;
                                                          end else begin
                                                            _T_18065_25 <= 8'h0;
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_25 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_26) begin
        if (_T_12675) begin
          _T_18065_26 <= _T_10366_0;
        end else begin
          if (_T_12673) begin
            _T_18065_26 <= _T_10366_1;
          end else begin
            if (_T_12671) begin
              _T_18065_26 <= _T_10366_2;
            end else begin
              if (_T_12669) begin
                _T_18065_26 <= _T_10366_3;
              end else begin
                if (_T_12667) begin
                  _T_18065_26 <= _T_10366_4;
                end else begin
                  if (_T_12665) begin
                    _T_18065_26 <= _T_10366_5;
                  end else begin
                    if (_T_12663) begin
                      _T_18065_26 <= _T_10366_6;
                    end else begin
                      if (_T_12661) begin
                        _T_18065_26 <= _T_10366_7;
                      end else begin
                        if (_T_12659) begin
                          _T_18065_26 <= _T_10366_8;
                        end else begin
                          if (_T_12657) begin
                            _T_18065_26 <= _T_10366_9;
                          end else begin
                            if (_T_12655) begin
                              _T_18065_26 <= _T_10366_10;
                            end else begin
                              if (_T_12653) begin
                                _T_18065_26 <= _T_10366_11;
                              end else begin
                                if (_T_12651) begin
                                  _T_18065_26 <= _T_10366_12;
                                end else begin
                                  if (_T_12649) begin
                                    _T_18065_26 <= _T_10366_13;
                                  end else begin
                                    if (_T_12647) begin
                                      _T_18065_26 <= _T_10366_14;
                                    end else begin
                                      if (_T_12645) begin
                                        _T_18065_26 <= _T_10366_15;
                                      end else begin
                                        if (_T_12643) begin
                                          _T_18065_26 <= _T_10366_16;
                                        end else begin
                                          if (_T_12641) begin
                                            _T_18065_26 <= _T_10366_17;
                                          end else begin
                                            if (_T_12639) begin
                                              _T_18065_26 <= _T_10366_18;
                                            end else begin
                                              if (_T_12637) begin
                                                _T_18065_26 <= _T_10366_19;
                                              end else begin
                                                if (_T_12635) begin
                                                  _T_18065_26 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12633) begin
                                                    _T_18065_26 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12631) begin
                                                      _T_18065_26 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_12629) begin
                                                        _T_18065_26 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_12627) begin
                                                          _T_18065_26 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_12625) begin
                                                            _T_18065_26 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_12623) begin
                                                              _T_18065_26 <= _T_10366_26;
                                                            end else begin
                                                              _T_18065_26 <= 8'h0;
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_26 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_27) begin
        if (_T_12760) begin
          _T_18065_27 <= _T_10366_0;
        end else begin
          if (_T_12758) begin
            _T_18065_27 <= _T_10366_1;
          end else begin
            if (_T_12756) begin
              _T_18065_27 <= _T_10366_2;
            end else begin
              if (_T_12754) begin
                _T_18065_27 <= _T_10366_3;
              end else begin
                if (_T_12752) begin
                  _T_18065_27 <= _T_10366_4;
                end else begin
                  if (_T_12750) begin
                    _T_18065_27 <= _T_10366_5;
                  end else begin
                    if (_T_12748) begin
                      _T_18065_27 <= _T_10366_6;
                    end else begin
                      if (_T_12746) begin
                        _T_18065_27 <= _T_10366_7;
                      end else begin
                        if (_T_12744) begin
                          _T_18065_27 <= _T_10366_8;
                        end else begin
                          if (_T_12742) begin
                            _T_18065_27 <= _T_10366_9;
                          end else begin
                            if (_T_12740) begin
                              _T_18065_27 <= _T_10366_10;
                            end else begin
                              if (_T_12738) begin
                                _T_18065_27 <= _T_10366_11;
                              end else begin
                                if (_T_12736) begin
                                  _T_18065_27 <= _T_10366_12;
                                end else begin
                                  if (_T_12734) begin
                                    _T_18065_27 <= _T_10366_13;
                                  end else begin
                                    if (_T_12732) begin
                                      _T_18065_27 <= _T_10366_14;
                                    end else begin
                                      if (_T_12730) begin
                                        _T_18065_27 <= _T_10366_15;
                                      end else begin
                                        if (_T_12728) begin
                                          _T_18065_27 <= _T_10366_16;
                                        end else begin
                                          if (_T_12726) begin
                                            _T_18065_27 <= _T_10366_17;
                                          end else begin
                                            if (_T_12724) begin
                                              _T_18065_27 <= _T_10366_18;
                                            end else begin
                                              if (_T_12722) begin
                                                _T_18065_27 <= _T_10366_19;
                                              end else begin
                                                if (_T_12720) begin
                                                  _T_18065_27 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12718) begin
                                                    _T_18065_27 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12716) begin
                                                      _T_18065_27 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_12714) begin
                                                        _T_18065_27 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_12712) begin
                                                          _T_18065_27 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_12710) begin
                                                            _T_18065_27 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_12708) begin
                                                              _T_18065_27 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_12706) begin
                                                                _T_18065_27 <= _T_10366_27;
                                                              end else begin
                                                                _T_18065_27 <= 8'h0;
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_27 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_28) begin
        if (_T_12848) begin
          _T_18065_28 <= _T_10366_0;
        end else begin
          if (_T_12846) begin
            _T_18065_28 <= _T_10366_1;
          end else begin
            if (_T_12844) begin
              _T_18065_28 <= _T_10366_2;
            end else begin
              if (_T_12842) begin
                _T_18065_28 <= _T_10366_3;
              end else begin
                if (_T_12840) begin
                  _T_18065_28 <= _T_10366_4;
                end else begin
                  if (_T_12838) begin
                    _T_18065_28 <= _T_10366_5;
                  end else begin
                    if (_T_12836) begin
                      _T_18065_28 <= _T_10366_6;
                    end else begin
                      if (_T_12834) begin
                        _T_18065_28 <= _T_10366_7;
                      end else begin
                        if (_T_12832) begin
                          _T_18065_28 <= _T_10366_8;
                        end else begin
                          if (_T_12830) begin
                            _T_18065_28 <= _T_10366_9;
                          end else begin
                            if (_T_12828) begin
                              _T_18065_28 <= _T_10366_10;
                            end else begin
                              if (_T_12826) begin
                                _T_18065_28 <= _T_10366_11;
                              end else begin
                                if (_T_12824) begin
                                  _T_18065_28 <= _T_10366_12;
                                end else begin
                                  if (_T_12822) begin
                                    _T_18065_28 <= _T_10366_13;
                                  end else begin
                                    if (_T_12820) begin
                                      _T_18065_28 <= _T_10366_14;
                                    end else begin
                                      if (_T_12818) begin
                                        _T_18065_28 <= _T_10366_15;
                                      end else begin
                                        if (_T_12816) begin
                                          _T_18065_28 <= _T_10366_16;
                                        end else begin
                                          if (_T_12814) begin
                                            _T_18065_28 <= _T_10366_17;
                                          end else begin
                                            if (_T_12812) begin
                                              _T_18065_28 <= _T_10366_18;
                                            end else begin
                                              if (_T_12810) begin
                                                _T_18065_28 <= _T_10366_19;
                                              end else begin
                                                if (_T_12808) begin
                                                  _T_18065_28 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12806) begin
                                                    _T_18065_28 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12804) begin
                                                      _T_18065_28 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_12802) begin
                                                        _T_18065_28 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_12800) begin
                                                          _T_18065_28 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_12798) begin
                                                            _T_18065_28 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_12796) begin
                                                              _T_18065_28 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_12794) begin
                                                                _T_18065_28 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_12792) begin
                                                                  _T_18065_28 <= _T_10366_28;
                                                                end else begin
                                                                  _T_18065_28 <= 8'h0;
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_28 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_29) begin
        if (_T_12939) begin
          _T_18065_29 <= _T_10366_0;
        end else begin
          if (_T_12937) begin
            _T_18065_29 <= _T_10366_1;
          end else begin
            if (_T_12935) begin
              _T_18065_29 <= _T_10366_2;
            end else begin
              if (_T_12933) begin
                _T_18065_29 <= _T_10366_3;
              end else begin
                if (_T_12931) begin
                  _T_18065_29 <= _T_10366_4;
                end else begin
                  if (_T_12929) begin
                    _T_18065_29 <= _T_10366_5;
                  end else begin
                    if (_T_12927) begin
                      _T_18065_29 <= _T_10366_6;
                    end else begin
                      if (_T_12925) begin
                        _T_18065_29 <= _T_10366_7;
                      end else begin
                        if (_T_12923) begin
                          _T_18065_29 <= _T_10366_8;
                        end else begin
                          if (_T_12921) begin
                            _T_18065_29 <= _T_10366_9;
                          end else begin
                            if (_T_12919) begin
                              _T_18065_29 <= _T_10366_10;
                            end else begin
                              if (_T_12917) begin
                                _T_18065_29 <= _T_10366_11;
                              end else begin
                                if (_T_12915) begin
                                  _T_18065_29 <= _T_10366_12;
                                end else begin
                                  if (_T_12913) begin
                                    _T_18065_29 <= _T_10366_13;
                                  end else begin
                                    if (_T_12911) begin
                                      _T_18065_29 <= _T_10366_14;
                                    end else begin
                                      if (_T_12909) begin
                                        _T_18065_29 <= _T_10366_15;
                                      end else begin
                                        if (_T_12907) begin
                                          _T_18065_29 <= _T_10366_16;
                                        end else begin
                                          if (_T_12905) begin
                                            _T_18065_29 <= _T_10366_17;
                                          end else begin
                                            if (_T_12903) begin
                                              _T_18065_29 <= _T_10366_18;
                                            end else begin
                                              if (_T_12901) begin
                                                _T_18065_29 <= _T_10366_19;
                                              end else begin
                                                if (_T_12899) begin
                                                  _T_18065_29 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12897) begin
                                                    _T_18065_29 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12895) begin
                                                      _T_18065_29 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_12893) begin
                                                        _T_18065_29 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_12891) begin
                                                          _T_18065_29 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_12889) begin
                                                            _T_18065_29 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_12887) begin
                                                              _T_18065_29 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_12885) begin
                                                                _T_18065_29 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_12883) begin
                                                                  _T_18065_29 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_12881) begin
                                                                    _T_18065_29 <= _T_10366_29;
                                                                  end else begin
                                                                    _T_18065_29 <= 8'h0;
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_29 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_30) begin
        if (_T_13033) begin
          _T_18065_30 <= _T_10366_0;
        end else begin
          if (_T_13031) begin
            _T_18065_30 <= _T_10366_1;
          end else begin
            if (_T_13029) begin
              _T_18065_30 <= _T_10366_2;
            end else begin
              if (_T_13027) begin
                _T_18065_30 <= _T_10366_3;
              end else begin
                if (_T_13025) begin
                  _T_18065_30 <= _T_10366_4;
                end else begin
                  if (_T_13023) begin
                    _T_18065_30 <= _T_10366_5;
                  end else begin
                    if (_T_13021) begin
                      _T_18065_30 <= _T_10366_6;
                    end else begin
                      if (_T_13019) begin
                        _T_18065_30 <= _T_10366_7;
                      end else begin
                        if (_T_13017) begin
                          _T_18065_30 <= _T_10366_8;
                        end else begin
                          if (_T_13015) begin
                            _T_18065_30 <= _T_10366_9;
                          end else begin
                            if (_T_13013) begin
                              _T_18065_30 <= _T_10366_10;
                            end else begin
                              if (_T_13011) begin
                                _T_18065_30 <= _T_10366_11;
                              end else begin
                                if (_T_13009) begin
                                  _T_18065_30 <= _T_10366_12;
                                end else begin
                                  if (_T_13007) begin
                                    _T_18065_30 <= _T_10366_13;
                                  end else begin
                                    if (_T_13005) begin
                                      _T_18065_30 <= _T_10366_14;
                                    end else begin
                                      if (_T_13003) begin
                                        _T_18065_30 <= _T_10366_15;
                                      end else begin
                                        if (_T_13001) begin
                                          _T_18065_30 <= _T_10366_16;
                                        end else begin
                                          if (_T_12999) begin
                                            _T_18065_30 <= _T_10366_17;
                                          end else begin
                                            if (_T_12997) begin
                                              _T_18065_30 <= _T_10366_18;
                                            end else begin
                                              if (_T_12995) begin
                                                _T_18065_30 <= _T_10366_19;
                                              end else begin
                                                if (_T_12993) begin
                                                  _T_18065_30 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12991) begin
                                                    _T_18065_30 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12989) begin
                                                      _T_18065_30 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_12987) begin
                                                        _T_18065_30 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_12985) begin
                                                          _T_18065_30 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_12983) begin
                                                            _T_18065_30 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_12981) begin
                                                              _T_18065_30 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_12979) begin
                                                                _T_18065_30 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_12977) begin
                                                                  _T_18065_30 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_12975) begin
                                                                    _T_18065_30 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_12973) begin
                                                                      _T_18065_30 <= _T_10366_30;
                                                                    end else begin
                                                                      _T_18065_30 <= 8'h0;
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_30 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_31) begin
        if (_T_13130) begin
          _T_18065_31 <= _T_10366_0;
        end else begin
          if (_T_13128) begin
            _T_18065_31 <= _T_10366_1;
          end else begin
            if (_T_13126) begin
              _T_18065_31 <= _T_10366_2;
            end else begin
              if (_T_13124) begin
                _T_18065_31 <= _T_10366_3;
              end else begin
                if (_T_13122) begin
                  _T_18065_31 <= _T_10366_4;
                end else begin
                  if (_T_13120) begin
                    _T_18065_31 <= _T_10366_5;
                  end else begin
                    if (_T_13118) begin
                      _T_18065_31 <= _T_10366_6;
                    end else begin
                      if (_T_13116) begin
                        _T_18065_31 <= _T_10366_7;
                      end else begin
                        if (_T_13114) begin
                          _T_18065_31 <= _T_10366_8;
                        end else begin
                          if (_T_13112) begin
                            _T_18065_31 <= _T_10366_9;
                          end else begin
                            if (_T_13110) begin
                              _T_18065_31 <= _T_10366_10;
                            end else begin
                              if (_T_13108) begin
                                _T_18065_31 <= _T_10366_11;
                              end else begin
                                if (_T_13106) begin
                                  _T_18065_31 <= _T_10366_12;
                                end else begin
                                  if (_T_13104) begin
                                    _T_18065_31 <= _T_10366_13;
                                  end else begin
                                    if (_T_13102) begin
                                      _T_18065_31 <= _T_10366_14;
                                    end else begin
                                      if (_T_13100) begin
                                        _T_18065_31 <= _T_10366_15;
                                      end else begin
                                        if (_T_13098) begin
                                          _T_18065_31 <= _T_10366_16;
                                        end else begin
                                          if (_T_13096) begin
                                            _T_18065_31 <= _T_10366_17;
                                          end else begin
                                            if (_T_13094) begin
                                              _T_18065_31 <= _T_10366_18;
                                            end else begin
                                              if (_T_13092) begin
                                                _T_18065_31 <= _T_10366_19;
                                              end else begin
                                                if (_T_13090) begin
                                                  _T_18065_31 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13088) begin
                                                    _T_18065_31 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13086) begin
                                                      _T_18065_31 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13084) begin
                                                        _T_18065_31 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13082) begin
                                                          _T_18065_31 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13080) begin
                                                            _T_18065_31 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13078) begin
                                                              _T_18065_31 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13076) begin
                                                                _T_18065_31 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13074) begin
                                                                  _T_18065_31 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13072) begin
                                                                    _T_18065_31 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13070) begin
                                                                      _T_18065_31 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13068) begin
                                                                        _T_18065_31 <= _T_10366_31;
                                                                      end else begin
                                                                        _T_18065_31 <= 8'h0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_31 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_32) begin
        if (_T_13230) begin
          _T_18065_32 <= _T_10366_0;
        end else begin
          if (_T_13228) begin
            _T_18065_32 <= _T_10366_1;
          end else begin
            if (_T_13226) begin
              _T_18065_32 <= _T_10366_2;
            end else begin
              if (_T_13224) begin
                _T_18065_32 <= _T_10366_3;
              end else begin
                if (_T_13222) begin
                  _T_18065_32 <= _T_10366_4;
                end else begin
                  if (_T_13220) begin
                    _T_18065_32 <= _T_10366_5;
                  end else begin
                    if (_T_13218) begin
                      _T_18065_32 <= _T_10366_6;
                    end else begin
                      if (_T_13216) begin
                        _T_18065_32 <= _T_10366_7;
                      end else begin
                        if (_T_13214) begin
                          _T_18065_32 <= _T_10366_8;
                        end else begin
                          if (_T_13212) begin
                            _T_18065_32 <= _T_10366_9;
                          end else begin
                            if (_T_13210) begin
                              _T_18065_32 <= _T_10366_10;
                            end else begin
                              if (_T_13208) begin
                                _T_18065_32 <= _T_10366_11;
                              end else begin
                                if (_T_13206) begin
                                  _T_18065_32 <= _T_10366_12;
                                end else begin
                                  if (_T_13204) begin
                                    _T_18065_32 <= _T_10366_13;
                                  end else begin
                                    if (_T_13202) begin
                                      _T_18065_32 <= _T_10366_14;
                                    end else begin
                                      if (_T_13200) begin
                                        _T_18065_32 <= _T_10366_15;
                                      end else begin
                                        if (_T_13198) begin
                                          _T_18065_32 <= _T_10366_16;
                                        end else begin
                                          if (_T_13196) begin
                                            _T_18065_32 <= _T_10366_17;
                                          end else begin
                                            if (_T_13194) begin
                                              _T_18065_32 <= _T_10366_18;
                                            end else begin
                                              if (_T_13192) begin
                                                _T_18065_32 <= _T_10366_19;
                                              end else begin
                                                if (_T_13190) begin
                                                  _T_18065_32 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13188) begin
                                                    _T_18065_32 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13186) begin
                                                      _T_18065_32 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13184) begin
                                                        _T_18065_32 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13182) begin
                                                          _T_18065_32 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13180) begin
                                                            _T_18065_32 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13178) begin
                                                              _T_18065_32 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13176) begin
                                                                _T_18065_32 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13174) begin
                                                                  _T_18065_32 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13172) begin
                                                                    _T_18065_32 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13170) begin
                                                                      _T_18065_32 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13168) begin
                                                                        _T_18065_32 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_13166) begin
                                                                          _T_18065_32 <= _T_10366_32;
                                                                        end else begin
                                                                          _T_18065_32 <= 8'h0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_32 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_33) begin
        if (_T_13333) begin
          _T_18065_33 <= _T_10366_0;
        end else begin
          if (_T_13331) begin
            _T_18065_33 <= _T_10366_1;
          end else begin
            if (_T_13329) begin
              _T_18065_33 <= _T_10366_2;
            end else begin
              if (_T_13327) begin
                _T_18065_33 <= _T_10366_3;
              end else begin
                if (_T_13325) begin
                  _T_18065_33 <= _T_10366_4;
                end else begin
                  if (_T_13323) begin
                    _T_18065_33 <= _T_10366_5;
                  end else begin
                    if (_T_13321) begin
                      _T_18065_33 <= _T_10366_6;
                    end else begin
                      if (_T_13319) begin
                        _T_18065_33 <= _T_10366_7;
                      end else begin
                        if (_T_13317) begin
                          _T_18065_33 <= _T_10366_8;
                        end else begin
                          if (_T_13315) begin
                            _T_18065_33 <= _T_10366_9;
                          end else begin
                            if (_T_13313) begin
                              _T_18065_33 <= _T_10366_10;
                            end else begin
                              if (_T_13311) begin
                                _T_18065_33 <= _T_10366_11;
                              end else begin
                                if (_T_13309) begin
                                  _T_18065_33 <= _T_10366_12;
                                end else begin
                                  if (_T_13307) begin
                                    _T_18065_33 <= _T_10366_13;
                                  end else begin
                                    if (_T_13305) begin
                                      _T_18065_33 <= _T_10366_14;
                                    end else begin
                                      if (_T_13303) begin
                                        _T_18065_33 <= _T_10366_15;
                                      end else begin
                                        if (_T_13301) begin
                                          _T_18065_33 <= _T_10366_16;
                                        end else begin
                                          if (_T_13299) begin
                                            _T_18065_33 <= _T_10366_17;
                                          end else begin
                                            if (_T_13297) begin
                                              _T_18065_33 <= _T_10366_18;
                                            end else begin
                                              if (_T_13295) begin
                                                _T_18065_33 <= _T_10366_19;
                                              end else begin
                                                if (_T_13293) begin
                                                  _T_18065_33 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13291) begin
                                                    _T_18065_33 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13289) begin
                                                      _T_18065_33 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13287) begin
                                                        _T_18065_33 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13285) begin
                                                          _T_18065_33 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13283) begin
                                                            _T_18065_33 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13281) begin
                                                              _T_18065_33 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13279) begin
                                                                _T_18065_33 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13277) begin
                                                                  _T_18065_33 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13275) begin
                                                                    _T_18065_33 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13273) begin
                                                                      _T_18065_33 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13271) begin
                                                                        _T_18065_33 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_13269) begin
                                                                          _T_18065_33 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_13267) begin
                                                                            _T_18065_33 <= _T_10366_33;
                                                                          end else begin
                                                                            _T_18065_33 <= 8'h0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_33 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_34) begin
        if (_T_13439) begin
          _T_18065_34 <= _T_10366_0;
        end else begin
          if (_T_13437) begin
            _T_18065_34 <= _T_10366_1;
          end else begin
            if (_T_13435) begin
              _T_18065_34 <= _T_10366_2;
            end else begin
              if (_T_13433) begin
                _T_18065_34 <= _T_10366_3;
              end else begin
                if (_T_13431) begin
                  _T_18065_34 <= _T_10366_4;
                end else begin
                  if (_T_13429) begin
                    _T_18065_34 <= _T_10366_5;
                  end else begin
                    if (_T_13427) begin
                      _T_18065_34 <= _T_10366_6;
                    end else begin
                      if (_T_13425) begin
                        _T_18065_34 <= _T_10366_7;
                      end else begin
                        if (_T_13423) begin
                          _T_18065_34 <= _T_10366_8;
                        end else begin
                          if (_T_13421) begin
                            _T_18065_34 <= _T_10366_9;
                          end else begin
                            if (_T_13419) begin
                              _T_18065_34 <= _T_10366_10;
                            end else begin
                              if (_T_13417) begin
                                _T_18065_34 <= _T_10366_11;
                              end else begin
                                if (_T_13415) begin
                                  _T_18065_34 <= _T_10366_12;
                                end else begin
                                  if (_T_13413) begin
                                    _T_18065_34 <= _T_10366_13;
                                  end else begin
                                    if (_T_13411) begin
                                      _T_18065_34 <= _T_10366_14;
                                    end else begin
                                      if (_T_13409) begin
                                        _T_18065_34 <= _T_10366_15;
                                      end else begin
                                        if (_T_13407) begin
                                          _T_18065_34 <= _T_10366_16;
                                        end else begin
                                          if (_T_13405) begin
                                            _T_18065_34 <= _T_10366_17;
                                          end else begin
                                            if (_T_13403) begin
                                              _T_18065_34 <= _T_10366_18;
                                            end else begin
                                              if (_T_13401) begin
                                                _T_18065_34 <= _T_10366_19;
                                              end else begin
                                                if (_T_13399) begin
                                                  _T_18065_34 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13397) begin
                                                    _T_18065_34 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13395) begin
                                                      _T_18065_34 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13393) begin
                                                        _T_18065_34 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13391) begin
                                                          _T_18065_34 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13389) begin
                                                            _T_18065_34 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13387) begin
                                                              _T_18065_34 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13385) begin
                                                                _T_18065_34 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13383) begin
                                                                  _T_18065_34 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13381) begin
                                                                    _T_18065_34 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13379) begin
                                                                      _T_18065_34 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13377) begin
                                                                        _T_18065_34 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_13375) begin
                                                                          _T_18065_34 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_13373) begin
                                                                            _T_18065_34 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_13371) begin
                                                                              _T_18065_34 <= _T_10366_34;
                                                                            end else begin
                                                                              _T_18065_34 <= 8'h0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_34 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_35) begin
        if (_T_13548) begin
          _T_18065_35 <= _T_10366_0;
        end else begin
          if (_T_13546) begin
            _T_18065_35 <= _T_10366_1;
          end else begin
            if (_T_13544) begin
              _T_18065_35 <= _T_10366_2;
            end else begin
              if (_T_13542) begin
                _T_18065_35 <= _T_10366_3;
              end else begin
                if (_T_13540) begin
                  _T_18065_35 <= _T_10366_4;
                end else begin
                  if (_T_13538) begin
                    _T_18065_35 <= _T_10366_5;
                  end else begin
                    if (_T_13536) begin
                      _T_18065_35 <= _T_10366_6;
                    end else begin
                      if (_T_13534) begin
                        _T_18065_35 <= _T_10366_7;
                      end else begin
                        if (_T_13532) begin
                          _T_18065_35 <= _T_10366_8;
                        end else begin
                          if (_T_13530) begin
                            _T_18065_35 <= _T_10366_9;
                          end else begin
                            if (_T_13528) begin
                              _T_18065_35 <= _T_10366_10;
                            end else begin
                              if (_T_13526) begin
                                _T_18065_35 <= _T_10366_11;
                              end else begin
                                if (_T_13524) begin
                                  _T_18065_35 <= _T_10366_12;
                                end else begin
                                  if (_T_13522) begin
                                    _T_18065_35 <= _T_10366_13;
                                  end else begin
                                    if (_T_13520) begin
                                      _T_18065_35 <= _T_10366_14;
                                    end else begin
                                      if (_T_13518) begin
                                        _T_18065_35 <= _T_10366_15;
                                      end else begin
                                        if (_T_13516) begin
                                          _T_18065_35 <= _T_10366_16;
                                        end else begin
                                          if (_T_13514) begin
                                            _T_18065_35 <= _T_10366_17;
                                          end else begin
                                            if (_T_13512) begin
                                              _T_18065_35 <= _T_10366_18;
                                            end else begin
                                              if (_T_13510) begin
                                                _T_18065_35 <= _T_10366_19;
                                              end else begin
                                                if (_T_13508) begin
                                                  _T_18065_35 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13506) begin
                                                    _T_18065_35 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13504) begin
                                                      _T_18065_35 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13502) begin
                                                        _T_18065_35 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13500) begin
                                                          _T_18065_35 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13498) begin
                                                            _T_18065_35 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13496) begin
                                                              _T_18065_35 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13494) begin
                                                                _T_18065_35 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13492) begin
                                                                  _T_18065_35 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13490) begin
                                                                    _T_18065_35 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13488) begin
                                                                      _T_18065_35 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13486) begin
                                                                        _T_18065_35 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_13484) begin
                                                                          _T_18065_35 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_13482) begin
                                                                            _T_18065_35 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_13480) begin
                                                                              _T_18065_35 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_13478) begin
                                                                                _T_18065_35 <= _T_10366_35;
                                                                              end else begin
                                                                                _T_18065_35 <= 8'h0;
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_35 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_36) begin
        if (_T_13660) begin
          _T_18065_36 <= _T_10366_0;
        end else begin
          if (_T_13658) begin
            _T_18065_36 <= _T_10366_1;
          end else begin
            if (_T_13656) begin
              _T_18065_36 <= _T_10366_2;
            end else begin
              if (_T_13654) begin
                _T_18065_36 <= _T_10366_3;
              end else begin
                if (_T_13652) begin
                  _T_18065_36 <= _T_10366_4;
                end else begin
                  if (_T_13650) begin
                    _T_18065_36 <= _T_10366_5;
                  end else begin
                    if (_T_13648) begin
                      _T_18065_36 <= _T_10366_6;
                    end else begin
                      if (_T_13646) begin
                        _T_18065_36 <= _T_10366_7;
                      end else begin
                        if (_T_13644) begin
                          _T_18065_36 <= _T_10366_8;
                        end else begin
                          if (_T_13642) begin
                            _T_18065_36 <= _T_10366_9;
                          end else begin
                            if (_T_13640) begin
                              _T_18065_36 <= _T_10366_10;
                            end else begin
                              if (_T_13638) begin
                                _T_18065_36 <= _T_10366_11;
                              end else begin
                                if (_T_13636) begin
                                  _T_18065_36 <= _T_10366_12;
                                end else begin
                                  if (_T_13634) begin
                                    _T_18065_36 <= _T_10366_13;
                                  end else begin
                                    if (_T_13632) begin
                                      _T_18065_36 <= _T_10366_14;
                                    end else begin
                                      if (_T_13630) begin
                                        _T_18065_36 <= _T_10366_15;
                                      end else begin
                                        if (_T_13628) begin
                                          _T_18065_36 <= _T_10366_16;
                                        end else begin
                                          if (_T_13626) begin
                                            _T_18065_36 <= _T_10366_17;
                                          end else begin
                                            if (_T_13624) begin
                                              _T_18065_36 <= _T_10366_18;
                                            end else begin
                                              if (_T_13622) begin
                                                _T_18065_36 <= _T_10366_19;
                                              end else begin
                                                if (_T_13620) begin
                                                  _T_18065_36 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13618) begin
                                                    _T_18065_36 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13616) begin
                                                      _T_18065_36 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13614) begin
                                                        _T_18065_36 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13612) begin
                                                          _T_18065_36 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13610) begin
                                                            _T_18065_36 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13608) begin
                                                              _T_18065_36 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13606) begin
                                                                _T_18065_36 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13604) begin
                                                                  _T_18065_36 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13602) begin
                                                                    _T_18065_36 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13600) begin
                                                                      _T_18065_36 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13598) begin
                                                                        _T_18065_36 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_13596) begin
                                                                          _T_18065_36 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_13594) begin
                                                                            _T_18065_36 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_13592) begin
                                                                              _T_18065_36 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_13590) begin
                                                                                _T_18065_36 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_13588) begin
                                                                                  _T_18065_36 <= _T_10366_36;
                                                                                end else begin
                                                                                  _T_18065_36 <= 8'h0;
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_36 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_37) begin
        if (_T_13775) begin
          _T_18065_37 <= _T_10366_0;
        end else begin
          if (_T_13773) begin
            _T_18065_37 <= _T_10366_1;
          end else begin
            if (_T_13771) begin
              _T_18065_37 <= _T_10366_2;
            end else begin
              if (_T_13769) begin
                _T_18065_37 <= _T_10366_3;
              end else begin
                if (_T_13767) begin
                  _T_18065_37 <= _T_10366_4;
                end else begin
                  if (_T_13765) begin
                    _T_18065_37 <= _T_10366_5;
                  end else begin
                    if (_T_13763) begin
                      _T_18065_37 <= _T_10366_6;
                    end else begin
                      if (_T_13761) begin
                        _T_18065_37 <= _T_10366_7;
                      end else begin
                        if (_T_13759) begin
                          _T_18065_37 <= _T_10366_8;
                        end else begin
                          if (_T_13757) begin
                            _T_18065_37 <= _T_10366_9;
                          end else begin
                            if (_T_13755) begin
                              _T_18065_37 <= _T_10366_10;
                            end else begin
                              if (_T_13753) begin
                                _T_18065_37 <= _T_10366_11;
                              end else begin
                                if (_T_13751) begin
                                  _T_18065_37 <= _T_10366_12;
                                end else begin
                                  if (_T_13749) begin
                                    _T_18065_37 <= _T_10366_13;
                                  end else begin
                                    if (_T_13747) begin
                                      _T_18065_37 <= _T_10366_14;
                                    end else begin
                                      if (_T_13745) begin
                                        _T_18065_37 <= _T_10366_15;
                                      end else begin
                                        if (_T_13743) begin
                                          _T_18065_37 <= _T_10366_16;
                                        end else begin
                                          if (_T_13741) begin
                                            _T_18065_37 <= _T_10366_17;
                                          end else begin
                                            if (_T_13739) begin
                                              _T_18065_37 <= _T_10366_18;
                                            end else begin
                                              if (_T_13737) begin
                                                _T_18065_37 <= _T_10366_19;
                                              end else begin
                                                if (_T_13735) begin
                                                  _T_18065_37 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13733) begin
                                                    _T_18065_37 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13731) begin
                                                      _T_18065_37 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13729) begin
                                                        _T_18065_37 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13727) begin
                                                          _T_18065_37 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13725) begin
                                                            _T_18065_37 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13723) begin
                                                              _T_18065_37 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13721) begin
                                                                _T_18065_37 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13719) begin
                                                                  _T_18065_37 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13717) begin
                                                                    _T_18065_37 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13715) begin
                                                                      _T_18065_37 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13713) begin
                                                                        _T_18065_37 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_13711) begin
                                                                          _T_18065_37 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_13709) begin
                                                                            _T_18065_37 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_13707) begin
                                                                              _T_18065_37 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_13705) begin
                                                                                _T_18065_37 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_13703) begin
                                                                                  _T_18065_37 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_13701) begin
                                                                                    _T_18065_37 <= _T_10366_37;
                                                                                  end else begin
                                                                                    _T_18065_37 <= 8'h0;
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_37 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_38) begin
        if (_T_13893) begin
          _T_18065_38 <= _T_10366_0;
        end else begin
          if (_T_13891) begin
            _T_18065_38 <= _T_10366_1;
          end else begin
            if (_T_13889) begin
              _T_18065_38 <= _T_10366_2;
            end else begin
              if (_T_13887) begin
                _T_18065_38 <= _T_10366_3;
              end else begin
                if (_T_13885) begin
                  _T_18065_38 <= _T_10366_4;
                end else begin
                  if (_T_13883) begin
                    _T_18065_38 <= _T_10366_5;
                  end else begin
                    if (_T_13881) begin
                      _T_18065_38 <= _T_10366_6;
                    end else begin
                      if (_T_13879) begin
                        _T_18065_38 <= _T_10366_7;
                      end else begin
                        if (_T_13877) begin
                          _T_18065_38 <= _T_10366_8;
                        end else begin
                          if (_T_13875) begin
                            _T_18065_38 <= _T_10366_9;
                          end else begin
                            if (_T_13873) begin
                              _T_18065_38 <= _T_10366_10;
                            end else begin
                              if (_T_13871) begin
                                _T_18065_38 <= _T_10366_11;
                              end else begin
                                if (_T_13869) begin
                                  _T_18065_38 <= _T_10366_12;
                                end else begin
                                  if (_T_13867) begin
                                    _T_18065_38 <= _T_10366_13;
                                  end else begin
                                    if (_T_13865) begin
                                      _T_18065_38 <= _T_10366_14;
                                    end else begin
                                      if (_T_13863) begin
                                        _T_18065_38 <= _T_10366_15;
                                      end else begin
                                        if (_T_13861) begin
                                          _T_18065_38 <= _T_10366_16;
                                        end else begin
                                          if (_T_13859) begin
                                            _T_18065_38 <= _T_10366_17;
                                          end else begin
                                            if (_T_13857) begin
                                              _T_18065_38 <= _T_10366_18;
                                            end else begin
                                              if (_T_13855) begin
                                                _T_18065_38 <= _T_10366_19;
                                              end else begin
                                                if (_T_13853) begin
                                                  _T_18065_38 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13851) begin
                                                    _T_18065_38 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13849) begin
                                                      _T_18065_38 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13847) begin
                                                        _T_18065_38 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13845) begin
                                                          _T_18065_38 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13843) begin
                                                            _T_18065_38 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13841) begin
                                                              _T_18065_38 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13839) begin
                                                                _T_18065_38 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13837) begin
                                                                  _T_18065_38 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13835) begin
                                                                    _T_18065_38 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13833) begin
                                                                      _T_18065_38 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13831) begin
                                                                        _T_18065_38 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_13829) begin
                                                                          _T_18065_38 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_13827) begin
                                                                            _T_18065_38 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_13825) begin
                                                                              _T_18065_38 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_13823) begin
                                                                                _T_18065_38 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_13821) begin
                                                                                  _T_18065_38 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_13819) begin
                                                                                    _T_18065_38 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_13817) begin
                                                                                      _T_18065_38 <= _T_10366_38;
                                                                                    end else begin
                                                                                      _T_18065_38 <= 8'h0;
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_38 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_39) begin
        if (_T_14014) begin
          _T_18065_39 <= _T_10366_0;
        end else begin
          if (_T_14012) begin
            _T_18065_39 <= _T_10366_1;
          end else begin
            if (_T_14010) begin
              _T_18065_39 <= _T_10366_2;
            end else begin
              if (_T_14008) begin
                _T_18065_39 <= _T_10366_3;
              end else begin
                if (_T_14006) begin
                  _T_18065_39 <= _T_10366_4;
                end else begin
                  if (_T_14004) begin
                    _T_18065_39 <= _T_10366_5;
                  end else begin
                    if (_T_14002) begin
                      _T_18065_39 <= _T_10366_6;
                    end else begin
                      if (_T_14000) begin
                        _T_18065_39 <= _T_10366_7;
                      end else begin
                        if (_T_13998) begin
                          _T_18065_39 <= _T_10366_8;
                        end else begin
                          if (_T_13996) begin
                            _T_18065_39 <= _T_10366_9;
                          end else begin
                            if (_T_13994) begin
                              _T_18065_39 <= _T_10366_10;
                            end else begin
                              if (_T_13992) begin
                                _T_18065_39 <= _T_10366_11;
                              end else begin
                                if (_T_13990) begin
                                  _T_18065_39 <= _T_10366_12;
                                end else begin
                                  if (_T_13988) begin
                                    _T_18065_39 <= _T_10366_13;
                                  end else begin
                                    if (_T_13986) begin
                                      _T_18065_39 <= _T_10366_14;
                                    end else begin
                                      if (_T_13984) begin
                                        _T_18065_39 <= _T_10366_15;
                                      end else begin
                                        if (_T_13982) begin
                                          _T_18065_39 <= _T_10366_16;
                                        end else begin
                                          if (_T_13980) begin
                                            _T_18065_39 <= _T_10366_17;
                                          end else begin
                                            if (_T_13978) begin
                                              _T_18065_39 <= _T_10366_18;
                                            end else begin
                                              if (_T_13976) begin
                                                _T_18065_39 <= _T_10366_19;
                                              end else begin
                                                if (_T_13974) begin
                                                  _T_18065_39 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13972) begin
                                                    _T_18065_39 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13970) begin
                                                      _T_18065_39 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13968) begin
                                                        _T_18065_39 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13966) begin
                                                          _T_18065_39 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13964) begin
                                                            _T_18065_39 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13962) begin
                                                              _T_18065_39 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13960) begin
                                                                _T_18065_39 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13958) begin
                                                                  _T_18065_39 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13956) begin
                                                                    _T_18065_39 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13954) begin
                                                                      _T_18065_39 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13952) begin
                                                                        _T_18065_39 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_13950) begin
                                                                          _T_18065_39 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_13948) begin
                                                                            _T_18065_39 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_13946) begin
                                                                              _T_18065_39 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_13944) begin
                                                                                _T_18065_39 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_13942) begin
                                                                                  _T_18065_39 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_13940) begin
                                                                                    _T_18065_39 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_13938) begin
                                                                                      _T_18065_39 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_13936) begin
                                                                                        _T_18065_39 <= _T_10366_39;
                                                                                      end else begin
                                                                                        _T_18065_39 <= 8'h0;
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_39 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_40) begin
        if (_T_14138) begin
          _T_18065_40 <= _T_10366_0;
        end else begin
          if (_T_14136) begin
            _T_18065_40 <= _T_10366_1;
          end else begin
            if (_T_14134) begin
              _T_18065_40 <= _T_10366_2;
            end else begin
              if (_T_14132) begin
                _T_18065_40 <= _T_10366_3;
              end else begin
                if (_T_14130) begin
                  _T_18065_40 <= _T_10366_4;
                end else begin
                  if (_T_14128) begin
                    _T_18065_40 <= _T_10366_5;
                  end else begin
                    if (_T_14126) begin
                      _T_18065_40 <= _T_10366_6;
                    end else begin
                      if (_T_14124) begin
                        _T_18065_40 <= _T_10366_7;
                      end else begin
                        if (_T_14122) begin
                          _T_18065_40 <= _T_10366_8;
                        end else begin
                          if (_T_14120) begin
                            _T_18065_40 <= _T_10366_9;
                          end else begin
                            if (_T_14118) begin
                              _T_18065_40 <= _T_10366_10;
                            end else begin
                              if (_T_14116) begin
                                _T_18065_40 <= _T_10366_11;
                              end else begin
                                if (_T_14114) begin
                                  _T_18065_40 <= _T_10366_12;
                                end else begin
                                  if (_T_14112) begin
                                    _T_18065_40 <= _T_10366_13;
                                  end else begin
                                    if (_T_14110) begin
                                      _T_18065_40 <= _T_10366_14;
                                    end else begin
                                      if (_T_14108) begin
                                        _T_18065_40 <= _T_10366_15;
                                      end else begin
                                        if (_T_14106) begin
                                          _T_18065_40 <= _T_10366_16;
                                        end else begin
                                          if (_T_14104) begin
                                            _T_18065_40 <= _T_10366_17;
                                          end else begin
                                            if (_T_14102) begin
                                              _T_18065_40 <= _T_10366_18;
                                            end else begin
                                              if (_T_14100) begin
                                                _T_18065_40 <= _T_10366_19;
                                              end else begin
                                                if (_T_14098) begin
                                                  _T_18065_40 <= _T_10366_20;
                                                end else begin
                                                  if (_T_14096) begin
                                                    _T_18065_40 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_14094) begin
                                                      _T_18065_40 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_14092) begin
                                                        _T_18065_40 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_14090) begin
                                                          _T_18065_40 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_14088) begin
                                                            _T_18065_40 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_14086) begin
                                                              _T_18065_40 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_14084) begin
                                                                _T_18065_40 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_14082) begin
                                                                  _T_18065_40 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_14080) begin
                                                                    _T_18065_40 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_14078) begin
                                                                      _T_18065_40 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_14076) begin
                                                                        _T_18065_40 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_14074) begin
                                                                          _T_18065_40 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_14072) begin
                                                                            _T_18065_40 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_14070) begin
                                                                              _T_18065_40 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_14068) begin
                                                                                _T_18065_40 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_14066) begin
                                                                                  _T_18065_40 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_14064) begin
                                                                                    _T_18065_40 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_14062) begin
                                                                                      _T_18065_40 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_14060) begin
                                                                                        _T_18065_40 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_14058) begin
                                                                                          _T_18065_40 <= _T_10366_40;
                                                                                        end else begin
                                                                                          _T_18065_40 <= 8'h0;
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_40 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_41) begin
        if (_T_14265) begin
          _T_18065_41 <= _T_10366_0;
        end else begin
          if (_T_14263) begin
            _T_18065_41 <= _T_10366_1;
          end else begin
            if (_T_14261) begin
              _T_18065_41 <= _T_10366_2;
            end else begin
              if (_T_14259) begin
                _T_18065_41 <= _T_10366_3;
              end else begin
                if (_T_14257) begin
                  _T_18065_41 <= _T_10366_4;
                end else begin
                  if (_T_14255) begin
                    _T_18065_41 <= _T_10366_5;
                  end else begin
                    if (_T_14253) begin
                      _T_18065_41 <= _T_10366_6;
                    end else begin
                      if (_T_14251) begin
                        _T_18065_41 <= _T_10366_7;
                      end else begin
                        if (_T_14249) begin
                          _T_18065_41 <= _T_10366_8;
                        end else begin
                          if (_T_14247) begin
                            _T_18065_41 <= _T_10366_9;
                          end else begin
                            if (_T_14245) begin
                              _T_18065_41 <= _T_10366_10;
                            end else begin
                              if (_T_14243) begin
                                _T_18065_41 <= _T_10366_11;
                              end else begin
                                if (_T_14241) begin
                                  _T_18065_41 <= _T_10366_12;
                                end else begin
                                  if (_T_14239) begin
                                    _T_18065_41 <= _T_10366_13;
                                  end else begin
                                    if (_T_14237) begin
                                      _T_18065_41 <= _T_10366_14;
                                    end else begin
                                      if (_T_14235) begin
                                        _T_18065_41 <= _T_10366_15;
                                      end else begin
                                        if (_T_14233) begin
                                          _T_18065_41 <= _T_10366_16;
                                        end else begin
                                          if (_T_14231) begin
                                            _T_18065_41 <= _T_10366_17;
                                          end else begin
                                            if (_T_14229) begin
                                              _T_18065_41 <= _T_10366_18;
                                            end else begin
                                              if (_T_14227) begin
                                                _T_18065_41 <= _T_10366_19;
                                              end else begin
                                                if (_T_14225) begin
                                                  _T_18065_41 <= _T_10366_20;
                                                end else begin
                                                  if (_T_14223) begin
                                                    _T_18065_41 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_14221) begin
                                                      _T_18065_41 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_14219) begin
                                                        _T_18065_41 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_14217) begin
                                                          _T_18065_41 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_14215) begin
                                                            _T_18065_41 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_14213) begin
                                                              _T_18065_41 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_14211) begin
                                                                _T_18065_41 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_14209) begin
                                                                  _T_18065_41 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_14207) begin
                                                                    _T_18065_41 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_14205) begin
                                                                      _T_18065_41 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_14203) begin
                                                                        _T_18065_41 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_14201) begin
                                                                          _T_18065_41 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_14199) begin
                                                                            _T_18065_41 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_14197) begin
                                                                              _T_18065_41 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_14195) begin
                                                                                _T_18065_41 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_14193) begin
                                                                                  _T_18065_41 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_14191) begin
                                                                                    _T_18065_41 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_14189) begin
                                                                                      _T_18065_41 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_14187) begin
                                                                                        _T_18065_41 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_14185) begin
                                                                                          _T_18065_41 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_14183) begin
                                                                                            _T_18065_41 <= _T_10366_41;
                                                                                          end else begin
                                                                                            _T_18065_41 <= 8'h0;
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_41 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_42) begin
        if (_T_14395) begin
          _T_18065_42 <= _T_10366_0;
        end else begin
          if (_T_14393) begin
            _T_18065_42 <= _T_10366_1;
          end else begin
            if (_T_14391) begin
              _T_18065_42 <= _T_10366_2;
            end else begin
              if (_T_14389) begin
                _T_18065_42 <= _T_10366_3;
              end else begin
                if (_T_14387) begin
                  _T_18065_42 <= _T_10366_4;
                end else begin
                  if (_T_14385) begin
                    _T_18065_42 <= _T_10366_5;
                  end else begin
                    if (_T_14383) begin
                      _T_18065_42 <= _T_10366_6;
                    end else begin
                      if (_T_14381) begin
                        _T_18065_42 <= _T_10366_7;
                      end else begin
                        if (_T_14379) begin
                          _T_18065_42 <= _T_10366_8;
                        end else begin
                          if (_T_14377) begin
                            _T_18065_42 <= _T_10366_9;
                          end else begin
                            if (_T_14375) begin
                              _T_18065_42 <= _T_10366_10;
                            end else begin
                              if (_T_14373) begin
                                _T_18065_42 <= _T_10366_11;
                              end else begin
                                if (_T_14371) begin
                                  _T_18065_42 <= _T_10366_12;
                                end else begin
                                  if (_T_14369) begin
                                    _T_18065_42 <= _T_10366_13;
                                  end else begin
                                    if (_T_14367) begin
                                      _T_18065_42 <= _T_10366_14;
                                    end else begin
                                      if (_T_14365) begin
                                        _T_18065_42 <= _T_10366_15;
                                      end else begin
                                        if (_T_14363) begin
                                          _T_18065_42 <= _T_10366_16;
                                        end else begin
                                          if (_T_14361) begin
                                            _T_18065_42 <= _T_10366_17;
                                          end else begin
                                            if (_T_14359) begin
                                              _T_18065_42 <= _T_10366_18;
                                            end else begin
                                              if (_T_14357) begin
                                                _T_18065_42 <= _T_10366_19;
                                              end else begin
                                                if (_T_14355) begin
                                                  _T_18065_42 <= _T_10366_20;
                                                end else begin
                                                  if (_T_14353) begin
                                                    _T_18065_42 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_14351) begin
                                                      _T_18065_42 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_14349) begin
                                                        _T_18065_42 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_14347) begin
                                                          _T_18065_42 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_14345) begin
                                                            _T_18065_42 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_14343) begin
                                                              _T_18065_42 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_14341) begin
                                                                _T_18065_42 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_14339) begin
                                                                  _T_18065_42 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_14337) begin
                                                                    _T_18065_42 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_14335) begin
                                                                      _T_18065_42 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_14333) begin
                                                                        _T_18065_42 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_14331) begin
                                                                          _T_18065_42 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_14329) begin
                                                                            _T_18065_42 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_14327) begin
                                                                              _T_18065_42 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_14325) begin
                                                                                _T_18065_42 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_14323) begin
                                                                                  _T_18065_42 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_14321) begin
                                                                                    _T_18065_42 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_14319) begin
                                                                                      _T_18065_42 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_14317) begin
                                                                                        _T_18065_42 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_14315) begin
                                                                                          _T_18065_42 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_14313) begin
                                                                                            _T_18065_42 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_14311) begin
                                                                                              _T_18065_42 <= _T_10366_42;
                                                                                            end else begin
                                                                                              _T_18065_42 <= 8'h0;
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_42 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_43) begin
        if (_T_14528) begin
          _T_18065_43 <= _T_10366_0;
        end else begin
          if (_T_14526) begin
            _T_18065_43 <= _T_10366_1;
          end else begin
            if (_T_14524) begin
              _T_18065_43 <= _T_10366_2;
            end else begin
              if (_T_14522) begin
                _T_18065_43 <= _T_10366_3;
              end else begin
                if (_T_14520) begin
                  _T_18065_43 <= _T_10366_4;
                end else begin
                  if (_T_14518) begin
                    _T_18065_43 <= _T_10366_5;
                  end else begin
                    if (_T_14516) begin
                      _T_18065_43 <= _T_10366_6;
                    end else begin
                      if (_T_14514) begin
                        _T_18065_43 <= _T_10366_7;
                      end else begin
                        if (_T_14512) begin
                          _T_18065_43 <= _T_10366_8;
                        end else begin
                          if (_T_14510) begin
                            _T_18065_43 <= _T_10366_9;
                          end else begin
                            if (_T_14508) begin
                              _T_18065_43 <= _T_10366_10;
                            end else begin
                              if (_T_14506) begin
                                _T_18065_43 <= _T_10366_11;
                              end else begin
                                if (_T_14504) begin
                                  _T_18065_43 <= _T_10366_12;
                                end else begin
                                  if (_T_14502) begin
                                    _T_18065_43 <= _T_10366_13;
                                  end else begin
                                    if (_T_14500) begin
                                      _T_18065_43 <= _T_10366_14;
                                    end else begin
                                      if (_T_14498) begin
                                        _T_18065_43 <= _T_10366_15;
                                      end else begin
                                        if (_T_14496) begin
                                          _T_18065_43 <= _T_10366_16;
                                        end else begin
                                          if (_T_14494) begin
                                            _T_18065_43 <= _T_10366_17;
                                          end else begin
                                            if (_T_14492) begin
                                              _T_18065_43 <= _T_10366_18;
                                            end else begin
                                              if (_T_14490) begin
                                                _T_18065_43 <= _T_10366_19;
                                              end else begin
                                                if (_T_14488) begin
                                                  _T_18065_43 <= _T_10366_20;
                                                end else begin
                                                  if (_T_14486) begin
                                                    _T_18065_43 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_14484) begin
                                                      _T_18065_43 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_14482) begin
                                                        _T_18065_43 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_14480) begin
                                                          _T_18065_43 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_14478) begin
                                                            _T_18065_43 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_14476) begin
                                                              _T_18065_43 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_14474) begin
                                                                _T_18065_43 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_14472) begin
                                                                  _T_18065_43 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_14470) begin
                                                                    _T_18065_43 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_14468) begin
                                                                      _T_18065_43 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_14466) begin
                                                                        _T_18065_43 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_14464) begin
                                                                          _T_18065_43 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_14462) begin
                                                                            _T_18065_43 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_14460) begin
                                                                              _T_18065_43 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_14458) begin
                                                                                _T_18065_43 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_14456) begin
                                                                                  _T_18065_43 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_14454) begin
                                                                                    _T_18065_43 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_14452) begin
                                                                                      _T_18065_43 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_14450) begin
                                                                                        _T_18065_43 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_14448) begin
                                                                                          _T_18065_43 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_14446) begin
                                                                                            _T_18065_43 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_14444) begin
                                                                                              _T_18065_43 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_14442) begin
                                                                                                _T_18065_43 <= _T_10366_43;
                                                                                              end else begin
                                                                                                _T_18065_43 <= 8'h0;
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_43 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_44) begin
        if (_T_14664) begin
          _T_18065_44 <= _T_10366_0;
        end else begin
          if (_T_14662) begin
            _T_18065_44 <= _T_10366_1;
          end else begin
            if (_T_14660) begin
              _T_18065_44 <= _T_10366_2;
            end else begin
              if (_T_14658) begin
                _T_18065_44 <= _T_10366_3;
              end else begin
                if (_T_14656) begin
                  _T_18065_44 <= _T_10366_4;
                end else begin
                  if (_T_14654) begin
                    _T_18065_44 <= _T_10366_5;
                  end else begin
                    if (_T_14652) begin
                      _T_18065_44 <= _T_10366_6;
                    end else begin
                      if (_T_14650) begin
                        _T_18065_44 <= _T_10366_7;
                      end else begin
                        if (_T_14648) begin
                          _T_18065_44 <= _T_10366_8;
                        end else begin
                          if (_T_14646) begin
                            _T_18065_44 <= _T_10366_9;
                          end else begin
                            if (_T_14644) begin
                              _T_18065_44 <= _T_10366_10;
                            end else begin
                              if (_T_14642) begin
                                _T_18065_44 <= _T_10366_11;
                              end else begin
                                if (_T_14640) begin
                                  _T_18065_44 <= _T_10366_12;
                                end else begin
                                  if (_T_14638) begin
                                    _T_18065_44 <= _T_10366_13;
                                  end else begin
                                    if (_T_14636) begin
                                      _T_18065_44 <= _T_10366_14;
                                    end else begin
                                      if (_T_14634) begin
                                        _T_18065_44 <= _T_10366_15;
                                      end else begin
                                        if (_T_14632) begin
                                          _T_18065_44 <= _T_10366_16;
                                        end else begin
                                          if (_T_14630) begin
                                            _T_18065_44 <= _T_10366_17;
                                          end else begin
                                            if (_T_14628) begin
                                              _T_18065_44 <= _T_10366_18;
                                            end else begin
                                              if (_T_14626) begin
                                                _T_18065_44 <= _T_10366_19;
                                              end else begin
                                                if (_T_14624) begin
                                                  _T_18065_44 <= _T_10366_20;
                                                end else begin
                                                  if (_T_14622) begin
                                                    _T_18065_44 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_14620) begin
                                                      _T_18065_44 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_14618) begin
                                                        _T_18065_44 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_14616) begin
                                                          _T_18065_44 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_14614) begin
                                                            _T_18065_44 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_14612) begin
                                                              _T_18065_44 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_14610) begin
                                                                _T_18065_44 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_14608) begin
                                                                  _T_18065_44 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_14606) begin
                                                                    _T_18065_44 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_14604) begin
                                                                      _T_18065_44 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_14602) begin
                                                                        _T_18065_44 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_14600) begin
                                                                          _T_18065_44 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_14598) begin
                                                                            _T_18065_44 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_14596) begin
                                                                              _T_18065_44 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_14594) begin
                                                                                _T_18065_44 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_14592) begin
                                                                                  _T_18065_44 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_14590) begin
                                                                                    _T_18065_44 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_14588) begin
                                                                                      _T_18065_44 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_14586) begin
                                                                                        _T_18065_44 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_14584) begin
                                                                                          _T_18065_44 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_14582) begin
                                                                                            _T_18065_44 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_14580) begin
                                                                                              _T_18065_44 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_14578) begin
                                                                                                _T_18065_44 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_14576) begin
                                                                                                  _T_18065_44 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  _T_18065_44 <= 8'h0;
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_44 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_45) begin
        if (_T_14803) begin
          _T_18065_45 <= _T_10366_0;
        end else begin
          if (_T_14801) begin
            _T_18065_45 <= _T_10366_1;
          end else begin
            if (_T_14799) begin
              _T_18065_45 <= _T_10366_2;
            end else begin
              if (_T_14797) begin
                _T_18065_45 <= _T_10366_3;
              end else begin
                if (_T_14795) begin
                  _T_18065_45 <= _T_10366_4;
                end else begin
                  if (_T_14793) begin
                    _T_18065_45 <= _T_10366_5;
                  end else begin
                    if (_T_14791) begin
                      _T_18065_45 <= _T_10366_6;
                    end else begin
                      if (_T_14789) begin
                        _T_18065_45 <= _T_10366_7;
                      end else begin
                        if (_T_14787) begin
                          _T_18065_45 <= _T_10366_8;
                        end else begin
                          if (_T_14785) begin
                            _T_18065_45 <= _T_10366_9;
                          end else begin
                            if (_T_14783) begin
                              _T_18065_45 <= _T_10366_10;
                            end else begin
                              if (_T_14781) begin
                                _T_18065_45 <= _T_10366_11;
                              end else begin
                                if (_T_14779) begin
                                  _T_18065_45 <= _T_10366_12;
                                end else begin
                                  if (_T_14777) begin
                                    _T_18065_45 <= _T_10366_13;
                                  end else begin
                                    if (_T_14775) begin
                                      _T_18065_45 <= _T_10366_14;
                                    end else begin
                                      if (_T_14773) begin
                                        _T_18065_45 <= _T_10366_15;
                                      end else begin
                                        if (_T_14771) begin
                                          _T_18065_45 <= _T_10366_16;
                                        end else begin
                                          if (_T_14769) begin
                                            _T_18065_45 <= _T_10366_17;
                                          end else begin
                                            if (_T_14767) begin
                                              _T_18065_45 <= _T_10366_18;
                                            end else begin
                                              if (_T_14765) begin
                                                _T_18065_45 <= _T_10366_19;
                                              end else begin
                                                if (_T_14763) begin
                                                  _T_18065_45 <= _T_10366_20;
                                                end else begin
                                                  if (_T_14761) begin
                                                    _T_18065_45 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_14759) begin
                                                      _T_18065_45 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_14757) begin
                                                        _T_18065_45 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_14755) begin
                                                          _T_18065_45 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_14753) begin
                                                            _T_18065_45 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_14751) begin
                                                              _T_18065_45 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_14749) begin
                                                                _T_18065_45 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_14747) begin
                                                                  _T_18065_45 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_14745) begin
                                                                    _T_18065_45 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_14743) begin
                                                                      _T_18065_45 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_14741) begin
                                                                        _T_18065_45 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_14739) begin
                                                                          _T_18065_45 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_14737) begin
                                                                            _T_18065_45 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_14735) begin
                                                                              _T_18065_45 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_14733) begin
                                                                                _T_18065_45 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_14731) begin
                                                                                  _T_18065_45 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_14729) begin
                                                                                    _T_18065_45 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_14727) begin
                                                                                      _T_18065_45 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_14725) begin
                                                                                        _T_18065_45 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_14723) begin
                                                                                          _T_18065_45 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_14721) begin
                                                                                            _T_18065_45 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_14719) begin
                                                                                              _T_18065_45 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_14717) begin
                                                                                                _T_18065_45 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_14715) begin
                                                                                                  _T_18065_45 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_14713) begin
                                                                                                    _T_18065_45 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    _T_18065_45 <= 8'h0;
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_45 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_46) begin
        if (_T_14945) begin
          _T_18065_46 <= _T_10366_0;
        end else begin
          if (_T_14943) begin
            _T_18065_46 <= _T_10366_1;
          end else begin
            if (_T_14941) begin
              _T_18065_46 <= _T_10366_2;
            end else begin
              if (_T_14939) begin
                _T_18065_46 <= _T_10366_3;
              end else begin
                if (_T_14937) begin
                  _T_18065_46 <= _T_10366_4;
                end else begin
                  if (_T_14935) begin
                    _T_18065_46 <= _T_10366_5;
                  end else begin
                    if (_T_14933) begin
                      _T_18065_46 <= _T_10366_6;
                    end else begin
                      if (_T_14931) begin
                        _T_18065_46 <= _T_10366_7;
                      end else begin
                        if (_T_14929) begin
                          _T_18065_46 <= _T_10366_8;
                        end else begin
                          if (_T_14927) begin
                            _T_18065_46 <= _T_10366_9;
                          end else begin
                            if (_T_14925) begin
                              _T_18065_46 <= _T_10366_10;
                            end else begin
                              if (_T_14923) begin
                                _T_18065_46 <= _T_10366_11;
                              end else begin
                                if (_T_14921) begin
                                  _T_18065_46 <= _T_10366_12;
                                end else begin
                                  if (_T_14919) begin
                                    _T_18065_46 <= _T_10366_13;
                                  end else begin
                                    if (_T_14917) begin
                                      _T_18065_46 <= _T_10366_14;
                                    end else begin
                                      if (_T_14915) begin
                                        _T_18065_46 <= _T_10366_15;
                                      end else begin
                                        if (_T_14913) begin
                                          _T_18065_46 <= _T_10366_16;
                                        end else begin
                                          if (_T_14911) begin
                                            _T_18065_46 <= _T_10366_17;
                                          end else begin
                                            if (_T_14909) begin
                                              _T_18065_46 <= _T_10366_18;
                                            end else begin
                                              if (_T_14907) begin
                                                _T_18065_46 <= _T_10366_19;
                                              end else begin
                                                if (_T_14905) begin
                                                  _T_18065_46 <= _T_10366_20;
                                                end else begin
                                                  if (_T_14903) begin
                                                    _T_18065_46 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_14901) begin
                                                      _T_18065_46 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_14899) begin
                                                        _T_18065_46 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_14897) begin
                                                          _T_18065_46 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_14895) begin
                                                            _T_18065_46 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_14893) begin
                                                              _T_18065_46 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_14891) begin
                                                                _T_18065_46 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_14889) begin
                                                                  _T_18065_46 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_14887) begin
                                                                    _T_18065_46 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_14885) begin
                                                                      _T_18065_46 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_14883) begin
                                                                        _T_18065_46 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_14881) begin
                                                                          _T_18065_46 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_14879) begin
                                                                            _T_18065_46 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_14877) begin
                                                                              _T_18065_46 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_14875) begin
                                                                                _T_18065_46 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_14873) begin
                                                                                  _T_18065_46 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_14871) begin
                                                                                    _T_18065_46 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_14869) begin
                                                                                      _T_18065_46 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_14867) begin
                                                                                        _T_18065_46 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_14865) begin
                                                                                          _T_18065_46 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_14863) begin
                                                                                            _T_18065_46 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_14861) begin
                                                                                              _T_18065_46 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_14859) begin
                                                                                                _T_18065_46 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_14857) begin
                                                                                                  _T_18065_46 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_14855) begin
                                                                                                    _T_18065_46 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_14853) begin
                                                                                                      _T_18065_46 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      _T_18065_46 <= 8'h0;
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_46 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_47) begin
        if (_T_15090) begin
          _T_18065_47 <= _T_10366_0;
        end else begin
          if (_T_15088) begin
            _T_18065_47 <= _T_10366_1;
          end else begin
            if (_T_15086) begin
              _T_18065_47 <= _T_10366_2;
            end else begin
              if (_T_15084) begin
                _T_18065_47 <= _T_10366_3;
              end else begin
                if (_T_15082) begin
                  _T_18065_47 <= _T_10366_4;
                end else begin
                  if (_T_15080) begin
                    _T_18065_47 <= _T_10366_5;
                  end else begin
                    if (_T_15078) begin
                      _T_18065_47 <= _T_10366_6;
                    end else begin
                      if (_T_15076) begin
                        _T_18065_47 <= _T_10366_7;
                      end else begin
                        if (_T_15074) begin
                          _T_18065_47 <= _T_10366_8;
                        end else begin
                          if (_T_15072) begin
                            _T_18065_47 <= _T_10366_9;
                          end else begin
                            if (_T_15070) begin
                              _T_18065_47 <= _T_10366_10;
                            end else begin
                              if (_T_15068) begin
                                _T_18065_47 <= _T_10366_11;
                              end else begin
                                if (_T_15066) begin
                                  _T_18065_47 <= _T_10366_12;
                                end else begin
                                  if (_T_15064) begin
                                    _T_18065_47 <= _T_10366_13;
                                  end else begin
                                    if (_T_15062) begin
                                      _T_18065_47 <= _T_10366_14;
                                    end else begin
                                      if (_T_15060) begin
                                        _T_18065_47 <= _T_10366_15;
                                      end else begin
                                        if (_T_15058) begin
                                          _T_18065_47 <= _T_10366_16;
                                        end else begin
                                          if (_T_15056) begin
                                            _T_18065_47 <= _T_10366_17;
                                          end else begin
                                            if (_T_15054) begin
                                              _T_18065_47 <= _T_10366_18;
                                            end else begin
                                              if (_T_15052) begin
                                                _T_18065_47 <= _T_10366_19;
                                              end else begin
                                                if (_T_15050) begin
                                                  _T_18065_47 <= _T_10366_20;
                                                end else begin
                                                  if (_T_15048) begin
                                                    _T_18065_47 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_15046) begin
                                                      _T_18065_47 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_15044) begin
                                                        _T_18065_47 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_15042) begin
                                                          _T_18065_47 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_15040) begin
                                                            _T_18065_47 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_15038) begin
                                                              _T_18065_47 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_15036) begin
                                                                _T_18065_47 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_15034) begin
                                                                  _T_18065_47 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_15032) begin
                                                                    _T_18065_47 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_15030) begin
                                                                      _T_18065_47 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_15028) begin
                                                                        _T_18065_47 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_15026) begin
                                                                          _T_18065_47 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_15024) begin
                                                                            _T_18065_47 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_15022) begin
                                                                              _T_18065_47 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_15020) begin
                                                                                _T_18065_47 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_15018) begin
                                                                                  _T_18065_47 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_15016) begin
                                                                                    _T_18065_47 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_15014) begin
                                                                                      _T_18065_47 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_15012) begin
                                                                                        _T_18065_47 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_15010) begin
                                                                                          _T_18065_47 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_15008) begin
                                                                                            _T_18065_47 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_15006) begin
                                                                                              _T_18065_47 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_15004) begin
                                                                                                _T_18065_47 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_15002) begin
                                                                                                  _T_18065_47 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_15000) begin
                                                                                                    _T_18065_47 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_14998) begin
                                                                                                      _T_18065_47 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_14996) begin
                                                                                                        _T_18065_47 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        _T_18065_47 <= 8'h0;
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_47 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_48) begin
        if (_T_15238) begin
          _T_18065_48 <= _T_10366_0;
        end else begin
          if (_T_15236) begin
            _T_18065_48 <= _T_10366_1;
          end else begin
            if (_T_15234) begin
              _T_18065_48 <= _T_10366_2;
            end else begin
              if (_T_15232) begin
                _T_18065_48 <= _T_10366_3;
              end else begin
                if (_T_15230) begin
                  _T_18065_48 <= _T_10366_4;
                end else begin
                  if (_T_15228) begin
                    _T_18065_48 <= _T_10366_5;
                  end else begin
                    if (_T_15226) begin
                      _T_18065_48 <= _T_10366_6;
                    end else begin
                      if (_T_15224) begin
                        _T_18065_48 <= _T_10366_7;
                      end else begin
                        if (_T_15222) begin
                          _T_18065_48 <= _T_10366_8;
                        end else begin
                          if (_T_15220) begin
                            _T_18065_48 <= _T_10366_9;
                          end else begin
                            if (_T_15218) begin
                              _T_18065_48 <= _T_10366_10;
                            end else begin
                              if (_T_15216) begin
                                _T_18065_48 <= _T_10366_11;
                              end else begin
                                if (_T_15214) begin
                                  _T_18065_48 <= _T_10366_12;
                                end else begin
                                  if (_T_15212) begin
                                    _T_18065_48 <= _T_10366_13;
                                  end else begin
                                    if (_T_15210) begin
                                      _T_18065_48 <= _T_10366_14;
                                    end else begin
                                      if (_T_15208) begin
                                        _T_18065_48 <= _T_10366_15;
                                      end else begin
                                        if (_T_15206) begin
                                          _T_18065_48 <= _T_10366_16;
                                        end else begin
                                          if (_T_15204) begin
                                            _T_18065_48 <= _T_10366_17;
                                          end else begin
                                            if (_T_15202) begin
                                              _T_18065_48 <= _T_10366_18;
                                            end else begin
                                              if (_T_15200) begin
                                                _T_18065_48 <= _T_10366_19;
                                              end else begin
                                                if (_T_15198) begin
                                                  _T_18065_48 <= _T_10366_20;
                                                end else begin
                                                  if (_T_15196) begin
                                                    _T_18065_48 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_15194) begin
                                                      _T_18065_48 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_15192) begin
                                                        _T_18065_48 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_15190) begin
                                                          _T_18065_48 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_15188) begin
                                                            _T_18065_48 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_15186) begin
                                                              _T_18065_48 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_15184) begin
                                                                _T_18065_48 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_15182) begin
                                                                  _T_18065_48 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_15180) begin
                                                                    _T_18065_48 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_15178) begin
                                                                      _T_18065_48 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_15176) begin
                                                                        _T_18065_48 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_15174) begin
                                                                          _T_18065_48 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_15172) begin
                                                                            _T_18065_48 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_15170) begin
                                                                              _T_18065_48 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_15168) begin
                                                                                _T_18065_48 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_15166) begin
                                                                                  _T_18065_48 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_15164) begin
                                                                                    _T_18065_48 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_15162) begin
                                                                                      _T_18065_48 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_15160) begin
                                                                                        _T_18065_48 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_15158) begin
                                                                                          _T_18065_48 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_15156) begin
                                                                                            _T_18065_48 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_15154) begin
                                                                                              _T_18065_48 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_15152) begin
                                                                                                _T_18065_48 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_15150) begin
                                                                                                  _T_18065_48 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_15148) begin
                                                                                                    _T_18065_48 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_15146) begin
                                                                                                      _T_18065_48 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_15144) begin
                                                                                                        _T_18065_48 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_15142) begin
                                                                                                          _T_18065_48 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          _T_18065_48 <= 8'h0;
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_48 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_49) begin
        if (_T_15389) begin
          _T_18065_49 <= _T_10366_0;
        end else begin
          if (_T_15387) begin
            _T_18065_49 <= _T_10366_1;
          end else begin
            if (_T_15385) begin
              _T_18065_49 <= _T_10366_2;
            end else begin
              if (_T_15383) begin
                _T_18065_49 <= _T_10366_3;
              end else begin
                if (_T_15381) begin
                  _T_18065_49 <= _T_10366_4;
                end else begin
                  if (_T_15379) begin
                    _T_18065_49 <= _T_10366_5;
                  end else begin
                    if (_T_15377) begin
                      _T_18065_49 <= _T_10366_6;
                    end else begin
                      if (_T_15375) begin
                        _T_18065_49 <= _T_10366_7;
                      end else begin
                        if (_T_15373) begin
                          _T_18065_49 <= _T_10366_8;
                        end else begin
                          if (_T_15371) begin
                            _T_18065_49 <= _T_10366_9;
                          end else begin
                            if (_T_15369) begin
                              _T_18065_49 <= _T_10366_10;
                            end else begin
                              if (_T_15367) begin
                                _T_18065_49 <= _T_10366_11;
                              end else begin
                                if (_T_15365) begin
                                  _T_18065_49 <= _T_10366_12;
                                end else begin
                                  if (_T_15363) begin
                                    _T_18065_49 <= _T_10366_13;
                                  end else begin
                                    if (_T_15361) begin
                                      _T_18065_49 <= _T_10366_14;
                                    end else begin
                                      if (_T_15359) begin
                                        _T_18065_49 <= _T_10366_15;
                                      end else begin
                                        if (_T_15357) begin
                                          _T_18065_49 <= _T_10366_16;
                                        end else begin
                                          if (_T_15355) begin
                                            _T_18065_49 <= _T_10366_17;
                                          end else begin
                                            if (_T_15353) begin
                                              _T_18065_49 <= _T_10366_18;
                                            end else begin
                                              if (_T_15351) begin
                                                _T_18065_49 <= _T_10366_19;
                                              end else begin
                                                if (_T_15349) begin
                                                  _T_18065_49 <= _T_10366_20;
                                                end else begin
                                                  if (_T_15347) begin
                                                    _T_18065_49 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_15345) begin
                                                      _T_18065_49 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_15343) begin
                                                        _T_18065_49 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_15341) begin
                                                          _T_18065_49 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_15339) begin
                                                            _T_18065_49 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_15337) begin
                                                              _T_18065_49 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_15335) begin
                                                                _T_18065_49 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_15333) begin
                                                                  _T_18065_49 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_15331) begin
                                                                    _T_18065_49 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_15329) begin
                                                                      _T_18065_49 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_15327) begin
                                                                        _T_18065_49 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_15325) begin
                                                                          _T_18065_49 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_15323) begin
                                                                            _T_18065_49 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_15321) begin
                                                                              _T_18065_49 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_15319) begin
                                                                                _T_18065_49 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_15317) begin
                                                                                  _T_18065_49 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_15315) begin
                                                                                    _T_18065_49 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_15313) begin
                                                                                      _T_18065_49 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_15311) begin
                                                                                        _T_18065_49 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_15309) begin
                                                                                          _T_18065_49 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_15307) begin
                                                                                            _T_18065_49 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_15305) begin
                                                                                              _T_18065_49 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_15303) begin
                                                                                                _T_18065_49 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_15301) begin
                                                                                                  _T_18065_49 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_15299) begin
                                                                                                    _T_18065_49 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_15297) begin
                                                                                                      _T_18065_49 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_15295) begin
                                                                                                        _T_18065_49 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_15293) begin
                                                                                                          _T_18065_49 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_15291) begin
                                                                                                            _T_18065_49 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            _T_18065_49 <= 8'h0;
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_49 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_50) begin
        if (_T_15543) begin
          _T_18065_50 <= _T_10366_0;
        end else begin
          if (_T_15541) begin
            _T_18065_50 <= _T_10366_1;
          end else begin
            if (_T_15539) begin
              _T_18065_50 <= _T_10366_2;
            end else begin
              if (_T_15537) begin
                _T_18065_50 <= _T_10366_3;
              end else begin
                if (_T_15535) begin
                  _T_18065_50 <= _T_10366_4;
                end else begin
                  if (_T_15533) begin
                    _T_18065_50 <= _T_10366_5;
                  end else begin
                    if (_T_15531) begin
                      _T_18065_50 <= _T_10366_6;
                    end else begin
                      if (_T_15529) begin
                        _T_18065_50 <= _T_10366_7;
                      end else begin
                        if (_T_15527) begin
                          _T_18065_50 <= _T_10366_8;
                        end else begin
                          if (_T_15525) begin
                            _T_18065_50 <= _T_10366_9;
                          end else begin
                            if (_T_15523) begin
                              _T_18065_50 <= _T_10366_10;
                            end else begin
                              if (_T_15521) begin
                                _T_18065_50 <= _T_10366_11;
                              end else begin
                                if (_T_15519) begin
                                  _T_18065_50 <= _T_10366_12;
                                end else begin
                                  if (_T_15517) begin
                                    _T_18065_50 <= _T_10366_13;
                                  end else begin
                                    if (_T_15515) begin
                                      _T_18065_50 <= _T_10366_14;
                                    end else begin
                                      if (_T_15513) begin
                                        _T_18065_50 <= _T_10366_15;
                                      end else begin
                                        if (_T_15511) begin
                                          _T_18065_50 <= _T_10366_16;
                                        end else begin
                                          if (_T_15509) begin
                                            _T_18065_50 <= _T_10366_17;
                                          end else begin
                                            if (_T_15507) begin
                                              _T_18065_50 <= _T_10366_18;
                                            end else begin
                                              if (_T_15505) begin
                                                _T_18065_50 <= _T_10366_19;
                                              end else begin
                                                if (_T_15503) begin
                                                  _T_18065_50 <= _T_10366_20;
                                                end else begin
                                                  if (_T_15501) begin
                                                    _T_18065_50 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_15499) begin
                                                      _T_18065_50 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_15497) begin
                                                        _T_18065_50 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_15495) begin
                                                          _T_18065_50 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_15493) begin
                                                            _T_18065_50 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_15491) begin
                                                              _T_18065_50 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_15489) begin
                                                                _T_18065_50 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_15487) begin
                                                                  _T_18065_50 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_15485) begin
                                                                    _T_18065_50 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_15483) begin
                                                                      _T_18065_50 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_15481) begin
                                                                        _T_18065_50 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_15479) begin
                                                                          _T_18065_50 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_15477) begin
                                                                            _T_18065_50 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_15475) begin
                                                                              _T_18065_50 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_15473) begin
                                                                                _T_18065_50 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_15471) begin
                                                                                  _T_18065_50 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_15469) begin
                                                                                    _T_18065_50 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_15467) begin
                                                                                      _T_18065_50 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_15465) begin
                                                                                        _T_18065_50 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_15463) begin
                                                                                          _T_18065_50 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_15461) begin
                                                                                            _T_18065_50 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_15459) begin
                                                                                              _T_18065_50 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_15457) begin
                                                                                                _T_18065_50 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_15455) begin
                                                                                                  _T_18065_50 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_15453) begin
                                                                                                    _T_18065_50 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_15451) begin
                                                                                                      _T_18065_50 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_15449) begin
                                                                                                        _T_18065_50 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_15447) begin
                                                                                                          _T_18065_50 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_15445) begin
                                                                                                            _T_18065_50 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_15443) begin
                                                                                                              _T_18065_50 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              _T_18065_50 <= 8'h0;
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_50 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_51) begin
        if (_T_15700) begin
          _T_18065_51 <= _T_10366_0;
        end else begin
          if (_T_15698) begin
            _T_18065_51 <= _T_10366_1;
          end else begin
            if (_T_15696) begin
              _T_18065_51 <= _T_10366_2;
            end else begin
              if (_T_15694) begin
                _T_18065_51 <= _T_10366_3;
              end else begin
                if (_T_15692) begin
                  _T_18065_51 <= _T_10366_4;
                end else begin
                  if (_T_15690) begin
                    _T_18065_51 <= _T_10366_5;
                  end else begin
                    if (_T_15688) begin
                      _T_18065_51 <= _T_10366_6;
                    end else begin
                      if (_T_15686) begin
                        _T_18065_51 <= _T_10366_7;
                      end else begin
                        if (_T_15684) begin
                          _T_18065_51 <= _T_10366_8;
                        end else begin
                          if (_T_15682) begin
                            _T_18065_51 <= _T_10366_9;
                          end else begin
                            if (_T_15680) begin
                              _T_18065_51 <= _T_10366_10;
                            end else begin
                              if (_T_15678) begin
                                _T_18065_51 <= _T_10366_11;
                              end else begin
                                if (_T_15676) begin
                                  _T_18065_51 <= _T_10366_12;
                                end else begin
                                  if (_T_15674) begin
                                    _T_18065_51 <= _T_10366_13;
                                  end else begin
                                    if (_T_15672) begin
                                      _T_18065_51 <= _T_10366_14;
                                    end else begin
                                      if (_T_15670) begin
                                        _T_18065_51 <= _T_10366_15;
                                      end else begin
                                        if (_T_15668) begin
                                          _T_18065_51 <= _T_10366_16;
                                        end else begin
                                          if (_T_15666) begin
                                            _T_18065_51 <= _T_10366_17;
                                          end else begin
                                            if (_T_15664) begin
                                              _T_18065_51 <= _T_10366_18;
                                            end else begin
                                              if (_T_15662) begin
                                                _T_18065_51 <= _T_10366_19;
                                              end else begin
                                                if (_T_15660) begin
                                                  _T_18065_51 <= _T_10366_20;
                                                end else begin
                                                  if (_T_15658) begin
                                                    _T_18065_51 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_15656) begin
                                                      _T_18065_51 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_15654) begin
                                                        _T_18065_51 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_15652) begin
                                                          _T_18065_51 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_15650) begin
                                                            _T_18065_51 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_15648) begin
                                                              _T_18065_51 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_15646) begin
                                                                _T_18065_51 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_15644) begin
                                                                  _T_18065_51 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_15642) begin
                                                                    _T_18065_51 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_15640) begin
                                                                      _T_18065_51 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_15638) begin
                                                                        _T_18065_51 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_15636) begin
                                                                          _T_18065_51 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_15634) begin
                                                                            _T_18065_51 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_15632) begin
                                                                              _T_18065_51 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_15630) begin
                                                                                _T_18065_51 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_15628) begin
                                                                                  _T_18065_51 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_15626) begin
                                                                                    _T_18065_51 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_15624) begin
                                                                                      _T_18065_51 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_15622) begin
                                                                                        _T_18065_51 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_15620) begin
                                                                                          _T_18065_51 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_15618) begin
                                                                                            _T_18065_51 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_15616) begin
                                                                                              _T_18065_51 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_15614) begin
                                                                                                _T_18065_51 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_15612) begin
                                                                                                  _T_18065_51 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_15610) begin
                                                                                                    _T_18065_51 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_15608) begin
                                                                                                      _T_18065_51 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_15606) begin
                                                                                                        _T_18065_51 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_15604) begin
                                                                                                          _T_18065_51 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_15602) begin
                                                                                                            _T_18065_51 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_15600) begin
                                                                                                              _T_18065_51 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_15598) begin
                                                                                                                _T_18065_51 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                _T_18065_51 <= 8'h0;
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_51 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_52) begin
        if (_T_15860) begin
          _T_18065_52 <= _T_10366_0;
        end else begin
          if (_T_15858) begin
            _T_18065_52 <= _T_10366_1;
          end else begin
            if (_T_15856) begin
              _T_18065_52 <= _T_10366_2;
            end else begin
              if (_T_15854) begin
                _T_18065_52 <= _T_10366_3;
              end else begin
                if (_T_15852) begin
                  _T_18065_52 <= _T_10366_4;
                end else begin
                  if (_T_15850) begin
                    _T_18065_52 <= _T_10366_5;
                  end else begin
                    if (_T_15848) begin
                      _T_18065_52 <= _T_10366_6;
                    end else begin
                      if (_T_15846) begin
                        _T_18065_52 <= _T_10366_7;
                      end else begin
                        if (_T_15844) begin
                          _T_18065_52 <= _T_10366_8;
                        end else begin
                          if (_T_15842) begin
                            _T_18065_52 <= _T_10366_9;
                          end else begin
                            if (_T_15840) begin
                              _T_18065_52 <= _T_10366_10;
                            end else begin
                              if (_T_15838) begin
                                _T_18065_52 <= _T_10366_11;
                              end else begin
                                if (_T_15836) begin
                                  _T_18065_52 <= _T_10366_12;
                                end else begin
                                  if (_T_15834) begin
                                    _T_18065_52 <= _T_10366_13;
                                  end else begin
                                    if (_T_15832) begin
                                      _T_18065_52 <= _T_10366_14;
                                    end else begin
                                      if (_T_15830) begin
                                        _T_18065_52 <= _T_10366_15;
                                      end else begin
                                        if (_T_15828) begin
                                          _T_18065_52 <= _T_10366_16;
                                        end else begin
                                          if (_T_15826) begin
                                            _T_18065_52 <= _T_10366_17;
                                          end else begin
                                            if (_T_15824) begin
                                              _T_18065_52 <= _T_10366_18;
                                            end else begin
                                              if (_T_15822) begin
                                                _T_18065_52 <= _T_10366_19;
                                              end else begin
                                                if (_T_15820) begin
                                                  _T_18065_52 <= _T_10366_20;
                                                end else begin
                                                  if (_T_15818) begin
                                                    _T_18065_52 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_15816) begin
                                                      _T_18065_52 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_15814) begin
                                                        _T_18065_52 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_15812) begin
                                                          _T_18065_52 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_15810) begin
                                                            _T_18065_52 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_15808) begin
                                                              _T_18065_52 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_15806) begin
                                                                _T_18065_52 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_15804) begin
                                                                  _T_18065_52 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_15802) begin
                                                                    _T_18065_52 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_15800) begin
                                                                      _T_18065_52 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_15798) begin
                                                                        _T_18065_52 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_15796) begin
                                                                          _T_18065_52 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_15794) begin
                                                                            _T_18065_52 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_15792) begin
                                                                              _T_18065_52 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_15790) begin
                                                                                _T_18065_52 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_15788) begin
                                                                                  _T_18065_52 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_15786) begin
                                                                                    _T_18065_52 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_15784) begin
                                                                                      _T_18065_52 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_15782) begin
                                                                                        _T_18065_52 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_15780) begin
                                                                                          _T_18065_52 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_15778) begin
                                                                                            _T_18065_52 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_15776) begin
                                                                                              _T_18065_52 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_15774) begin
                                                                                                _T_18065_52 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_15772) begin
                                                                                                  _T_18065_52 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_15770) begin
                                                                                                    _T_18065_52 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_15768) begin
                                                                                                      _T_18065_52 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_15766) begin
                                                                                                        _T_18065_52 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_15764) begin
                                                                                                          _T_18065_52 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_15762) begin
                                                                                                            _T_18065_52 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_15760) begin
                                                                                                              _T_18065_52 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_15758) begin
                                                                                                                _T_18065_52 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_15756) begin
                                                                                                                  _T_18065_52 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  _T_18065_52 <= 8'h0;
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_52 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_53) begin
        if (_T_16023) begin
          _T_18065_53 <= _T_10366_0;
        end else begin
          if (_T_16021) begin
            _T_18065_53 <= _T_10366_1;
          end else begin
            if (_T_16019) begin
              _T_18065_53 <= _T_10366_2;
            end else begin
              if (_T_16017) begin
                _T_18065_53 <= _T_10366_3;
              end else begin
                if (_T_16015) begin
                  _T_18065_53 <= _T_10366_4;
                end else begin
                  if (_T_16013) begin
                    _T_18065_53 <= _T_10366_5;
                  end else begin
                    if (_T_16011) begin
                      _T_18065_53 <= _T_10366_6;
                    end else begin
                      if (_T_16009) begin
                        _T_18065_53 <= _T_10366_7;
                      end else begin
                        if (_T_16007) begin
                          _T_18065_53 <= _T_10366_8;
                        end else begin
                          if (_T_16005) begin
                            _T_18065_53 <= _T_10366_9;
                          end else begin
                            if (_T_16003) begin
                              _T_18065_53 <= _T_10366_10;
                            end else begin
                              if (_T_16001) begin
                                _T_18065_53 <= _T_10366_11;
                              end else begin
                                if (_T_15999) begin
                                  _T_18065_53 <= _T_10366_12;
                                end else begin
                                  if (_T_15997) begin
                                    _T_18065_53 <= _T_10366_13;
                                  end else begin
                                    if (_T_15995) begin
                                      _T_18065_53 <= _T_10366_14;
                                    end else begin
                                      if (_T_15993) begin
                                        _T_18065_53 <= _T_10366_15;
                                      end else begin
                                        if (_T_15991) begin
                                          _T_18065_53 <= _T_10366_16;
                                        end else begin
                                          if (_T_15989) begin
                                            _T_18065_53 <= _T_10366_17;
                                          end else begin
                                            if (_T_15987) begin
                                              _T_18065_53 <= _T_10366_18;
                                            end else begin
                                              if (_T_15985) begin
                                                _T_18065_53 <= _T_10366_19;
                                              end else begin
                                                if (_T_15983) begin
                                                  _T_18065_53 <= _T_10366_20;
                                                end else begin
                                                  if (_T_15981) begin
                                                    _T_18065_53 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_15979) begin
                                                      _T_18065_53 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_15977) begin
                                                        _T_18065_53 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_15975) begin
                                                          _T_18065_53 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_15973) begin
                                                            _T_18065_53 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_15971) begin
                                                              _T_18065_53 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_15969) begin
                                                                _T_18065_53 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_15967) begin
                                                                  _T_18065_53 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_15965) begin
                                                                    _T_18065_53 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_15963) begin
                                                                      _T_18065_53 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_15961) begin
                                                                        _T_18065_53 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_15959) begin
                                                                          _T_18065_53 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_15957) begin
                                                                            _T_18065_53 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_15955) begin
                                                                              _T_18065_53 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_15953) begin
                                                                                _T_18065_53 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_15951) begin
                                                                                  _T_18065_53 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_15949) begin
                                                                                    _T_18065_53 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_15947) begin
                                                                                      _T_18065_53 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_15945) begin
                                                                                        _T_18065_53 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_15943) begin
                                                                                          _T_18065_53 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_15941) begin
                                                                                            _T_18065_53 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_15939) begin
                                                                                              _T_18065_53 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_15937) begin
                                                                                                _T_18065_53 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_15935) begin
                                                                                                  _T_18065_53 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_15933) begin
                                                                                                    _T_18065_53 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_15931) begin
                                                                                                      _T_18065_53 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_15929) begin
                                                                                                        _T_18065_53 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_15927) begin
                                                                                                          _T_18065_53 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_15925) begin
                                                                                                            _T_18065_53 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_15923) begin
                                                                                                              _T_18065_53 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_15921) begin
                                                                                                                _T_18065_53 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_15919) begin
                                                                                                                  _T_18065_53 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_15917) begin
                                                                                                                    _T_18065_53 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    _T_18065_53 <= 8'h0;
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_53 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_54) begin
        if (_T_16189) begin
          _T_18065_54 <= _T_10366_0;
        end else begin
          if (_T_16187) begin
            _T_18065_54 <= _T_10366_1;
          end else begin
            if (_T_16185) begin
              _T_18065_54 <= _T_10366_2;
            end else begin
              if (_T_16183) begin
                _T_18065_54 <= _T_10366_3;
              end else begin
                if (_T_16181) begin
                  _T_18065_54 <= _T_10366_4;
                end else begin
                  if (_T_16179) begin
                    _T_18065_54 <= _T_10366_5;
                  end else begin
                    if (_T_16177) begin
                      _T_18065_54 <= _T_10366_6;
                    end else begin
                      if (_T_16175) begin
                        _T_18065_54 <= _T_10366_7;
                      end else begin
                        if (_T_16173) begin
                          _T_18065_54 <= _T_10366_8;
                        end else begin
                          if (_T_16171) begin
                            _T_18065_54 <= _T_10366_9;
                          end else begin
                            if (_T_16169) begin
                              _T_18065_54 <= _T_10366_10;
                            end else begin
                              if (_T_16167) begin
                                _T_18065_54 <= _T_10366_11;
                              end else begin
                                if (_T_16165) begin
                                  _T_18065_54 <= _T_10366_12;
                                end else begin
                                  if (_T_16163) begin
                                    _T_18065_54 <= _T_10366_13;
                                  end else begin
                                    if (_T_16161) begin
                                      _T_18065_54 <= _T_10366_14;
                                    end else begin
                                      if (_T_16159) begin
                                        _T_18065_54 <= _T_10366_15;
                                      end else begin
                                        if (_T_16157) begin
                                          _T_18065_54 <= _T_10366_16;
                                        end else begin
                                          if (_T_16155) begin
                                            _T_18065_54 <= _T_10366_17;
                                          end else begin
                                            if (_T_16153) begin
                                              _T_18065_54 <= _T_10366_18;
                                            end else begin
                                              if (_T_16151) begin
                                                _T_18065_54 <= _T_10366_19;
                                              end else begin
                                                if (_T_16149) begin
                                                  _T_18065_54 <= _T_10366_20;
                                                end else begin
                                                  if (_T_16147) begin
                                                    _T_18065_54 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_16145) begin
                                                      _T_18065_54 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_16143) begin
                                                        _T_18065_54 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_16141) begin
                                                          _T_18065_54 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_16139) begin
                                                            _T_18065_54 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_16137) begin
                                                              _T_18065_54 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_16135) begin
                                                                _T_18065_54 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_16133) begin
                                                                  _T_18065_54 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_16131) begin
                                                                    _T_18065_54 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_16129) begin
                                                                      _T_18065_54 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_16127) begin
                                                                        _T_18065_54 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_16125) begin
                                                                          _T_18065_54 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_16123) begin
                                                                            _T_18065_54 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_16121) begin
                                                                              _T_18065_54 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_16119) begin
                                                                                _T_18065_54 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_16117) begin
                                                                                  _T_18065_54 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_16115) begin
                                                                                    _T_18065_54 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_16113) begin
                                                                                      _T_18065_54 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_16111) begin
                                                                                        _T_18065_54 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_16109) begin
                                                                                          _T_18065_54 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_16107) begin
                                                                                            _T_18065_54 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_16105) begin
                                                                                              _T_18065_54 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_16103) begin
                                                                                                _T_18065_54 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_16101) begin
                                                                                                  _T_18065_54 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_16099) begin
                                                                                                    _T_18065_54 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_16097) begin
                                                                                                      _T_18065_54 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_16095) begin
                                                                                                        _T_18065_54 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_16093) begin
                                                                                                          _T_18065_54 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_16091) begin
                                                                                                            _T_18065_54 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_16089) begin
                                                                                                              _T_18065_54 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_16087) begin
                                                                                                                _T_18065_54 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_16085) begin
                                                                                                                  _T_18065_54 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_16083) begin
                                                                                                                    _T_18065_54 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_16081) begin
                                                                                                                      _T_18065_54 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      _T_18065_54 <= 8'h0;
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_54 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_55) begin
        if (_T_16358) begin
          _T_18065_55 <= _T_10366_0;
        end else begin
          if (_T_16356) begin
            _T_18065_55 <= _T_10366_1;
          end else begin
            if (_T_16354) begin
              _T_18065_55 <= _T_10366_2;
            end else begin
              if (_T_16352) begin
                _T_18065_55 <= _T_10366_3;
              end else begin
                if (_T_16350) begin
                  _T_18065_55 <= _T_10366_4;
                end else begin
                  if (_T_16348) begin
                    _T_18065_55 <= _T_10366_5;
                  end else begin
                    if (_T_16346) begin
                      _T_18065_55 <= _T_10366_6;
                    end else begin
                      if (_T_16344) begin
                        _T_18065_55 <= _T_10366_7;
                      end else begin
                        if (_T_16342) begin
                          _T_18065_55 <= _T_10366_8;
                        end else begin
                          if (_T_16340) begin
                            _T_18065_55 <= _T_10366_9;
                          end else begin
                            if (_T_16338) begin
                              _T_18065_55 <= _T_10366_10;
                            end else begin
                              if (_T_16336) begin
                                _T_18065_55 <= _T_10366_11;
                              end else begin
                                if (_T_16334) begin
                                  _T_18065_55 <= _T_10366_12;
                                end else begin
                                  if (_T_16332) begin
                                    _T_18065_55 <= _T_10366_13;
                                  end else begin
                                    if (_T_16330) begin
                                      _T_18065_55 <= _T_10366_14;
                                    end else begin
                                      if (_T_16328) begin
                                        _T_18065_55 <= _T_10366_15;
                                      end else begin
                                        if (_T_16326) begin
                                          _T_18065_55 <= _T_10366_16;
                                        end else begin
                                          if (_T_16324) begin
                                            _T_18065_55 <= _T_10366_17;
                                          end else begin
                                            if (_T_16322) begin
                                              _T_18065_55 <= _T_10366_18;
                                            end else begin
                                              if (_T_16320) begin
                                                _T_18065_55 <= _T_10366_19;
                                              end else begin
                                                if (_T_16318) begin
                                                  _T_18065_55 <= _T_10366_20;
                                                end else begin
                                                  if (_T_16316) begin
                                                    _T_18065_55 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_16314) begin
                                                      _T_18065_55 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_16312) begin
                                                        _T_18065_55 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_16310) begin
                                                          _T_18065_55 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_16308) begin
                                                            _T_18065_55 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_16306) begin
                                                              _T_18065_55 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_16304) begin
                                                                _T_18065_55 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_16302) begin
                                                                  _T_18065_55 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_16300) begin
                                                                    _T_18065_55 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_16298) begin
                                                                      _T_18065_55 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_16296) begin
                                                                        _T_18065_55 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_16294) begin
                                                                          _T_18065_55 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_16292) begin
                                                                            _T_18065_55 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_16290) begin
                                                                              _T_18065_55 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_16288) begin
                                                                                _T_18065_55 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_16286) begin
                                                                                  _T_18065_55 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_16284) begin
                                                                                    _T_18065_55 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_16282) begin
                                                                                      _T_18065_55 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_16280) begin
                                                                                        _T_18065_55 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_16278) begin
                                                                                          _T_18065_55 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_16276) begin
                                                                                            _T_18065_55 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_16274) begin
                                                                                              _T_18065_55 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_16272) begin
                                                                                                _T_18065_55 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_16270) begin
                                                                                                  _T_18065_55 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_16268) begin
                                                                                                    _T_18065_55 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_16266) begin
                                                                                                      _T_18065_55 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_16264) begin
                                                                                                        _T_18065_55 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_16262) begin
                                                                                                          _T_18065_55 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_16260) begin
                                                                                                            _T_18065_55 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_16258) begin
                                                                                                              _T_18065_55 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_16256) begin
                                                                                                                _T_18065_55 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_16254) begin
                                                                                                                  _T_18065_55 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_16252) begin
                                                                                                                    _T_18065_55 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_16250) begin
                                                                                                                      _T_18065_55 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_16248) begin
                                                                                                                        _T_18065_55 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        _T_18065_55 <= 8'h0;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_55 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_56) begin
        if (_T_16530) begin
          _T_18065_56 <= _T_10366_0;
        end else begin
          if (_T_16528) begin
            _T_18065_56 <= _T_10366_1;
          end else begin
            if (_T_16526) begin
              _T_18065_56 <= _T_10366_2;
            end else begin
              if (_T_16524) begin
                _T_18065_56 <= _T_10366_3;
              end else begin
                if (_T_16522) begin
                  _T_18065_56 <= _T_10366_4;
                end else begin
                  if (_T_16520) begin
                    _T_18065_56 <= _T_10366_5;
                  end else begin
                    if (_T_16518) begin
                      _T_18065_56 <= _T_10366_6;
                    end else begin
                      if (_T_16516) begin
                        _T_18065_56 <= _T_10366_7;
                      end else begin
                        if (_T_16514) begin
                          _T_18065_56 <= _T_10366_8;
                        end else begin
                          if (_T_16512) begin
                            _T_18065_56 <= _T_10366_9;
                          end else begin
                            if (_T_16510) begin
                              _T_18065_56 <= _T_10366_10;
                            end else begin
                              if (_T_16508) begin
                                _T_18065_56 <= _T_10366_11;
                              end else begin
                                if (_T_16506) begin
                                  _T_18065_56 <= _T_10366_12;
                                end else begin
                                  if (_T_16504) begin
                                    _T_18065_56 <= _T_10366_13;
                                  end else begin
                                    if (_T_16502) begin
                                      _T_18065_56 <= _T_10366_14;
                                    end else begin
                                      if (_T_16500) begin
                                        _T_18065_56 <= _T_10366_15;
                                      end else begin
                                        if (_T_16498) begin
                                          _T_18065_56 <= _T_10366_16;
                                        end else begin
                                          if (_T_16496) begin
                                            _T_18065_56 <= _T_10366_17;
                                          end else begin
                                            if (_T_16494) begin
                                              _T_18065_56 <= _T_10366_18;
                                            end else begin
                                              if (_T_16492) begin
                                                _T_18065_56 <= _T_10366_19;
                                              end else begin
                                                if (_T_16490) begin
                                                  _T_18065_56 <= _T_10366_20;
                                                end else begin
                                                  if (_T_16488) begin
                                                    _T_18065_56 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_16486) begin
                                                      _T_18065_56 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_16484) begin
                                                        _T_18065_56 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_16482) begin
                                                          _T_18065_56 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_16480) begin
                                                            _T_18065_56 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_16478) begin
                                                              _T_18065_56 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_16476) begin
                                                                _T_18065_56 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_16474) begin
                                                                  _T_18065_56 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_16472) begin
                                                                    _T_18065_56 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_16470) begin
                                                                      _T_18065_56 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_16468) begin
                                                                        _T_18065_56 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_16466) begin
                                                                          _T_18065_56 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_16464) begin
                                                                            _T_18065_56 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_16462) begin
                                                                              _T_18065_56 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_16460) begin
                                                                                _T_18065_56 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_16458) begin
                                                                                  _T_18065_56 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_16456) begin
                                                                                    _T_18065_56 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_16454) begin
                                                                                      _T_18065_56 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_16452) begin
                                                                                        _T_18065_56 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_16450) begin
                                                                                          _T_18065_56 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_16448) begin
                                                                                            _T_18065_56 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_16446) begin
                                                                                              _T_18065_56 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_16444) begin
                                                                                                _T_18065_56 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_16442) begin
                                                                                                  _T_18065_56 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_16440) begin
                                                                                                    _T_18065_56 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_16438) begin
                                                                                                      _T_18065_56 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_16436) begin
                                                                                                        _T_18065_56 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_16434) begin
                                                                                                          _T_18065_56 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_16432) begin
                                                                                                            _T_18065_56 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_16430) begin
                                                                                                              _T_18065_56 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_16428) begin
                                                                                                                _T_18065_56 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_16426) begin
                                                                                                                  _T_18065_56 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_16424) begin
                                                                                                                    _T_18065_56 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_16422) begin
                                                                                                                      _T_18065_56 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_16420) begin
                                                                                                                        _T_18065_56 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_16418) begin
                                                                                                                          _T_18065_56 <= _T_10366_56;
                                                                                                                        end else begin
                                                                                                                          _T_18065_56 <= 8'h0;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_56 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_57) begin
        if (_T_16705) begin
          _T_18065_57 <= _T_10366_0;
        end else begin
          if (_T_16703) begin
            _T_18065_57 <= _T_10366_1;
          end else begin
            if (_T_16701) begin
              _T_18065_57 <= _T_10366_2;
            end else begin
              if (_T_16699) begin
                _T_18065_57 <= _T_10366_3;
              end else begin
                if (_T_16697) begin
                  _T_18065_57 <= _T_10366_4;
                end else begin
                  if (_T_16695) begin
                    _T_18065_57 <= _T_10366_5;
                  end else begin
                    if (_T_16693) begin
                      _T_18065_57 <= _T_10366_6;
                    end else begin
                      if (_T_16691) begin
                        _T_18065_57 <= _T_10366_7;
                      end else begin
                        if (_T_16689) begin
                          _T_18065_57 <= _T_10366_8;
                        end else begin
                          if (_T_16687) begin
                            _T_18065_57 <= _T_10366_9;
                          end else begin
                            if (_T_16685) begin
                              _T_18065_57 <= _T_10366_10;
                            end else begin
                              if (_T_16683) begin
                                _T_18065_57 <= _T_10366_11;
                              end else begin
                                if (_T_16681) begin
                                  _T_18065_57 <= _T_10366_12;
                                end else begin
                                  if (_T_16679) begin
                                    _T_18065_57 <= _T_10366_13;
                                  end else begin
                                    if (_T_16677) begin
                                      _T_18065_57 <= _T_10366_14;
                                    end else begin
                                      if (_T_16675) begin
                                        _T_18065_57 <= _T_10366_15;
                                      end else begin
                                        if (_T_16673) begin
                                          _T_18065_57 <= _T_10366_16;
                                        end else begin
                                          if (_T_16671) begin
                                            _T_18065_57 <= _T_10366_17;
                                          end else begin
                                            if (_T_16669) begin
                                              _T_18065_57 <= _T_10366_18;
                                            end else begin
                                              if (_T_16667) begin
                                                _T_18065_57 <= _T_10366_19;
                                              end else begin
                                                if (_T_16665) begin
                                                  _T_18065_57 <= _T_10366_20;
                                                end else begin
                                                  if (_T_16663) begin
                                                    _T_18065_57 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_16661) begin
                                                      _T_18065_57 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_16659) begin
                                                        _T_18065_57 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_16657) begin
                                                          _T_18065_57 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_16655) begin
                                                            _T_18065_57 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_16653) begin
                                                              _T_18065_57 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_16651) begin
                                                                _T_18065_57 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_16649) begin
                                                                  _T_18065_57 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_16647) begin
                                                                    _T_18065_57 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_16645) begin
                                                                      _T_18065_57 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_16643) begin
                                                                        _T_18065_57 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_16641) begin
                                                                          _T_18065_57 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_16639) begin
                                                                            _T_18065_57 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_16637) begin
                                                                              _T_18065_57 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_16635) begin
                                                                                _T_18065_57 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_16633) begin
                                                                                  _T_18065_57 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_16631) begin
                                                                                    _T_18065_57 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_16629) begin
                                                                                      _T_18065_57 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_16627) begin
                                                                                        _T_18065_57 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_16625) begin
                                                                                          _T_18065_57 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_16623) begin
                                                                                            _T_18065_57 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_16621) begin
                                                                                              _T_18065_57 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_16619) begin
                                                                                                _T_18065_57 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_16617) begin
                                                                                                  _T_18065_57 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_16615) begin
                                                                                                    _T_18065_57 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_16613) begin
                                                                                                      _T_18065_57 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_16611) begin
                                                                                                        _T_18065_57 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_16609) begin
                                                                                                          _T_18065_57 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_16607) begin
                                                                                                            _T_18065_57 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_16605) begin
                                                                                                              _T_18065_57 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_16603) begin
                                                                                                                _T_18065_57 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_16601) begin
                                                                                                                  _T_18065_57 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_16599) begin
                                                                                                                    _T_18065_57 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_16597) begin
                                                                                                                      _T_18065_57 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_16595) begin
                                                                                                                        _T_18065_57 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_16593) begin
                                                                                                                          _T_18065_57 <= _T_10366_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_16591) begin
                                                                                                                            _T_18065_57 <= _T_10366_57;
                                                                                                                          end else begin
                                                                                                                            _T_18065_57 <= 8'h0;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_57 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_58) begin
        if (_T_16883) begin
          _T_18065_58 <= _T_10366_0;
        end else begin
          if (_T_16881) begin
            _T_18065_58 <= _T_10366_1;
          end else begin
            if (_T_16879) begin
              _T_18065_58 <= _T_10366_2;
            end else begin
              if (_T_16877) begin
                _T_18065_58 <= _T_10366_3;
              end else begin
                if (_T_16875) begin
                  _T_18065_58 <= _T_10366_4;
                end else begin
                  if (_T_16873) begin
                    _T_18065_58 <= _T_10366_5;
                  end else begin
                    if (_T_16871) begin
                      _T_18065_58 <= _T_10366_6;
                    end else begin
                      if (_T_16869) begin
                        _T_18065_58 <= _T_10366_7;
                      end else begin
                        if (_T_16867) begin
                          _T_18065_58 <= _T_10366_8;
                        end else begin
                          if (_T_16865) begin
                            _T_18065_58 <= _T_10366_9;
                          end else begin
                            if (_T_16863) begin
                              _T_18065_58 <= _T_10366_10;
                            end else begin
                              if (_T_16861) begin
                                _T_18065_58 <= _T_10366_11;
                              end else begin
                                if (_T_16859) begin
                                  _T_18065_58 <= _T_10366_12;
                                end else begin
                                  if (_T_16857) begin
                                    _T_18065_58 <= _T_10366_13;
                                  end else begin
                                    if (_T_16855) begin
                                      _T_18065_58 <= _T_10366_14;
                                    end else begin
                                      if (_T_16853) begin
                                        _T_18065_58 <= _T_10366_15;
                                      end else begin
                                        if (_T_16851) begin
                                          _T_18065_58 <= _T_10366_16;
                                        end else begin
                                          if (_T_16849) begin
                                            _T_18065_58 <= _T_10366_17;
                                          end else begin
                                            if (_T_16847) begin
                                              _T_18065_58 <= _T_10366_18;
                                            end else begin
                                              if (_T_16845) begin
                                                _T_18065_58 <= _T_10366_19;
                                              end else begin
                                                if (_T_16843) begin
                                                  _T_18065_58 <= _T_10366_20;
                                                end else begin
                                                  if (_T_16841) begin
                                                    _T_18065_58 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_16839) begin
                                                      _T_18065_58 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_16837) begin
                                                        _T_18065_58 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_16835) begin
                                                          _T_18065_58 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_16833) begin
                                                            _T_18065_58 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_16831) begin
                                                              _T_18065_58 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_16829) begin
                                                                _T_18065_58 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_16827) begin
                                                                  _T_18065_58 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_16825) begin
                                                                    _T_18065_58 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_16823) begin
                                                                      _T_18065_58 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_16821) begin
                                                                        _T_18065_58 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_16819) begin
                                                                          _T_18065_58 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_16817) begin
                                                                            _T_18065_58 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_16815) begin
                                                                              _T_18065_58 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_16813) begin
                                                                                _T_18065_58 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_16811) begin
                                                                                  _T_18065_58 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_16809) begin
                                                                                    _T_18065_58 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_16807) begin
                                                                                      _T_18065_58 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_16805) begin
                                                                                        _T_18065_58 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_16803) begin
                                                                                          _T_18065_58 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_16801) begin
                                                                                            _T_18065_58 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_16799) begin
                                                                                              _T_18065_58 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_16797) begin
                                                                                                _T_18065_58 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_16795) begin
                                                                                                  _T_18065_58 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_16793) begin
                                                                                                    _T_18065_58 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_16791) begin
                                                                                                      _T_18065_58 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_16789) begin
                                                                                                        _T_18065_58 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_16787) begin
                                                                                                          _T_18065_58 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_16785) begin
                                                                                                            _T_18065_58 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_16783) begin
                                                                                                              _T_18065_58 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_16781) begin
                                                                                                                _T_18065_58 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_16779) begin
                                                                                                                  _T_18065_58 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_16777) begin
                                                                                                                    _T_18065_58 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_16775) begin
                                                                                                                      _T_18065_58 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_16773) begin
                                                                                                                        _T_18065_58 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_16771) begin
                                                                                                                          _T_18065_58 <= _T_10366_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_16769) begin
                                                                                                                            _T_18065_58 <= _T_10366_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_16767) begin
                                                                                                                              _T_18065_58 <= _T_10366_58;
                                                                                                                            end else begin
                                                                                                                              _T_18065_58 <= 8'h0;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_58 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_59) begin
        if (_T_17064) begin
          _T_18065_59 <= _T_10366_0;
        end else begin
          if (_T_17062) begin
            _T_18065_59 <= _T_10366_1;
          end else begin
            if (_T_17060) begin
              _T_18065_59 <= _T_10366_2;
            end else begin
              if (_T_17058) begin
                _T_18065_59 <= _T_10366_3;
              end else begin
                if (_T_17056) begin
                  _T_18065_59 <= _T_10366_4;
                end else begin
                  if (_T_17054) begin
                    _T_18065_59 <= _T_10366_5;
                  end else begin
                    if (_T_17052) begin
                      _T_18065_59 <= _T_10366_6;
                    end else begin
                      if (_T_17050) begin
                        _T_18065_59 <= _T_10366_7;
                      end else begin
                        if (_T_17048) begin
                          _T_18065_59 <= _T_10366_8;
                        end else begin
                          if (_T_17046) begin
                            _T_18065_59 <= _T_10366_9;
                          end else begin
                            if (_T_17044) begin
                              _T_18065_59 <= _T_10366_10;
                            end else begin
                              if (_T_17042) begin
                                _T_18065_59 <= _T_10366_11;
                              end else begin
                                if (_T_17040) begin
                                  _T_18065_59 <= _T_10366_12;
                                end else begin
                                  if (_T_17038) begin
                                    _T_18065_59 <= _T_10366_13;
                                  end else begin
                                    if (_T_17036) begin
                                      _T_18065_59 <= _T_10366_14;
                                    end else begin
                                      if (_T_17034) begin
                                        _T_18065_59 <= _T_10366_15;
                                      end else begin
                                        if (_T_17032) begin
                                          _T_18065_59 <= _T_10366_16;
                                        end else begin
                                          if (_T_17030) begin
                                            _T_18065_59 <= _T_10366_17;
                                          end else begin
                                            if (_T_17028) begin
                                              _T_18065_59 <= _T_10366_18;
                                            end else begin
                                              if (_T_17026) begin
                                                _T_18065_59 <= _T_10366_19;
                                              end else begin
                                                if (_T_17024) begin
                                                  _T_18065_59 <= _T_10366_20;
                                                end else begin
                                                  if (_T_17022) begin
                                                    _T_18065_59 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_17020) begin
                                                      _T_18065_59 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_17018) begin
                                                        _T_18065_59 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_17016) begin
                                                          _T_18065_59 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_17014) begin
                                                            _T_18065_59 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_17012) begin
                                                              _T_18065_59 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_17010) begin
                                                                _T_18065_59 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_17008) begin
                                                                  _T_18065_59 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_17006) begin
                                                                    _T_18065_59 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_17004) begin
                                                                      _T_18065_59 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_17002) begin
                                                                        _T_18065_59 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_17000) begin
                                                                          _T_18065_59 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_16998) begin
                                                                            _T_18065_59 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_16996) begin
                                                                              _T_18065_59 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_16994) begin
                                                                                _T_18065_59 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_16992) begin
                                                                                  _T_18065_59 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_16990) begin
                                                                                    _T_18065_59 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_16988) begin
                                                                                      _T_18065_59 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_16986) begin
                                                                                        _T_18065_59 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_16984) begin
                                                                                          _T_18065_59 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_16982) begin
                                                                                            _T_18065_59 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_16980) begin
                                                                                              _T_18065_59 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_16978) begin
                                                                                                _T_18065_59 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_16976) begin
                                                                                                  _T_18065_59 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_16974) begin
                                                                                                    _T_18065_59 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_16972) begin
                                                                                                      _T_18065_59 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_16970) begin
                                                                                                        _T_18065_59 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_16968) begin
                                                                                                          _T_18065_59 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_16966) begin
                                                                                                            _T_18065_59 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_16964) begin
                                                                                                              _T_18065_59 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_16962) begin
                                                                                                                _T_18065_59 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_16960) begin
                                                                                                                  _T_18065_59 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_16958) begin
                                                                                                                    _T_18065_59 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_16956) begin
                                                                                                                      _T_18065_59 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_16954) begin
                                                                                                                        _T_18065_59 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_16952) begin
                                                                                                                          _T_18065_59 <= _T_10366_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_16950) begin
                                                                                                                            _T_18065_59 <= _T_10366_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_16948) begin
                                                                                                                              _T_18065_59 <= _T_10366_58;
                                                                                                                            end else begin
                                                                                                                              if (_T_16946) begin
                                                                                                                                _T_18065_59 <= _T_10366_59;
                                                                                                                              end else begin
                                                                                                                                _T_18065_59 <= 8'h0;
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_59 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_60) begin
        if (_T_17248) begin
          _T_18065_60 <= _T_10366_0;
        end else begin
          if (_T_17246) begin
            _T_18065_60 <= _T_10366_1;
          end else begin
            if (_T_17244) begin
              _T_18065_60 <= _T_10366_2;
            end else begin
              if (_T_17242) begin
                _T_18065_60 <= _T_10366_3;
              end else begin
                if (_T_17240) begin
                  _T_18065_60 <= _T_10366_4;
                end else begin
                  if (_T_17238) begin
                    _T_18065_60 <= _T_10366_5;
                  end else begin
                    if (_T_17236) begin
                      _T_18065_60 <= _T_10366_6;
                    end else begin
                      if (_T_17234) begin
                        _T_18065_60 <= _T_10366_7;
                      end else begin
                        if (_T_17232) begin
                          _T_18065_60 <= _T_10366_8;
                        end else begin
                          if (_T_17230) begin
                            _T_18065_60 <= _T_10366_9;
                          end else begin
                            if (_T_17228) begin
                              _T_18065_60 <= _T_10366_10;
                            end else begin
                              if (_T_17226) begin
                                _T_18065_60 <= _T_10366_11;
                              end else begin
                                if (_T_17224) begin
                                  _T_18065_60 <= _T_10366_12;
                                end else begin
                                  if (_T_17222) begin
                                    _T_18065_60 <= _T_10366_13;
                                  end else begin
                                    if (_T_17220) begin
                                      _T_18065_60 <= _T_10366_14;
                                    end else begin
                                      if (_T_17218) begin
                                        _T_18065_60 <= _T_10366_15;
                                      end else begin
                                        if (_T_17216) begin
                                          _T_18065_60 <= _T_10366_16;
                                        end else begin
                                          if (_T_17214) begin
                                            _T_18065_60 <= _T_10366_17;
                                          end else begin
                                            if (_T_17212) begin
                                              _T_18065_60 <= _T_10366_18;
                                            end else begin
                                              if (_T_17210) begin
                                                _T_18065_60 <= _T_10366_19;
                                              end else begin
                                                if (_T_17208) begin
                                                  _T_18065_60 <= _T_10366_20;
                                                end else begin
                                                  if (_T_17206) begin
                                                    _T_18065_60 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_17204) begin
                                                      _T_18065_60 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_17202) begin
                                                        _T_18065_60 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_17200) begin
                                                          _T_18065_60 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_17198) begin
                                                            _T_18065_60 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_17196) begin
                                                              _T_18065_60 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_17194) begin
                                                                _T_18065_60 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_17192) begin
                                                                  _T_18065_60 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_17190) begin
                                                                    _T_18065_60 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_17188) begin
                                                                      _T_18065_60 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_17186) begin
                                                                        _T_18065_60 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_17184) begin
                                                                          _T_18065_60 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_17182) begin
                                                                            _T_18065_60 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_17180) begin
                                                                              _T_18065_60 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_17178) begin
                                                                                _T_18065_60 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_17176) begin
                                                                                  _T_18065_60 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_17174) begin
                                                                                    _T_18065_60 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_17172) begin
                                                                                      _T_18065_60 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_17170) begin
                                                                                        _T_18065_60 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_17168) begin
                                                                                          _T_18065_60 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_17166) begin
                                                                                            _T_18065_60 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_17164) begin
                                                                                              _T_18065_60 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_17162) begin
                                                                                                _T_18065_60 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_17160) begin
                                                                                                  _T_18065_60 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_17158) begin
                                                                                                    _T_18065_60 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_17156) begin
                                                                                                      _T_18065_60 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_17154) begin
                                                                                                        _T_18065_60 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_17152) begin
                                                                                                          _T_18065_60 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_17150) begin
                                                                                                            _T_18065_60 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_17148) begin
                                                                                                              _T_18065_60 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_17146) begin
                                                                                                                _T_18065_60 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_17144) begin
                                                                                                                  _T_18065_60 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_17142) begin
                                                                                                                    _T_18065_60 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_17140) begin
                                                                                                                      _T_18065_60 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_17138) begin
                                                                                                                        _T_18065_60 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_17136) begin
                                                                                                                          _T_18065_60 <= _T_10366_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_17134) begin
                                                                                                                            _T_18065_60 <= _T_10366_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_17132) begin
                                                                                                                              _T_18065_60 <= _T_10366_58;
                                                                                                                            end else begin
                                                                                                                              if (_T_17130) begin
                                                                                                                                _T_18065_60 <= _T_10366_59;
                                                                                                                              end else begin
                                                                                                                                if (_T_17128) begin
                                                                                                                                  _T_18065_60 <= _T_10366_60;
                                                                                                                                end else begin
                                                                                                                                  _T_18065_60 <= 8'h0;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_60 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_61) begin
        if (_T_17435) begin
          _T_18065_61 <= _T_10366_0;
        end else begin
          if (_T_17433) begin
            _T_18065_61 <= _T_10366_1;
          end else begin
            if (_T_17431) begin
              _T_18065_61 <= _T_10366_2;
            end else begin
              if (_T_17429) begin
                _T_18065_61 <= _T_10366_3;
              end else begin
                if (_T_17427) begin
                  _T_18065_61 <= _T_10366_4;
                end else begin
                  if (_T_17425) begin
                    _T_18065_61 <= _T_10366_5;
                  end else begin
                    if (_T_17423) begin
                      _T_18065_61 <= _T_10366_6;
                    end else begin
                      if (_T_17421) begin
                        _T_18065_61 <= _T_10366_7;
                      end else begin
                        if (_T_17419) begin
                          _T_18065_61 <= _T_10366_8;
                        end else begin
                          if (_T_17417) begin
                            _T_18065_61 <= _T_10366_9;
                          end else begin
                            if (_T_17415) begin
                              _T_18065_61 <= _T_10366_10;
                            end else begin
                              if (_T_17413) begin
                                _T_18065_61 <= _T_10366_11;
                              end else begin
                                if (_T_17411) begin
                                  _T_18065_61 <= _T_10366_12;
                                end else begin
                                  if (_T_17409) begin
                                    _T_18065_61 <= _T_10366_13;
                                  end else begin
                                    if (_T_17407) begin
                                      _T_18065_61 <= _T_10366_14;
                                    end else begin
                                      if (_T_17405) begin
                                        _T_18065_61 <= _T_10366_15;
                                      end else begin
                                        if (_T_17403) begin
                                          _T_18065_61 <= _T_10366_16;
                                        end else begin
                                          if (_T_17401) begin
                                            _T_18065_61 <= _T_10366_17;
                                          end else begin
                                            if (_T_17399) begin
                                              _T_18065_61 <= _T_10366_18;
                                            end else begin
                                              if (_T_17397) begin
                                                _T_18065_61 <= _T_10366_19;
                                              end else begin
                                                if (_T_17395) begin
                                                  _T_18065_61 <= _T_10366_20;
                                                end else begin
                                                  if (_T_17393) begin
                                                    _T_18065_61 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_17391) begin
                                                      _T_18065_61 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_17389) begin
                                                        _T_18065_61 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_17387) begin
                                                          _T_18065_61 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_17385) begin
                                                            _T_18065_61 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_17383) begin
                                                              _T_18065_61 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_17381) begin
                                                                _T_18065_61 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_17379) begin
                                                                  _T_18065_61 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_17377) begin
                                                                    _T_18065_61 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_17375) begin
                                                                      _T_18065_61 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_17373) begin
                                                                        _T_18065_61 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_17371) begin
                                                                          _T_18065_61 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_17369) begin
                                                                            _T_18065_61 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_17367) begin
                                                                              _T_18065_61 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_17365) begin
                                                                                _T_18065_61 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_17363) begin
                                                                                  _T_18065_61 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_17361) begin
                                                                                    _T_18065_61 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_17359) begin
                                                                                      _T_18065_61 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_17357) begin
                                                                                        _T_18065_61 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_17355) begin
                                                                                          _T_18065_61 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_17353) begin
                                                                                            _T_18065_61 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_17351) begin
                                                                                              _T_18065_61 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_17349) begin
                                                                                                _T_18065_61 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_17347) begin
                                                                                                  _T_18065_61 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_17345) begin
                                                                                                    _T_18065_61 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_17343) begin
                                                                                                      _T_18065_61 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_17341) begin
                                                                                                        _T_18065_61 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_17339) begin
                                                                                                          _T_18065_61 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_17337) begin
                                                                                                            _T_18065_61 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_17335) begin
                                                                                                              _T_18065_61 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_17333) begin
                                                                                                                _T_18065_61 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_17331) begin
                                                                                                                  _T_18065_61 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_17329) begin
                                                                                                                    _T_18065_61 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_17327) begin
                                                                                                                      _T_18065_61 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_17325) begin
                                                                                                                        _T_18065_61 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_17323) begin
                                                                                                                          _T_18065_61 <= _T_10366_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_17321) begin
                                                                                                                            _T_18065_61 <= _T_10366_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_17319) begin
                                                                                                                              _T_18065_61 <= _T_10366_58;
                                                                                                                            end else begin
                                                                                                                              if (_T_17317) begin
                                                                                                                                _T_18065_61 <= _T_10366_59;
                                                                                                                              end else begin
                                                                                                                                if (_T_17315) begin
                                                                                                                                  _T_18065_61 <= _T_10366_60;
                                                                                                                                end else begin
                                                                                                                                  if (_T_17313) begin
                                                                                                                                    _T_18065_61 <= _T_10366_61;
                                                                                                                                  end else begin
                                                                                                                                    _T_18065_61 <= 8'h0;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_61 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_62) begin
        if (_T_17625) begin
          _T_18065_62 <= _T_10366_0;
        end else begin
          if (_T_17623) begin
            _T_18065_62 <= _T_10366_1;
          end else begin
            if (_T_17621) begin
              _T_18065_62 <= _T_10366_2;
            end else begin
              if (_T_17619) begin
                _T_18065_62 <= _T_10366_3;
              end else begin
                if (_T_17617) begin
                  _T_18065_62 <= _T_10366_4;
                end else begin
                  if (_T_17615) begin
                    _T_18065_62 <= _T_10366_5;
                  end else begin
                    if (_T_17613) begin
                      _T_18065_62 <= _T_10366_6;
                    end else begin
                      if (_T_17611) begin
                        _T_18065_62 <= _T_10366_7;
                      end else begin
                        if (_T_17609) begin
                          _T_18065_62 <= _T_10366_8;
                        end else begin
                          if (_T_17607) begin
                            _T_18065_62 <= _T_10366_9;
                          end else begin
                            if (_T_17605) begin
                              _T_18065_62 <= _T_10366_10;
                            end else begin
                              if (_T_17603) begin
                                _T_18065_62 <= _T_10366_11;
                              end else begin
                                if (_T_17601) begin
                                  _T_18065_62 <= _T_10366_12;
                                end else begin
                                  if (_T_17599) begin
                                    _T_18065_62 <= _T_10366_13;
                                  end else begin
                                    if (_T_17597) begin
                                      _T_18065_62 <= _T_10366_14;
                                    end else begin
                                      if (_T_17595) begin
                                        _T_18065_62 <= _T_10366_15;
                                      end else begin
                                        if (_T_17593) begin
                                          _T_18065_62 <= _T_10366_16;
                                        end else begin
                                          if (_T_17591) begin
                                            _T_18065_62 <= _T_10366_17;
                                          end else begin
                                            if (_T_17589) begin
                                              _T_18065_62 <= _T_10366_18;
                                            end else begin
                                              if (_T_17587) begin
                                                _T_18065_62 <= _T_10366_19;
                                              end else begin
                                                if (_T_17585) begin
                                                  _T_18065_62 <= _T_10366_20;
                                                end else begin
                                                  if (_T_17583) begin
                                                    _T_18065_62 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_17581) begin
                                                      _T_18065_62 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_17579) begin
                                                        _T_18065_62 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_17577) begin
                                                          _T_18065_62 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_17575) begin
                                                            _T_18065_62 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_17573) begin
                                                              _T_18065_62 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_17571) begin
                                                                _T_18065_62 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_17569) begin
                                                                  _T_18065_62 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_17567) begin
                                                                    _T_18065_62 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_17565) begin
                                                                      _T_18065_62 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_17563) begin
                                                                        _T_18065_62 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_17561) begin
                                                                          _T_18065_62 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_17559) begin
                                                                            _T_18065_62 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_17557) begin
                                                                              _T_18065_62 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_17555) begin
                                                                                _T_18065_62 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_17553) begin
                                                                                  _T_18065_62 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_17551) begin
                                                                                    _T_18065_62 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_17549) begin
                                                                                      _T_18065_62 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_17547) begin
                                                                                        _T_18065_62 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_17545) begin
                                                                                          _T_18065_62 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_17543) begin
                                                                                            _T_18065_62 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_17541) begin
                                                                                              _T_18065_62 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_17539) begin
                                                                                                _T_18065_62 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_17537) begin
                                                                                                  _T_18065_62 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_17535) begin
                                                                                                    _T_18065_62 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_17533) begin
                                                                                                      _T_18065_62 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_17531) begin
                                                                                                        _T_18065_62 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_17529) begin
                                                                                                          _T_18065_62 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_17527) begin
                                                                                                            _T_18065_62 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_17525) begin
                                                                                                              _T_18065_62 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_17523) begin
                                                                                                                _T_18065_62 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_17521) begin
                                                                                                                  _T_18065_62 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_17519) begin
                                                                                                                    _T_18065_62 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_17517) begin
                                                                                                                      _T_18065_62 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_17515) begin
                                                                                                                        _T_18065_62 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_17513) begin
                                                                                                                          _T_18065_62 <= _T_10366_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_17511) begin
                                                                                                                            _T_18065_62 <= _T_10366_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_17509) begin
                                                                                                                              _T_18065_62 <= _T_10366_58;
                                                                                                                            end else begin
                                                                                                                              if (_T_17507) begin
                                                                                                                                _T_18065_62 <= _T_10366_59;
                                                                                                                              end else begin
                                                                                                                                if (_T_17505) begin
                                                                                                                                  _T_18065_62 <= _T_10366_60;
                                                                                                                                end else begin
                                                                                                                                  if (_T_17503) begin
                                                                                                                                    _T_18065_62 <= _T_10366_61;
                                                                                                                                  end else begin
                                                                                                                                    if (_T_17501) begin
                                                                                                                                      _T_18065_62 <= _T_10366_62;
                                                                                                                                    end else begin
                                                                                                                                      _T_18065_62 <= 8'h0;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_62 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_63) begin
        if (_T_17818) begin
          _T_18065_63 <= _T_10366_0;
        end else begin
          if (_T_17816) begin
            _T_18065_63 <= _T_10366_1;
          end else begin
            if (_T_17814) begin
              _T_18065_63 <= _T_10366_2;
            end else begin
              if (_T_17812) begin
                _T_18065_63 <= _T_10366_3;
              end else begin
                if (_T_17810) begin
                  _T_18065_63 <= _T_10366_4;
                end else begin
                  if (_T_17808) begin
                    _T_18065_63 <= _T_10366_5;
                  end else begin
                    if (_T_17806) begin
                      _T_18065_63 <= _T_10366_6;
                    end else begin
                      if (_T_17804) begin
                        _T_18065_63 <= _T_10366_7;
                      end else begin
                        if (_T_17802) begin
                          _T_18065_63 <= _T_10366_8;
                        end else begin
                          if (_T_17800) begin
                            _T_18065_63 <= _T_10366_9;
                          end else begin
                            if (_T_17798) begin
                              _T_18065_63 <= _T_10366_10;
                            end else begin
                              if (_T_17796) begin
                                _T_18065_63 <= _T_10366_11;
                              end else begin
                                if (_T_17794) begin
                                  _T_18065_63 <= _T_10366_12;
                                end else begin
                                  if (_T_17792) begin
                                    _T_18065_63 <= _T_10366_13;
                                  end else begin
                                    if (_T_17790) begin
                                      _T_18065_63 <= _T_10366_14;
                                    end else begin
                                      if (_T_17788) begin
                                        _T_18065_63 <= _T_10366_15;
                                      end else begin
                                        if (_T_17786) begin
                                          _T_18065_63 <= _T_10366_16;
                                        end else begin
                                          if (_T_17784) begin
                                            _T_18065_63 <= _T_10366_17;
                                          end else begin
                                            if (_T_17782) begin
                                              _T_18065_63 <= _T_10366_18;
                                            end else begin
                                              if (_T_17780) begin
                                                _T_18065_63 <= _T_10366_19;
                                              end else begin
                                                if (_T_17778) begin
                                                  _T_18065_63 <= _T_10366_20;
                                                end else begin
                                                  if (_T_17776) begin
                                                    _T_18065_63 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_17774) begin
                                                      _T_18065_63 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_17772) begin
                                                        _T_18065_63 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_17770) begin
                                                          _T_18065_63 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_17768) begin
                                                            _T_18065_63 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_17766) begin
                                                              _T_18065_63 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_17764) begin
                                                                _T_18065_63 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_17762) begin
                                                                  _T_18065_63 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_17760) begin
                                                                    _T_18065_63 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_17758) begin
                                                                      _T_18065_63 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_17756) begin
                                                                        _T_18065_63 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_17754) begin
                                                                          _T_18065_63 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_17752) begin
                                                                            _T_18065_63 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_17750) begin
                                                                              _T_18065_63 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_17748) begin
                                                                                _T_18065_63 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_17746) begin
                                                                                  _T_18065_63 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_17744) begin
                                                                                    _T_18065_63 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_17742) begin
                                                                                      _T_18065_63 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_17740) begin
                                                                                        _T_18065_63 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_17738) begin
                                                                                          _T_18065_63 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_17736) begin
                                                                                            _T_18065_63 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_17734) begin
                                                                                              _T_18065_63 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_17732) begin
                                                                                                _T_18065_63 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_17730) begin
                                                                                                  _T_18065_63 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_17728) begin
                                                                                                    _T_18065_63 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_17726) begin
                                                                                                      _T_18065_63 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_17724) begin
                                                                                                        _T_18065_63 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_17722) begin
                                                                                                          _T_18065_63 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_17720) begin
                                                                                                            _T_18065_63 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_17718) begin
                                                                                                              _T_18065_63 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_17716) begin
                                                                                                                _T_18065_63 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_17714) begin
                                                                                                                  _T_18065_63 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_17712) begin
                                                                                                                    _T_18065_63 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_17710) begin
                                                                                                                      _T_18065_63 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_17708) begin
                                                                                                                        _T_18065_63 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_17706) begin
                                                                                                                          _T_18065_63 <= _T_10366_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_17704) begin
                                                                                                                            _T_18065_63 <= _T_10366_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_17702) begin
                                                                                                                              _T_18065_63 <= _T_10366_58;
                                                                                                                            end else begin
                                                                                                                              if (_T_17700) begin
                                                                                                                                _T_18065_63 <= _T_10366_59;
                                                                                                                              end else begin
                                                                                                                                if (_T_17698) begin
                                                                                                                                  _T_18065_63 <= _T_10366_60;
                                                                                                                                end else begin
                                                                                                                                  if (_T_17696) begin
                                                                                                                                    _T_18065_63 <= _T_10366_61;
                                                                                                                                  end else begin
                                                                                                                                    if (_T_17694) begin
                                                                                                                                      _T_18065_63 <= _T_10366_62;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_17692) begin
                                                                                                                                        _T_18065_63 <= _T_10366_63;
                                                                                                                                      end else begin
                                                                                                                                        _T_18065_63 <= 8'h0;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_63 <= 8'h0;
      end
    end
    if (reset) begin
      _T_18396 <= 1'h0;
    end else begin
      _T_18396 <= _T_17822;
    end
    if (_T_17822) begin
      _T_18400_0 <= _T_18267;
    end
    if (_T_17822) begin
      _T_18400_1 <= _T_18269;
    end
    if (_T_17822) begin
      _T_18400_2 <= _T_18271;
    end
    if (_T_17822) begin
      _T_18400_3 <= _T_18273;
    end
    if (_T_17822) begin
      _T_18400_4 <= _T_18275;
    end
    if (_T_17822) begin
      _T_18400_5 <= _T_18277;
    end
    if (_T_17822) begin
      _T_18400_6 <= _T_18279;
    end
    if (_T_17822) begin
      _T_18400_7 <= _T_18281;
    end
    if (_T_17822) begin
      _T_18400_8 <= _T_18283;
    end
    if (_T_17822) begin
      _T_18400_9 <= _T_18285;
    end
    if (_T_17822) begin
      _T_18400_10 <= _T_18287;
    end
    if (_T_17822) begin
      _T_18400_11 <= _T_18289;
    end
    if (_T_17822) begin
      _T_18400_12 <= _T_18291;
    end
    if (_T_17822) begin
      _T_18400_13 <= _T_18293;
    end
    if (_T_17822) begin
      _T_18400_14 <= _T_18295;
    end
    if (_T_17822) begin
      _T_18400_15 <= _T_18297;
    end
    if (_T_17822) begin
      _T_18400_16 <= _T_18299;
    end
    if (_T_17822) begin
      _T_18400_17 <= _T_18301;
    end
    if (_T_17822) begin
      _T_18400_18 <= _T_18303;
    end
    if (_T_17822) begin
      _T_18400_19 <= _T_18305;
    end
    if (_T_17822) begin
      _T_18400_20 <= _T_18307;
    end
    if (_T_17822) begin
      _T_18400_21 <= _T_18309;
    end
    if (_T_17822) begin
      _T_18400_22 <= _T_18311;
    end
    if (_T_17822) begin
      _T_18400_23 <= _T_18313;
    end
    if (_T_17822) begin
      _T_18400_24 <= _T_18315;
    end
    if (_T_17822) begin
      _T_18400_25 <= _T_18317;
    end
    if (_T_17822) begin
      _T_18400_26 <= _T_18319;
    end
    if (_T_17822) begin
      _T_18400_27 <= _T_18321;
    end
    if (_T_17822) begin
      _T_18400_28 <= _T_18323;
    end
    if (_T_17822) begin
      _T_18400_29 <= _T_18325;
    end
    if (_T_17822) begin
      _T_18400_30 <= _T_18327;
    end
    if (_T_17822) begin
      _T_18400_31 <= _T_18329;
    end
    if (_T_17822) begin
      _T_18400_32 <= _T_18331;
    end
    if (_T_17822) begin
      _T_18400_33 <= _T_18333;
    end
    if (_T_17822) begin
      _T_18400_34 <= _T_18335;
    end
    if (_T_17822) begin
      _T_18400_35 <= _T_18337;
    end
    if (_T_17822) begin
      _T_18400_36 <= _T_18339;
    end
    if (_T_17822) begin
      _T_18400_37 <= _T_18341;
    end
    if (_T_17822) begin
      _T_18400_38 <= _T_18343;
    end
    if (_T_17822) begin
      _T_18400_39 <= _T_18345;
    end
    if (_T_17822) begin
      _T_18400_40 <= _T_18347;
    end
    if (_T_17822) begin
      _T_18400_41 <= _T_18349;
    end
    if (_T_17822) begin
      _T_18400_42 <= _T_18351;
    end
    if (_T_17822) begin
      _T_18400_43 <= _T_18353;
    end
    if (_T_17822) begin
      _T_18400_44 <= _T_18355;
    end
    if (_T_17822) begin
      _T_18400_45 <= _T_18357;
    end
    if (_T_17822) begin
      _T_18400_46 <= _T_18359;
    end
    if (_T_17822) begin
      _T_18400_47 <= _T_18361;
    end
    if (_T_17822) begin
      _T_18400_48 <= _T_18363;
    end
    if (_T_17822) begin
      _T_18400_49 <= _T_18365;
    end
    if (_T_17822) begin
      _T_18400_50 <= _T_18367;
    end
    if (_T_17822) begin
      _T_18400_51 <= _T_18369;
    end
    if (_T_17822) begin
      _T_18400_52 <= _T_18371;
    end
    if (_T_17822) begin
      _T_18400_53 <= _T_18373;
    end
    if (_T_17822) begin
      _T_18400_54 <= _T_18375;
    end
    if (_T_17822) begin
      _T_18400_55 <= _T_18377;
    end
    if (_T_17822) begin
      _T_18400_56 <= _T_18379;
    end
    if (_T_17822) begin
      _T_18400_57 <= _T_18381;
    end
    if (_T_17822) begin
      _T_18400_58 <= _T_18383;
    end
    if (_T_17822) begin
      _T_18400_59 <= _T_18385;
    end
    if (_T_17822) begin
      _T_18400_60 <= _T_18387;
    end
    if (_T_17822) begin
      _T_18400_61 <= _T_18389;
    end
    if (_T_17822) begin
      _T_18400_62 <= _T_18391;
    end
    if (_T_17822) begin
      _T_18400_63 <= _T_18393;
    end
    if (reset) begin
      _T_18605_0 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_0 <= _T_17961_0;
      end
    end
    if (reset) begin
      _T_18605_1 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_1 <= _T_17961_1;
      end
    end
    if (reset) begin
      _T_18605_2 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_2 <= _T_17961_2;
      end
    end
    if (reset) begin
      _T_18605_3 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_3 <= _T_17961_3;
      end
    end
    if (reset) begin
      _T_18605_4 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_4 <= _T_17961_4;
      end
    end
    if (reset) begin
      _T_18605_5 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_5 <= _T_17961_5;
      end
    end
    if (reset) begin
      _T_18605_6 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_6 <= _T_17961_6;
      end
    end
    if (reset) begin
      _T_18605_7 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_7 <= _T_17961_7;
      end
    end
    if (reset) begin
      _T_18605_8 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_8 <= _T_17961_8;
      end
    end
    if (reset) begin
      _T_18605_9 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_9 <= _T_17961_9;
      end
    end
    if (reset) begin
      _T_18605_10 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_10 <= _T_17961_10;
      end
    end
    if (reset) begin
      _T_18605_11 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_11 <= _T_17961_11;
      end
    end
    if (reset) begin
      _T_18605_12 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_12 <= _T_17961_12;
      end
    end
    if (reset) begin
      _T_18605_13 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_13 <= _T_17961_13;
      end
    end
    if (reset) begin
      _T_18605_14 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_14 <= _T_17961_14;
      end
    end
    if (reset) begin
      _T_18605_15 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_15 <= _T_17961_15;
      end
    end
    if (reset) begin
      _T_18605_16 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_16 <= _T_17961_16;
      end
    end
    if (reset) begin
      _T_18605_17 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_17 <= _T_17961_17;
      end
    end
    if (reset) begin
      _T_18605_18 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_18 <= _T_17961_18;
      end
    end
    if (reset) begin
      _T_18605_19 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_19 <= _T_17961_19;
      end
    end
    if (reset) begin
      _T_18605_20 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_20 <= _T_17961_20;
      end
    end
    if (reset) begin
      _T_18605_21 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_21 <= _T_17961_21;
      end
    end
    if (reset) begin
      _T_18605_22 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_22 <= _T_17961_22;
      end
    end
    if (reset) begin
      _T_18605_23 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_23 <= _T_17961_23;
      end
    end
    if (reset) begin
      _T_18605_24 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_24 <= _T_17961_24;
      end
    end
    if (reset) begin
      _T_18605_25 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_25 <= _T_17961_25;
      end
    end
    if (reset) begin
      _T_18605_26 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_26 <= _T_17961_26;
      end
    end
    if (reset) begin
      _T_18605_27 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_27 <= _T_17961_27;
      end
    end
    if (reset) begin
      _T_18605_28 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_28 <= _T_17961_28;
      end
    end
    if (reset) begin
      _T_18605_29 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_29 <= _T_17961_29;
      end
    end
    if (reset) begin
      _T_18605_30 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_30 <= _T_17961_30;
      end
    end
    if (reset) begin
      _T_18605_31 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_31 <= _T_17961_31;
      end
    end
    if (_T_17822) begin
      _T_18709_0 <= _T_18065_0;
    end
    if (_T_17822) begin
      _T_18709_1 <= _T_18065_1;
    end
    if (_T_17822) begin
      _T_18709_2 <= _T_18065_2;
    end
    if (_T_17822) begin
      _T_18709_3 <= _T_18065_3;
    end
    if (_T_17822) begin
      _T_18709_4 <= _T_18065_4;
    end
    if (_T_17822) begin
      _T_18709_5 <= _T_18065_5;
    end
    if (_T_17822) begin
      _T_18709_6 <= _T_18065_6;
    end
    if (_T_17822) begin
      _T_18709_7 <= _T_18065_7;
    end
    if (_T_17822) begin
      _T_18709_8 <= _T_18065_8;
    end
    if (_T_17822) begin
      _T_18709_9 <= _T_18065_9;
    end
    if (_T_17822) begin
      _T_18709_10 <= _T_18065_10;
    end
    if (_T_17822) begin
      _T_18709_11 <= _T_18065_11;
    end
    if (_T_17822) begin
      _T_18709_12 <= _T_18065_12;
    end
    if (_T_17822) begin
      _T_18709_13 <= _T_18065_13;
    end
    if (_T_17822) begin
      _T_18709_14 <= _T_18065_14;
    end
    if (_T_17822) begin
      _T_18709_15 <= _T_18065_15;
    end
    if (_T_17822) begin
      _T_18709_16 <= _T_18065_16;
    end
    if (_T_17822) begin
      _T_18709_17 <= _T_18065_17;
    end
    if (_T_17822) begin
      _T_18709_18 <= _T_18065_18;
    end
    if (_T_17822) begin
      _T_18709_19 <= _T_18065_19;
    end
    if (_T_17822) begin
      _T_18709_20 <= _T_18065_20;
    end
    if (_T_17822) begin
      _T_18709_21 <= _T_18065_21;
    end
    if (_T_17822) begin
      _T_18709_22 <= _T_18065_22;
    end
    if (_T_17822) begin
      _T_18709_23 <= _T_18065_23;
    end
    if (_T_17822) begin
      _T_18709_24 <= _T_18065_24;
    end
    if (_T_17822) begin
      _T_18709_25 <= _T_18065_25;
    end
    if (_T_17822) begin
      _T_18709_26 <= _T_18065_26;
    end
    if (_T_17822) begin
      _T_18709_27 <= _T_18065_27;
    end
    if (_T_17822) begin
      _T_18709_28 <= _T_18065_28;
    end
    if (_T_17822) begin
      _T_18709_29 <= _T_18065_29;
    end
    if (_T_17822) begin
      _T_18709_30 <= _T_18065_30;
    end
    if (_T_17822) begin
      _T_18709_31 <= _T_18065_31;
    end
    if (_T_17822) begin
      _T_18709_32 <= _T_18065_32;
    end
    if (_T_17822) begin
      _T_18709_33 <= _T_18065_33;
    end
    if (_T_17822) begin
      _T_18709_34 <= _T_18065_34;
    end
    if (_T_17822) begin
      _T_18709_35 <= _T_18065_35;
    end
    if (_T_17822) begin
      _T_18709_36 <= _T_18065_36;
    end
    if (_T_17822) begin
      _T_18709_37 <= _T_18065_37;
    end
    if (_T_17822) begin
      _T_18709_38 <= _T_18065_38;
    end
    if (_T_17822) begin
      _T_18709_39 <= _T_18065_39;
    end
    if (_T_17822) begin
      _T_18709_40 <= _T_18065_40;
    end
    if (_T_17822) begin
      _T_18709_41 <= _T_18065_41;
    end
    if (_T_17822) begin
      _T_18709_42 <= _T_18065_42;
    end
    if (_T_17822) begin
      _T_18709_43 <= _T_18065_43;
    end
    if (_T_17822) begin
      _T_18709_44 <= _T_18065_44;
    end
    if (_T_17822) begin
      _T_18709_45 <= _T_18065_45;
    end
    if (_T_17822) begin
      _T_18709_46 <= _T_18065_46;
    end
    if (_T_17822) begin
      _T_18709_47 <= _T_18065_47;
    end
    if (_T_17822) begin
      _T_18709_48 <= _T_18065_48;
    end
    if (_T_17822) begin
      _T_18709_49 <= _T_18065_49;
    end
    if (_T_17822) begin
      _T_18709_50 <= _T_18065_50;
    end
    if (_T_17822) begin
      _T_18709_51 <= _T_18065_51;
    end
    if (_T_17822) begin
      _T_18709_52 <= _T_18065_52;
    end
    if (_T_17822) begin
      _T_18709_53 <= _T_18065_53;
    end
    if (_T_17822) begin
      _T_18709_54 <= _T_18065_54;
    end
    if (_T_17822) begin
      _T_18709_55 <= _T_18065_55;
    end
    if (_T_17822) begin
      _T_18709_56 <= _T_18065_56;
    end
    if (_T_17822) begin
      _T_18709_57 <= _T_18065_57;
    end
    if (_T_17822) begin
      _T_18709_58 <= _T_18065_58;
    end
    if (_T_17822) begin
      _T_18709_59 <= _T_18065_59;
    end
    if (_T_17822) begin
      _T_18709_60 <= _T_18065_60;
    end
    if (_T_17822) begin
      _T_18709_61 <= _T_18065_61;
    end
    if (_T_17822) begin
      _T_18709_62 <= _T_18065_62;
    end
    if (_T_17822) begin
      _T_18709_63 <= _T_18065_63;
    end
  end
endmodule
module NV_NVDLA_CSC_wl( // @[:@16367.2]
  input          reset, // @[:@16369.4]
  input          io_nvdla_core_clk, // @[:@16370.4]
  input          io_nvdla_core_ng_clk, // @[:@16370.4]
  input          io_sg2wl_pd_valid, // @[:@16370.4]
  input  [17:0]  io_sg2wl_pd_bits, // @[:@16370.4]
  input          io_sg2wl_reuse_rls, // @[:@16370.4]
  input  [1:0]   io_sc_state, // @[:@16370.4]
  input          io_sc2cdma_wt_pending_req, // @[:@16370.4]
  output         io_sc2cdma_wt_updt_valid, // @[:@16370.4]
  output [14:0]  io_sc2cdma_wt_updt_bits_entries, // @[:@16370.4]
  output [8:0]   io_sc2cdma_wmb_entries, // @[:@16370.4]
  output         io_sc2buf_wt_rd_addr_valid, // @[:@16370.4]
  output [12:0]  io_sc2buf_wt_rd_addr_bits, // @[:@16370.4]
  input          io_sc2buf_wt_rd_data_valid, // @[:@16370.4]
  input  [511:0] io_sc2buf_wt_rd_data_bits, // @[:@16370.4]
  output         io_sc2mac_wt_a_valid, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_sel_0, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_sel_1, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_sel_2, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_sel_3, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_sel_4, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_sel_5, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_sel_6, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_sel_7, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_sel_8, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_sel_9, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_sel_10, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_sel_11, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_sel_12, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_sel_13, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_sel_14, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_sel_15, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_0, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_1, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_2, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_3, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_4, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_5, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_6, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_7, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_8, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_9, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_10, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_11, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_12, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_13, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_14, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_15, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_16, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_17, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_18, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_19, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_20, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_21, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_22, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_23, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_24, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_25, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_26, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_27, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_28, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_29, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_30, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_31, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_32, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_33, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_34, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_35, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_36, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_37, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_38, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_39, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_40, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_41, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_42, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_43, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_44, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_45, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_46, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_47, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_48, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_49, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_50, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_51, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_52, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_53, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_54, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_55, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_56, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_57, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_58, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_59, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_60, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_61, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_62, // @[:@16370.4]
  output         io_sc2mac_wt_a_bits_mask_63, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_0, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_1, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_2, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_3, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_4, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_5, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_6, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_7, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_8, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_9, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_10, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_11, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_12, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_13, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_14, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_15, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_16, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_17, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_18, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_19, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_20, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_21, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_22, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_23, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_24, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_25, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_26, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_27, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_28, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_29, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_30, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_31, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_32, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_33, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_34, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_35, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_36, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_37, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_38, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_39, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_40, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_41, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_42, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_43, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_44, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_45, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_46, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_47, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_48, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_49, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_50, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_51, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_52, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_53, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_54, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_55, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_56, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_57, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_58, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_59, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_60, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_61, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_62, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_63, // @[:@16370.4]
  output         io_sc2mac_wt_b_valid, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_sel_0, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_sel_1, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_sel_2, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_sel_3, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_sel_4, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_sel_5, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_sel_6, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_sel_7, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_sel_8, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_sel_9, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_sel_10, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_sel_11, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_sel_12, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_sel_13, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_sel_14, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_sel_15, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_0, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_1, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_2, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_3, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_4, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_5, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_6, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_7, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_8, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_9, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_10, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_11, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_12, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_13, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_14, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_15, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_16, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_17, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_18, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_19, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_20, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_21, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_22, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_23, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_24, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_25, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_26, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_27, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_28, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_29, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_30, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_31, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_32, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_33, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_34, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_35, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_36, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_37, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_38, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_39, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_40, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_41, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_42, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_43, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_44, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_45, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_46, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_47, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_48, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_49, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_50, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_51, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_52, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_53, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_54, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_55, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_56, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_57, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_58, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_59, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_60, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_61, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_62, // @[:@16370.4]
  output         io_sc2mac_wt_b_bits_mask_63, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_0, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_1, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_2, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_3, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_4, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_5, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_6, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_7, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_8, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_9, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_10, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_11, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_12, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_13, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_14, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_15, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_16, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_17, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_18, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_19, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_20, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_21, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_22, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_23, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_24, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_25, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_26, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_27, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_28, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_29, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_30, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_31, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_32, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_33, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_34, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_35, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_36, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_37, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_38, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_39, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_40, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_41, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_42, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_43, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_44, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_45, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_46, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_47, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_48, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_49, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_50, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_51, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_52, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_53, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_54, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_55, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_56, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_57, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_58, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_59, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_60, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_61, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_62, // @[:@16370.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_63, // @[:@16370.4]
  input          io_reg2dp_op_en, // @[:@16370.4]
  input  [1:0]   io_reg2dp_y_extension, // @[:@16370.4]
  input          io_reg2dp_skip_weight_rls, // @[:@16370.4]
  input          io_reg2dp_weight_format, // @[:@16370.4]
  input  [31:0]  io_reg2dp_weight_bytes, // @[:@16370.4]
  input  [27:0]  io_reg2dp_wmb_bytes, // @[:@16370.4]
  input  [4:0]   io_reg2dp_data_bank, // @[:@16370.4]
  input  [4:0]   io_reg2dp_weight_bank // @[:@16370.4]
);
  wire  NV_NVDLA_CSC_WL_dec_reset; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_nvdla_core_clk; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_valid; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_0; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_1; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_2; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_3; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_4; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_5; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_6; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_7; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_8; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_9; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_10; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_11; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_12; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_13; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_14; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_15; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_16; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_17; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_18; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_19; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_20; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_21; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_22; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_23; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_24; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_25; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_26; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_27; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_28; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_29; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_30; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_31; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_32; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_33; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_34; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_35; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_36; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_37; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_38; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_39; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_40; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_41; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_42; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_43; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_44; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_45; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_46; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_47; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_48; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_49; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_50; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_51; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_52; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_53; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_54; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_55; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_56; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_57; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_58; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_59; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_60; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_61; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_62; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_63; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_0; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_1; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_2; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_3; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_4; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_5; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_6; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_7; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_8; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_9; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_10; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_11; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_12; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_13; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_14; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_15; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_16; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_17; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_18; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_19; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_20; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_21; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_22; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_23; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_24; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_25; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_26; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_27; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_28; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_29; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_30; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_31; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_32; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_33; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_34; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_35; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_36; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_37; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_38; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_39; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_40; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_41; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_42; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_43; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_44; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_45; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_46; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_47; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_48; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_49; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_50; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_51; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_52; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_53; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_54; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_55; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_56; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_57; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_58; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_59; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_60; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_61; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_62; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_63; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_0; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_1; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_2; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_3; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_4; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_5; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_6; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_7; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_8; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_9; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_10; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_11; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_12; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_13; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_14; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_15; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_16; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_17; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_18; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_19; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_20; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_21; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_22; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_23; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_24; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_25; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_26; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_27; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_28; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_29; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_30; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_31; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [9:0] NV_NVDLA_CSC_WL_dec_io_input_mask_en; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_valid; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_0; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_1; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_2; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_3; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_4; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_5; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_6; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_7; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_8; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_9; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_10; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_11; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_12; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_13; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_14; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_15; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_16; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_17; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_18; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_19; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_20; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_21; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_22; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_23; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_24; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_25; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_26; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_27; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_28; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_29; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_30; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_31; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_32; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_33; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_34; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_35; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_36; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_37; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_38; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_39; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_40; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_41; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_42; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_43; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_44; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_45; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_46; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_47; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_48; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_49; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_50; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_51; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_52; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_53; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_54; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_55; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_56; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_57; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_58; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_59; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_60; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_61; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_62; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_63; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_0; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_1; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_2; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_3; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_4; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_5; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_6; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_7; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_8; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_9; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_10; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_11; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_12; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_13; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_14; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_15; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_16; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_17; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_18; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_19; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_20; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_21; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_22; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_23; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_24; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_25; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_26; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_27; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_28; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_29; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_30; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_31; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_32; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_33; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_34; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_35; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_36; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_37; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_38; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_39; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_40; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_41; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_42; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_43; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_44; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_45; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_46; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_47; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_48; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_49; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_50; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_51; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_52; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_53; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_54; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_55; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_56; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_57; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_58; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_59; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_60; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_61; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_62; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_63; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_0; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_1; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_2; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_3; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_4; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_5; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_6; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_7; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_8; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_9; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_10; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_11; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_12; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_13; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_14; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_15; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_16; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_17; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_18; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_19; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_20; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_21; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_22; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_23; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_24; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_25; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_26; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_27; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_28; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_29; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_30; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_31; // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
  reg  _T_698; // @[NV_NVDLA_CSC_wl.scala 95:35:@16373.4]
  reg [31:0] _RAND_0;
  wire  _T_700; // @[NV_NVDLA_CSC_wl.scala 97:35:@16374.4]
  wire  _T_704; // @[NV_NVDLA_CSC_wl.scala 99:38:@16376.4]
  wire  _T_706; // @[NV_NVDLA_CSC_wl.scala 100:35:@16377.4]
  wire  _T_707; // @[NV_NVDLA_CSC_wl.scala 101:37:@16378.4]
  wire  _T_708; // @[NV_NVDLA_CSC_wl.scala 101:35:@16379.4]
  reg [4:0] _T_715; // @[NV_NVDLA_CSC_wl.scala 108:28:@16382.4]
  reg [31:0] _RAND_1;
  reg [4:0] _T_722; // @[NV_NVDLA_CSC_wl.scala 109:30:@16384.4]
  reg [31:0] _RAND_2;
  reg [14:0] _T_729; // @[NV_NVDLA_CSC_wl.scala 110:38:@16386.4]
  reg [31:0] _RAND_3;
  reg [8:0] _T_736; // @[NV_NVDLA_CSC_wl.scala 111:35:@16388.4]
  reg [31:0] _RAND_4;
  reg [2:0] _T_739; // @[NV_NVDLA_CSC_wl.scala 112:30:@16389.4]
  reg [31:0] _RAND_5;
  reg  _T_742; // @[NV_NVDLA_CSC_wl.scala 113:35:@16390.4]
  reg [31:0] _RAND_6;
  wire  _T_743; // @[NV_NVDLA_CSC_wl.scala 115:36:@16391.4]
  wire [5:0] _T_749; // @[NV_NVDLA_CSC_wl.scala 120:42:@16395.6]
  wire [4:0] _T_750; // @[NV_NVDLA_CSC_wl.scala 120:42:@16396.6]
  wire [5:0] _T_752; // @[NV_NVDLA_CSC_wl.scala 121:46:@16398.6]
  wire [4:0] _T_753; // @[NV_NVDLA_CSC_wl.scala 121:46:@16399.6]
  wire [8:0] _T_755; // @[NV_NVDLA_CSC_wl.scala 122:42:@16401.6]
  wire [2:0] _T_756; // @[NV_NVDLA_CSC_wl.scala 122:67:@16402.6]
  wire [4:0] _GEN_0; // @[NV_NVDLA_CSC_wl.scala 119:19:@16394.4]
  wire [4:0] _GEN_1; // @[NV_NVDLA_CSC_wl.scala 119:19:@16394.4]
  wire [2:0] _GEN_2; // @[NV_NVDLA_CSC_wl.scala 119:19:@16394.4]
  wire  _GEN_3; // @[NV_NVDLA_CSC_wl.scala 119:19:@16394.4]
  wire  _T_757; // @[NV_NVDLA_CSC_wl.scala 125:21:@16406.4]
  wire [14:0] _T_758; // @[NV_NVDLA_CSC_wl.scala 126:54:@16408.6]
  wire [8:0] _T_759; // @[NV_NVDLA_CSC_wl.scala 127:70:@16410.6]
  wire [8:0] _T_761; // @[NV_NVDLA_CSC_wl.scala 127:32:@16411.6]
  wire [14:0] _GEN_4; // @[NV_NVDLA_CSC_wl.scala 125:49:@16407.4]
  wire [8:0] _GEN_5; // @[NV_NVDLA_CSC_wl.scala 125:49:@16407.4]
  reg  _T_1692; // @[NV_NVDLA_CSC_wl.scala 654:76:@17206.4]
  reg [31:0] _RAND_7;
  reg [35:0] _T_1712; // @[NV_NVDLA_CSC_wl.scala 656:75:@17213.4]
  reg [63:0] _RAND_8;
  wire  _T_1759; // @[NV_NVDLA_CSC_wl.scala 693:34:@17289.4]
  wire  _T_857; // @[NV_NVDLA_CSC_wl.scala 203:36:@16489.4]
  wire  _T_858; // @[NV_NVDLA_CSC_wl.scala 207:25:@16490.4]
  wire [14:0] _T_1755; // @[NV_NVDLA_CSC_wl.scala 689:44:@17284.4]
  wire [14:0] _T_859; // @[NV_NVDLA_CSC_wl.scala 208:29:@16492.4]
  wire [8:0] _T_1754; // @[NV_NVDLA_CSC_wl.scala 688:45:@17282.4]
  wire [8:0] _T_860; // @[NV_NVDLA_CSC_wl.scala 209:30:@16494.4]
  reg [14:0] _T_798; // @[NV_NVDLA_CSC_wl.scala 153:62:@16435.4]
  reg [31:0] _RAND_9;
  wire [15:0] _T_799; // @[NV_NVDLA_CSC_wl.scala 155:39:@16436.4]
  wire [14:0] _T_800; // @[NV_NVDLA_CSC_wl.scala 155:39:@16437.4]
  wire [13:0] _T_802; // @[Cat.scala 30:58:@16438.4]
  wire [14:0] _GEN_497; // @[NV_NVDLA_CSC_wl.scala 156:48:@16439.4]
  wire [15:0] _T_803; // @[NV_NVDLA_CSC_wl.scala 156:48:@16439.4]
  wire [15:0] _T_804; // @[NV_NVDLA_CSC_wl.scala 156:48:@16440.4]
  wire [14:0] _T_805; // @[NV_NVDLA_CSC_wl.scala 156:48:@16441.4]
  wire  _T_808; // @[NV_NVDLA_CSC_wl.scala 157:48:@16443.4]
  wire  _T_810; // @[NV_NVDLA_CSC_wl.scala 158:88:@16444.4]
  wire [14:0] _T_811; // @[NV_NVDLA_CSC_wl.scala 158:113:@16445.4]
  wire [14:0] _T_812; // @[NV_NVDLA_CSC_wl.scala 158:87:@16446.4]
  wire [14:0] _T_813; // @[NV_NVDLA_CSC_wl.scala 158:28:@16447.4]
  wire  _T_847; // @[NV_NVDLA_CSC_wl.scala 184:21:@16475.4]
  wire [14:0] _GEN_8; // @[NV_NVDLA_CSC_wl.scala 184:30:@16476.4]
  reg  _T_863; // @[NV_NVDLA_CSC_wl.scala 212:40:@16496.4]
  reg [31:0] _RAND_10;
  reg [14:0] _T_867; // @[Reg.scala 19:20:@16500.4]
  reg [31:0] _RAND_11;
  wire [14:0] _GEN_12; // @[Reg.scala 20:19:@16501.4]
  reg [8:0] _T_871; // @[Reg.scala 19:20:@16506.4]
  reg [31:0] _RAND_12;
  wire [8:0] _GEN_13; // @[Reg.scala 20:19:@16507.4]
  reg  _T_877; // @[NV_NVDLA_CSC_wl.scala 223:71:@16513.4]
  reg [31:0] _RAND_13;
  reg [17:0] _T_882; // @[NV_NVDLA_CSC_wl.scala 225:67:@16515.4]
  reg [31:0] _RAND_14;
  wire  _T_879; // @[NV_NVDLA_CSC_wl.scala 224:26:@16514.4 NV_NVDLA_CSC_wl.scala 228:19:@16517.4]
  wire [17:0] _GEN_14; // @[NV_NVDLA_CSC_wl.scala 232:30:@16519.4]
  wire [6:0] _T_883; // @[NV_NVDLA_CSC_wl.scala 241:31:@16522.4]
  wire [5:0] _T_884; // @[NV_NVDLA_CSC_wl.scala 242:31:@16523.4]
  wire [1:0] _T_885; // @[NV_NVDLA_CSC_wl.scala 243:29:@16524.4]
  wire  _T_886; // @[NV_NVDLA_CSC_wl.scala 244:31:@16525.4]
  wire  _T_887; // @[NV_NVDLA_CSC_wl.scala 245:29:@16526.4]
  wire  _T_888; // @[NV_NVDLA_CSC_wl.scala 246:30:@16527.4]
  reg [4:0] _T_893; // @[NV_NVDLA_CSC_wl.scala 254:29:@16529.4]
  reg [31:0] _RAND_15;
  reg  _T_896; // @[NV_NVDLA_CSC_wl.scala 255:36:@16530.4]
  reg [31:0] _RAND_16;
  wire [5:0] _T_898; // @[NV_NVDLA_CSC_wl.scala 257:37:@16531.4]
  wire [4:0] _T_899; // @[NV_NVDLA_CSC_wl.scala 257:37:@16532.4]
  wire [4:0] _T_904; // @[NV_NVDLA_CSC_wl.scala 259:39:@16535.4]
  wire  _T_905; // @[NV_NVDLA_CSC_wl.scala 260:38:@16536.4]
  wire [4:0] _T_902; // @[NV_NVDLA_CSC_wl.scala 258:59:@16533.4]
  wire [4:0] _T_903; // @[NV_NVDLA_CSC_wl.scala 258:27:@16534.4]
  wire  _T_908; // @[NV_NVDLA_CSC_wl.scala 262:64:@16538.4]
  wire  _T_909; // @[NV_NVDLA_CSC_wl.scala 262:51:@16539.4]
  wire  _T_911; // @[NV_NVDLA_CSC_wl.scala 262:50:@16540.4]
  wire  _T_912; // @[NV_NVDLA_CSC_wl.scala 262:29:@16541.4]
  wire  _T_913; // @[NV_NVDLA_CSC_wl.scala 263:38:@16542.4]
  wire [4:0] _GEN_15; // @[NV_NVDLA_CSC_wl.scala 265:28:@16543.4]
  reg [10:0] _T_920; // @[NV_NVDLA_CSC_wl.scala 272:34:@16548.4]
  reg [31:0] _RAND_17;
  reg [10:0] _T_923; // @[NV_NVDLA_CSC_wl.scala 273:39:@16549.4]
  reg [31:0] _RAND_18;
  wire  _T_966; // @[NV_NVDLA_CSC_wl.scala 289:37:@16580.4]
  wire  _T_964; // @[Mux.scala 46:19:@16577.4]
  wire [7:0] _T_942; // @[Cat.scala 30:58:@16563.4]
  wire  _T_962; // @[Mux.scala 46:19:@16575.4]
  wire [6:0] _T_951; // @[NV_NVDLA_CSC_wl.scala 285:101:@16567.4]
  wire [8:0] _T_954; // @[Cat.scala 30:58:@16569.4]
  wire  _T_960; // @[Mux.scala 46:19:@16573.4]
  wire [7:0] _T_958; // @[Cat.scala 30:58:@16571.4]
  wire [8:0] _T_959; // @[NV_NVDLA_CSC_wl.scala 286:109:@16572.4]
  wire [5:0] _T_944; // @[NV_NVDLA_CSC_wl.scala 282:92:@16564.4]
  wire [8:0] _T_947; // @[Cat.scala 30:58:@16566.4]
  wire [8:0] _T_961; // @[Mux.scala 46:16:@16574.4]
  wire [8:0] _T_963; // @[Mux.scala 46:16:@16576.4]
  wire [8:0] _T_965; // @[Mux.scala 46:16:@16578.4]
  wire [7:0] _T_917; // @[NV_NVDLA_CSC_wl.scala 271:31:@16547.4 NV_NVDLA_CSC_wl.scala 282:21:@16579.4]
  wire [10:0] _T_968; // @[Cat.scala 30:58:@16581.4]
  wire  _T_969; // @[NV_NVDLA_CSC_wl.scala 289:75:@16582.4]
  wire  _T_970; // @[NV_NVDLA_CSC_wl.scala 289:56:@16583.4]
  wire  _T_924; // @[NV_NVDLA_CSC_wl.scala 275:35:@16550.4]
  wire [10:0] _T_927; // @[NV_NVDLA_CSC_wl.scala 275:34:@16551.4]
  wire [7:0] _T_929; // @[NV_NVDLA_CSC_wl.scala 276:34:@16552.4]
  wire [11:0] _T_930; // @[NV_NVDLA_CSC_wl.scala 277:47:@16553.4]
  wire [10:0] _T_931; // @[NV_NVDLA_CSC_wl.scala 277:47:@16554.4]
  wire [10:0] _GEN_501; // @[NV_NVDLA_CSC_wl.scala 277:69:@16555.4]
  wire [11:0] _T_932; // @[NV_NVDLA_CSC_wl.scala 277:69:@16555.4]
  wire [11:0] _T_933; // @[NV_NVDLA_CSC_wl.scala 277:69:@16556.4]
  wire [10:0] _T_934; // @[NV_NVDLA_CSC_wl.scala 277:69:@16557.4]
  wire  _T_936; // @[NV_NVDLA_CSC_wl.scala 278:82:@16558.4]
  wire  _T_937; // @[NV_NVDLA_CSC_wl.scala 278:80:@16559.4]
  wire  _T_938; // @[NV_NVDLA_CSC_wl.scala 278:96:@16560.4]
  wire [10:0] _T_939; // @[NV_NVDLA_CSC_wl.scala 278:65:@16561.4]
  wire [10:0] _T_940; // @[NV_NVDLA_CSC_wl.scala 278:32:@16562.4]
  wire  _T_972; // @[NV_NVDLA_CSC_wl.scala 290:43:@16586.4]
  wire  _T_974; // @[NV_NVDLA_CSC_wl.scala 291:85:@16588.4]
  wire  _T_975; // @[NV_NVDLA_CSC_wl.scala 291:101:@16589.4]
  wire  _T_976; // @[NV_NVDLA_CSC_wl.scala 291:48:@16590.4]
  wire [10:0] _GEN_16; // @[NV_NVDLA_CSC_wl.scala 293:33:@16591.4]
  wire [10:0] _GEN_17; // @[NV_NVDLA_CSC_wl.scala 296:38:@16594.4]
  reg  _T_1003; // @[NV_NVDLA_CSC_wl.scala 318:34:@16622.4]
  reg [31:0] _RAND_19;
  reg [8:0] _T_1006; // @[NV_NVDLA_CSC_wl.scala 319:30:@16623.4]
  reg [31:0] _RAND_20;
  wire  _T_1007; // @[NV_NVDLA_CSC_wl.scala 321:58:@16624.4]
  wire  _T_1008; // @[NV_NVDLA_CSC_wl.scala 321:42:@16625.4]
  wire  _T_1010; // @[NV_NVDLA_CSC_wl.scala 322:48:@16626.4]
  wire  _T_1012; // @[NV_NVDLA_CSC_wl.scala 322:32:@16627.4]
  wire  _T_1013; // @[NV_NVDLA_CSC_wl.scala 321:32:@16628.4]
  wire [9:0] _T_1015; // @[NV_NVDLA_CSC_wl.scala 323:39:@16629.4]
  wire [8:0] _T_1016; // @[NV_NVDLA_CSC_wl.scala 323:39:@16630.4]
  wire  _T_1018; // @[NV_NVDLA_CSC_wl.scala 325:43:@16631.4]
  wire [8:0] _T_1020; // @[NV_NVDLA_CSC_wl.scala 325:28:@16632.4]
  wire [8:0] _T_1021; // @[NV_NVDLA_CSC_wl.scala 324:28:@16633.4]
  wire  _T_1022; // @[NV_NVDLA_CSC_wl.scala 326:58:@16634.4]
  wire  _T_1023; // @[NV_NVDLA_CSC_wl.scala 326:75:@16635.4]
  wire  _T_1024; // @[NV_NVDLA_CSC_wl.scala 326:91:@16636.4]
  wire  _T_1025; // @[NV_NVDLA_CSC_wl.scala 326:39:@16637.4]
  wire  _T_1026; // @[NV_NVDLA_CSC_wl.scala 326:126:@16638.4]
  wire  _T_1027; // @[NV_NVDLA_CSC_wl.scala 326:144:@16639.4]
  wire  _T_1028; // @[NV_NVDLA_CSC_wl.scala 326:142:@16640.4]
  wire  _T_1029; // @[NV_NVDLA_CSC_wl.scala 326:107:@16641.4]
  wire  _T_1031; // @[NV_NVDLA_CSC_wl.scala 327:47:@16643.4]
  wire [8:0] _T_1032; // @[NV_NVDLA_CSC_wl.scala 327:30:@16644.4]
  wire [8:0] _GEN_20; // @[NV_NVDLA_CSC_wl.scala 330:29:@16646.4]
  reg [6:0] _T_1041; // @[NV_NVDLA_CSC_wl.scala 337:41:@16651.4]
  reg [31:0] _RAND_21;
  reg [7:0] _T_1044; // @[NV_NVDLA_CSC_wl.scala 338:37:@16652.4]
  reg [31:0] _RAND_22;
  reg [8:0] _T_1047; // @[NV_NVDLA_CSC_wl.scala 339:41:@16653.4]
  reg [31:0] _RAND_23;
  reg  _T_1050; // @[NV_NVDLA_CSC_wl.scala 340:40:@16654.4]
  reg [31:0] _RAND_24;
  reg  _T_1053; // @[NV_NVDLA_CSC_wl.scala 341:41:@16655.4]
  reg [31:0] _RAND_25;
  reg  _T_1056; // @[NV_NVDLA_CSC_wl.scala 342:39:@16656.4]
  reg [31:0] _RAND_26;
  reg  _T_1059; // @[NV_NVDLA_CSC_wl.scala 343:33:@16657.4]
  reg [31:0] _RAND_27;
  reg [1:0] _T_1062; // @[NV_NVDLA_CSC_wl.scala 344:39:@16658.4]
  reg [31:0] _RAND_28;
  wire [6:0] _GEN_22; // @[NV_NVDLA_CSC_wl.scala 351:25:@16664.4]
  wire [7:0] _GEN_23; // @[NV_NVDLA_CSC_wl.scala 351:25:@16664.4]
  wire  _T_1063; // @[NV_NVDLA_CSC_wl.scala 355:25:@16668.4]
  wire  _T_1064; // @[NV_NVDLA_CSC_wl.scala 355:41:@16669.4]
  wire [8:0] _GEN_24; // @[NV_NVDLA_CSC_wl.scala 355:57:@16670.4]
  wire  _T_1067; // @[NV_NVDLA_CSC_wl.scala 362:41:@16679.6]
  wire  _GEN_25; // @[NV_NVDLA_CSC_wl.scala 358:25:@16673.4]
  wire  _GEN_26; // @[NV_NVDLA_CSC_wl.scala 358:25:@16673.4]
  wire  _GEN_27; // @[NV_NVDLA_CSC_wl.scala 358:25:@16673.4]
  wire  _GEN_28; // @[NV_NVDLA_CSC_wl.scala 358:25:@16673.4]
  wire [1:0] _GEN_29; // @[NV_NVDLA_CSC_wl.scala 358:25:@16673.4]
  wire [30:0] _T_1076; // @[Cat.scala 30:58:@16690.4]
  reg  _T_1081; // @[NV_NVDLA_CSC_wl.scala 385:77:@16692.4]
  reg [31:0] _RAND_29;
  reg  _T_1084; // @[NV_NVDLA_CSC_wl.scala 385:77:@16693.4]
  reg [31:0] _RAND_30;
  reg  _T_1087; // @[NV_NVDLA_CSC_wl.scala 385:77:@16694.4]
  reg [31:0] _RAND_31;
  reg  _T_1090; // @[NV_NVDLA_CSC_wl.scala 385:77:@16695.4]
  reg [31:0] _RAND_32;
  reg  _T_1093; // @[NV_NVDLA_CSC_wl.scala 385:77:@16696.4]
  reg [31:0] _RAND_33;
  reg  _T_1096; // @[NV_NVDLA_CSC_wl.scala 385:77:@16697.4]
  reg [31:0] _RAND_34;
  reg [30:0] _T_1101; // @[NV_NVDLA_CSC_wl.scala 387:75:@16699.4]
  reg [31:0] _RAND_35;
  reg [30:0] _T_1104; // @[NV_NVDLA_CSC_wl.scala 387:75:@16700.4]
  reg [31:0] _RAND_36;
  reg [30:0] _T_1107; // @[NV_NVDLA_CSC_wl.scala 387:75:@16701.4]
  reg [31:0] _RAND_37;
  reg [30:0] _T_1110; // @[NV_NVDLA_CSC_wl.scala 387:75:@16702.4]
  reg [31:0] _RAND_38;
  reg [30:0] _T_1113; // @[NV_NVDLA_CSC_wl.scala 387:75:@16703.4]
  reg [31:0] _RAND_39;
  reg [30:0] _T_1116; // @[NV_NVDLA_CSC_wl.scala 387:75:@16704.4]
  reg [31:0] _RAND_40;
  wire [30:0] _GEN_30; // @[NV_NVDLA_CSC_wl.scala 394:37:@16708.4]
  wire [30:0] _GEN_31; // @[NV_NVDLA_CSC_wl.scala 394:37:@16712.4]
  wire [30:0] _GEN_32; // @[NV_NVDLA_CSC_wl.scala 394:37:@16716.4]
  wire [30:0] _GEN_33; // @[NV_NVDLA_CSC_wl.scala 394:37:@16720.4]
  wire [30:0] _GEN_34; // @[NV_NVDLA_CSC_wl.scala 394:37:@16724.4]
  wire [30:0] _GEN_35; // @[NV_NVDLA_CSC_wl.scala 394:37:@16728.4]
  wire [6:0] _T_1117; // @[NV_NVDLA_CSC_wl.scala 404:46:@16731.4]
  wire [7:0] _T_1118; // @[NV_NVDLA_CSC_wl.scala 405:42:@16732.4]
  wire [8:0] _T_1119; // @[NV_NVDLA_CSC_wl.scala 406:46:@16733.4]
  wire  _T_1120; // @[NV_NVDLA_CSC_wl.scala 407:45:@16734.4]
  wire  _T_1121; // @[NV_NVDLA_CSC_wl.scala 408:46:@16735.4]
  wire  _T_1122; // @[NV_NVDLA_CSC_wl.scala 409:44:@16736.4]
  wire  _T_1123; // @[NV_NVDLA_CSC_wl.scala 410:38:@16737.4]
  wire [1:0] _T_1124; // @[NV_NVDLA_CSC_wl.scala 411:44:@16738.4]
  wire  _T_1137; // @[NV_NVDLA_CSC_wl.scala 421:91:@16743.4]
  wire  _T_1138; // @[NV_NVDLA_CSC_wl.scala 421:89:@16744.4]
  wire  _T_1145; // @[NV_NVDLA_CSC_wl.scala 422:72:@16751.4]
  wire  _T_1146; // @[NV_NVDLA_CSC_wl.scala 422:92:@16752.4]
  wire  _T_1147; // @[NV_NVDLA_CSC_wl.scala 422:51:@16753.4]
  wire  _T_1148; // @[NV_NVDLA_CSC_wl.scala 424:40:@16754.4]
  wire  _T_1149; // @[NV_NVDLA_CSC_wl.scala 424:19:@16755.4]
  reg [318:0] _T_1156; // @[NV_NVDLA_CSC_wl.scala 433:31:@16763.4]
  reg [319:0] _RAND_41;
  reg [511:0] _T_1163; // @[NV_NVDLA_CSC_wl.scala 434:35:@16765.4]
  reg [511:0] _RAND_42;
  wire [63:0] _T_1170; // @[NV_NVDLA_CSC_wl.scala 437:63:@16771.4]
  wire [190:0] _T_1171; // @[NV_NVDLA_CSC_wl.scala 437:45:@16772.4]
  wire  _T_1172; // @[NV_NVDLA_CSC_wl.scala 437:108:@16773.4]
  wire [63:0] _T_1176; // @[Bitwise.scala 72:12:@16775.4]
  wire [190:0] _GEN_503; // @[NV_NVDLA_CSC_wl.scala 437:85:@16776.4]
  wire [190:0] _T_1177; // @[NV_NVDLA_CSC_wl.scala 437:85:@16776.4]
  wire [318:0] _T_1183; // @[NV_NVDLA_CSC_wl.scala 438:56:@16778.4]
  wire [318:0] _T_1184; // @[NV_NVDLA_CSC_wl.scala 438:25:@16779.4]
  wire [63:0] _T_1185; // @[NV_NVDLA_CSC_wl.scala 439:41:@16780.4]
  wire [318:0] _GEN_504; // @[NV_NVDLA_CSC_wl.scala 439:63:@16781.4]
  wire [318:0] _T_1186; // @[NV_NVDLA_CSC_wl.scala 439:63:@16781.4]
  wire [318:0] _GEN_38; // @[NV_NVDLA_CSC_wl.scala 441:28:@16782.4]
  reg [511:0] _T_1193; // @[NV_NVDLA_CSC_wl.scala 447:40:@16786.4]
  reg [511:0] _RAND_43;
  wire [511:0] _T_1199; // @[NV_NVDLA_CSC_wl.scala 450:49:@16792.4]
  wire [511:0] _T_1208; // @[NV_NVDLA_CSC_wl.scala 453:84:@16797.4]
  wire [511:0] _T_1209; // @[NV_NVDLA_CSC_wl.scala 453:33:@16798.4]
  wire [4:0] _T_1215; // @[NV_NVDLA_CSC_wl.scala 456:52:@16804.4]
  wire [5:0] _T_1217; // @[Cat.scala 30:58:@16805.4]
  wire [5:0] _GEN_506; // @[NV_NVDLA_CSC_wl.scala 456:69:@16807.4]
  wire [6:0] _T_1219; // @[NV_NVDLA_CSC_wl.scala 456:69:@16807.4]
  wire [5:0] _T_1220; // @[NV_NVDLA_CSC_wl.scala 456:69:@16808.4]
  wire [511:0] _GEN_39; // @[NV_NVDLA_CSC_wl.scala 458:34:@16809.4]
  wire [511:0] _GEN_40; // @[NV_NVDLA_CSC_wl.scala 461:39:@16812.4]
  reg  _T_1223; // @[NV_NVDLA_CSC_wl.scala 466:36:@16815.4]
  reg [31:0] _RAND_44;
  reg [6:0] _T_1226; // @[NV_NVDLA_CSC_wl.scala 467:37:@16816.4]
  reg [31:0] _RAND_45;
  reg  _T_1229; // @[NV_NVDLA_CSC_wl.scala 468:36:@16817.4]
  reg [31:0] _RAND_46;
  reg  _T_1232; // @[NV_NVDLA_CSC_wl.scala 469:37:@16818.4]
  reg [31:0] _RAND_47;
  reg  _T_1235; // @[NV_NVDLA_CSC_wl.scala 470:35:@16819.4]
  reg [31:0] _RAND_48;
  reg  _T_1238; // @[NV_NVDLA_CSC_wl.scala 471:29:@16820.4]
  reg [31:0] _RAND_49;
  reg [8:0] _T_1241; // @[NV_NVDLA_CSC_wl.scala 472:41:@16821.4]
  reg [31:0] _RAND_50;
  reg [1:0] _T_1244; // @[NV_NVDLA_CSC_wl.scala 473:35:@16822.4]
  reg [31:0] _RAND_51;
  reg [6:0] _T_1247; // @[NV_NVDLA_CSC_wl.scala 474:35:@16823.4]
  reg [31:0] _RAND_52;
  wire [6:0] _GEN_41; // @[NV_NVDLA_CSC_wl.scala 477:28:@16825.4]
  wire  _GEN_42; // @[NV_NVDLA_CSC_wl.scala 477:28:@16825.4]
  wire  _GEN_43; // @[NV_NVDLA_CSC_wl.scala 477:28:@16825.4]
  wire  _GEN_44; // @[NV_NVDLA_CSC_wl.scala 477:28:@16825.4]
  wire  _GEN_45; // @[NV_NVDLA_CSC_wl.scala 477:28:@16825.4]
  wire [8:0] _GEN_46; // @[NV_NVDLA_CSC_wl.scala 477:28:@16825.4]
  wire [1:0] _GEN_47; // @[NV_NVDLA_CSC_wl.scala 477:28:@16825.4]
  wire [6:0] _GEN_48; // @[NV_NVDLA_CSC_wl.scala 477:28:@16825.4]
  wire  _T_1318; // @[NV_NVDLA_CSC_wl.scala 497:40:@16836.4]
  wire  _T_1319; // @[NV_NVDLA_CSC_wl.scala 497:40:@16838.4]
  wire  _T_1320; // @[NV_NVDLA_CSC_wl.scala 497:40:@16840.4]
  wire  _T_1321; // @[NV_NVDLA_CSC_wl.scala 497:40:@16842.4]
  wire  _T_1322; // @[NV_NVDLA_CSC_wl.scala 497:40:@16844.4]
  wire  _T_1323; // @[NV_NVDLA_CSC_wl.scala 497:40:@16846.4]
  wire  _T_1324; // @[NV_NVDLA_CSC_wl.scala 497:40:@16848.4]
  wire  _T_1325; // @[NV_NVDLA_CSC_wl.scala 497:40:@16850.4]
  wire  _T_1326; // @[NV_NVDLA_CSC_wl.scala 497:40:@16852.4]
  wire  _T_1327; // @[NV_NVDLA_CSC_wl.scala 497:40:@16854.4]
  wire  _T_1328; // @[NV_NVDLA_CSC_wl.scala 497:40:@16856.4]
  wire  _T_1329; // @[NV_NVDLA_CSC_wl.scala 497:40:@16858.4]
  wire  _T_1330; // @[NV_NVDLA_CSC_wl.scala 497:40:@16860.4]
  wire  _T_1331; // @[NV_NVDLA_CSC_wl.scala 497:40:@16862.4]
  wire  _T_1332; // @[NV_NVDLA_CSC_wl.scala 497:40:@16864.4]
  wire  _T_1333; // @[NV_NVDLA_CSC_wl.scala 497:40:@16866.4]
  wire  _T_1334; // @[NV_NVDLA_CSC_wl.scala 497:40:@16868.4]
  wire  _T_1335; // @[NV_NVDLA_CSC_wl.scala 497:40:@16870.4]
  wire  _T_1336; // @[NV_NVDLA_CSC_wl.scala 497:40:@16872.4]
  wire  _T_1337; // @[NV_NVDLA_CSC_wl.scala 497:40:@16874.4]
  wire  _T_1338; // @[NV_NVDLA_CSC_wl.scala 497:40:@16876.4]
  wire  _T_1339; // @[NV_NVDLA_CSC_wl.scala 497:40:@16878.4]
  wire  _T_1340; // @[NV_NVDLA_CSC_wl.scala 497:40:@16880.4]
  wire  _T_1341; // @[NV_NVDLA_CSC_wl.scala 497:40:@16882.4]
  wire  _T_1342; // @[NV_NVDLA_CSC_wl.scala 497:40:@16884.4]
  wire  _T_1343; // @[NV_NVDLA_CSC_wl.scala 497:40:@16886.4]
  wire  _T_1344; // @[NV_NVDLA_CSC_wl.scala 497:40:@16888.4]
  wire  _T_1345; // @[NV_NVDLA_CSC_wl.scala 497:40:@16890.4]
  wire  _T_1346; // @[NV_NVDLA_CSC_wl.scala 497:40:@16892.4]
  wire  _T_1347; // @[NV_NVDLA_CSC_wl.scala 497:40:@16894.4]
  wire  _T_1348; // @[NV_NVDLA_CSC_wl.scala 497:40:@16896.4]
  wire  _T_1349; // @[NV_NVDLA_CSC_wl.scala 497:40:@16898.4]
  wire  _T_1350; // @[NV_NVDLA_CSC_wl.scala 497:40:@16900.4]
  wire  _T_1351; // @[NV_NVDLA_CSC_wl.scala 497:40:@16902.4]
  wire  _T_1352; // @[NV_NVDLA_CSC_wl.scala 497:40:@16904.4]
  wire  _T_1353; // @[NV_NVDLA_CSC_wl.scala 497:40:@16906.4]
  wire  _T_1354; // @[NV_NVDLA_CSC_wl.scala 497:40:@16908.4]
  wire  _T_1355; // @[NV_NVDLA_CSC_wl.scala 497:40:@16910.4]
  wire  _T_1356; // @[NV_NVDLA_CSC_wl.scala 497:40:@16912.4]
  wire  _T_1357; // @[NV_NVDLA_CSC_wl.scala 497:40:@16914.4]
  wire  _T_1358; // @[NV_NVDLA_CSC_wl.scala 497:40:@16916.4]
  wire  _T_1359; // @[NV_NVDLA_CSC_wl.scala 497:40:@16918.4]
  wire  _T_1360; // @[NV_NVDLA_CSC_wl.scala 497:40:@16920.4]
  wire  _T_1361; // @[NV_NVDLA_CSC_wl.scala 497:40:@16922.4]
  wire  _T_1362; // @[NV_NVDLA_CSC_wl.scala 497:40:@16924.4]
  wire  _T_1363; // @[NV_NVDLA_CSC_wl.scala 497:40:@16926.4]
  wire  _T_1364; // @[NV_NVDLA_CSC_wl.scala 497:40:@16928.4]
  wire  _T_1365; // @[NV_NVDLA_CSC_wl.scala 497:40:@16930.4]
  wire  _T_1366; // @[NV_NVDLA_CSC_wl.scala 497:40:@16932.4]
  wire  _T_1367; // @[NV_NVDLA_CSC_wl.scala 497:40:@16934.4]
  wire  _T_1368; // @[NV_NVDLA_CSC_wl.scala 497:40:@16936.4]
  wire  _T_1369; // @[NV_NVDLA_CSC_wl.scala 497:40:@16938.4]
  wire  _T_1370; // @[NV_NVDLA_CSC_wl.scala 497:40:@16940.4]
  wire  _T_1371; // @[NV_NVDLA_CSC_wl.scala 497:40:@16942.4]
  wire  _T_1372; // @[NV_NVDLA_CSC_wl.scala 497:40:@16944.4]
  wire  _T_1373; // @[NV_NVDLA_CSC_wl.scala 497:40:@16946.4]
  wire  _T_1374; // @[NV_NVDLA_CSC_wl.scala 497:40:@16948.4]
  wire  _T_1375; // @[NV_NVDLA_CSC_wl.scala 497:40:@16950.4]
  wire  _T_1376; // @[NV_NVDLA_CSC_wl.scala 497:40:@16952.4]
  wire  _T_1377; // @[NV_NVDLA_CSC_wl.scala 497:40:@16954.4]
  wire  _T_1378; // @[NV_NVDLA_CSC_wl.scala 497:40:@16956.4]
  wire  _T_1379; // @[NV_NVDLA_CSC_wl.scala 497:40:@16958.4]
  wire  _T_1380; // @[NV_NVDLA_CSC_wl.scala 497:40:@16960.4]
  wire  _T_1381; // @[NV_NVDLA_CSC_wl.scala 497:40:@16962.4]
  wire [1:0] _T_1382; // @[NV_NVDLA_CSC_wl.scala 499:46:@16964.4]
  wire [1:0] _GEN_507; // @[NV_NVDLA_CSC_wl.scala 499:46:@16965.4]
  wire [2:0] _T_1383; // @[NV_NVDLA_CSC_wl.scala 499:46:@16965.4]
  wire [2:0] _GEN_508; // @[NV_NVDLA_CSC_wl.scala 499:46:@16966.4]
  wire [3:0] _T_1384; // @[NV_NVDLA_CSC_wl.scala 499:46:@16966.4]
  wire [3:0] _GEN_509; // @[NV_NVDLA_CSC_wl.scala 499:46:@16967.4]
  wire [4:0] _T_1385; // @[NV_NVDLA_CSC_wl.scala 499:46:@16967.4]
  wire [4:0] _GEN_510; // @[NV_NVDLA_CSC_wl.scala 499:46:@16968.4]
  wire [5:0] _T_1386; // @[NV_NVDLA_CSC_wl.scala 499:46:@16968.4]
  wire [5:0] _GEN_511; // @[NV_NVDLA_CSC_wl.scala 499:46:@16969.4]
  wire [6:0] _T_1387; // @[NV_NVDLA_CSC_wl.scala 499:46:@16969.4]
  wire [6:0] _GEN_512; // @[NV_NVDLA_CSC_wl.scala 499:46:@16970.4]
  wire [7:0] _T_1388; // @[NV_NVDLA_CSC_wl.scala 499:46:@16970.4]
  wire [7:0] _GEN_513; // @[NV_NVDLA_CSC_wl.scala 499:46:@16971.4]
  wire [8:0] _T_1389; // @[NV_NVDLA_CSC_wl.scala 499:46:@16971.4]
  wire [8:0] _GEN_514; // @[NV_NVDLA_CSC_wl.scala 499:46:@16972.4]
  wire [9:0] _T_1390; // @[NV_NVDLA_CSC_wl.scala 499:46:@16972.4]
  wire [9:0] _GEN_515; // @[NV_NVDLA_CSC_wl.scala 499:46:@16973.4]
  wire [10:0] _T_1391; // @[NV_NVDLA_CSC_wl.scala 499:46:@16973.4]
  wire [10:0] _GEN_516; // @[NV_NVDLA_CSC_wl.scala 499:46:@16974.4]
  wire [11:0] _T_1392; // @[NV_NVDLA_CSC_wl.scala 499:46:@16974.4]
  wire [11:0] _GEN_517; // @[NV_NVDLA_CSC_wl.scala 499:46:@16975.4]
  wire [12:0] _T_1393; // @[NV_NVDLA_CSC_wl.scala 499:46:@16975.4]
  wire [12:0] _GEN_518; // @[NV_NVDLA_CSC_wl.scala 499:46:@16976.4]
  wire [13:0] _T_1394; // @[NV_NVDLA_CSC_wl.scala 499:46:@16976.4]
  wire [13:0] _GEN_519; // @[NV_NVDLA_CSC_wl.scala 499:46:@16977.4]
  wire [14:0] _T_1395; // @[NV_NVDLA_CSC_wl.scala 499:46:@16977.4]
  wire [14:0] _GEN_520; // @[NV_NVDLA_CSC_wl.scala 499:46:@16978.4]
  wire [15:0] _T_1396; // @[NV_NVDLA_CSC_wl.scala 499:46:@16978.4]
  wire [15:0] _GEN_521; // @[NV_NVDLA_CSC_wl.scala 499:46:@16979.4]
  wire [16:0] _T_1397; // @[NV_NVDLA_CSC_wl.scala 499:46:@16979.4]
  wire [16:0] _GEN_522; // @[NV_NVDLA_CSC_wl.scala 499:46:@16980.4]
  wire [17:0] _T_1398; // @[NV_NVDLA_CSC_wl.scala 499:46:@16980.4]
  wire [17:0] _GEN_523; // @[NV_NVDLA_CSC_wl.scala 499:46:@16981.4]
  wire [18:0] _T_1399; // @[NV_NVDLA_CSC_wl.scala 499:46:@16981.4]
  wire [18:0] _GEN_524; // @[NV_NVDLA_CSC_wl.scala 499:46:@16982.4]
  wire [19:0] _T_1400; // @[NV_NVDLA_CSC_wl.scala 499:46:@16982.4]
  wire [19:0] _GEN_525; // @[NV_NVDLA_CSC_wl.scala 499:46:@16983.4]
  wire [20:0] _T_1401; // @[NV_NVDLA_CSC_wl.scala 499:46:@16983.4]
  wire [20:0] _GEN_526; // @[NV_NVDLA_CSC_wl.scala 499:46:@16984.4]
  wire [21:0] _T_1402; // @[NV_NVDLA_CSC_wl.scala 499:46:@16984.4]
  wire [21:0] _GEN_527; // @[NV_NVDLA_CSC_wl.scala 499:46:@16985.4]
  wire [22:0] _T_1403; // @[NV_NVDLA_CSC_wl.scala 499:46:@16985.4]
  wire [22:0] _GEN_528; // @[NV_NVDLA_CSC_wl.scala 499:46:@16986.4]
  wire [23:0] _T_1404; // @[NV_NVDLA_CSC_wl.scala 499:46:@16986.4]
  wire [23:0] _GEN_529; // @[NV_NVDLA_CSC_wl.scala 499:46:@16987.4]
  wire [24:0] _T_1405; // @[NV_NVDLA_CSC_wl.scala 499:46:@16987.4]
  wire [24:0] _GEN_530; // @[NV_NVDLA_CSC_wl.scala 499:46:@16988.4]
  wire [25:0] _T_1406; // @[NV_NVDLA_CSC_wl.scala 499:46:@16988.4]
  wire [25:0] _GEN_531; // @[NV_NVDLA_CSC_wl.scala 499:46:@16989.4]
  wire [26:0] _T_1407; // @[NV_NVDLA_CSC_wl.scala 499:46:@16989.4]
  wire [26:0] _GEN_532; // @[NV_NVDLA_CSC_wl.scala 499:46:@16990.4]
  wire [27:0] _T_1408; // @[NV_NVDLA_CSC_wl.scala 499:46:@16990.4]
  wire [27:0] _GEN_533; // @[NV_NVDLA_CSC_wl.scala 499:46:@16991.4]
  wire [28:0] _T_1409; // @[NV_NVDLA_CSC_wl.scala 499:46:@16991.4]
  wire [28:0] _GEN_534; // @[NV_NVDLA_CSC_wl.scala 499:46:@16992.4]
  wire [29:0] _T_1410; // @[NV_NVDLA_CSC_wl.scala 499:46:@16992.4]
  wire [29:0] _GEN_535; // @[NV_NVDLA_CSC_wl.scala 499:46:@16993.4]
  wire [30:0] _T_1411; // @[NV_NVDLA_CSC_wl.scala 499:46:@16993.4]
  wire [30:0] _GEN_536; // @[NV_NVDLA_CSC_wl.scala 499:46:@16994.4]
  wire [31:0] _T_1412; // @[NV_NVDLA_CSC_wl.scala 499:46:@16994.4]
  wire [31:0] _GEN_537; // @[NV_NVDLA_CSC_wl.scala 499:46:@16995.4]
  wire [32:0] _T_1413; // @[NV_NVDLA_CSC_wl.scala 499:46:@16995.4]
  wire [32:0] _GEN_538; // @[NV_NVDLA_CSC_wl.scala 499:46:@16996.4]
  wire [33:0] _T_1414; // @[NV_NVDLA_CSC_wl.scala 499:46:@16996.4]
  wire [33:0] _GEN_539; // @[NV_NVDLA_CSC_wl.scala 499:46:@16997.4]
  wire [34:0] _T_1415; // @[NV_NVDLA_CSC_wl.scala 499:46:@16997.4]
  wire [34:0] _GEN_540; // @[NV_NVDLA_CSC_wl.scala 499:46:@16998.4]
  wire [35:0] _T_1416; // @[NV_NVDLA_CSC_wl.scala 499:46:@16998.4]
  wire [35:0] _GEN_541; // @[NV_NVDLA_CSC_wl.scala 499:46:@16999.4]
  wire [36:0] _T_1417; // @[NV_NVDLA_CSC_wl.scala 499:46:@16999.4]
  wire [36:0] _GEN_542; // @[NV_NVDLA_CSC_wl.scala 499:46:@17000.4]
  wire [37:0] _T_1418; // @[NV_NVDLA_CSC_wl.scala 499:46:@17000.4]
  wire [37:0] _GEN_543; // @[NV_NVDLA_CSC_wl.scala 499:46:@17001.4]
  wire [38:0] _T_1419; // @[NV_NVDLA_CSC_wl.scala 499:46:@17001.4]
  wire [38:0] _GEN_544; // @[NV_NVDLA_CSC_wl.scala 499:46:@17002.4]
  wire [39:0] _T_1420; // @[NV_NVDLA_CSC_wl.scala 499:46:@17002.4]
  wire [39:0] _GEN_545; // @[NV_NVDLA_CSC_wl.scala 499:46:@17003.4]
  wire [40:0] _T_1421; // @[NV_NVDLA_CSC_wl.scala 499:46:@17003.4]
  wire [40:0] _GEN_546; // @[NV_NVDLA_CSC_wl.scala 499:46:@17004.4]
  wire [41:0] _T_1422; // @[NV_NVDLA_CSC_wl.scala 499:46:@17004.4]
  wire [41:0] _GEN_547; // @[NV_NVDLA_CSC_wl.scala 499:46:@17005.4]
  wire [42:0] _T_1423; // @[NV_NVDLA_CSC_wl.scala 499:46:@17005.4]
  wire [42:0] _GEN_548; // @[NV_NVDLA_CSC_wl.scala 499:46:@17006.4]
  wire [43:0] _T_1424; // @[NV_NVDLA_CSC_wl.scala 499:46:@17006.4]
  wire [43:0] _GEN_549; // @[NV_NVDLA_CSC_wl.scala 499:46:@17007.4]
  wire [44:0] _T_1425; // @[NV_NVDLA_CSC_wl.scala 499:46:@17007.4]
  wire [44:0] _GEN_550; // @[NV_NVDLA_CSC_wl.scala 499:46:@17008.4]
  wire [45:0] _T_1426; // @[NV_NVDLA_CSC_wl.scala 499:46:@17008.4]
  wire [45:0] _GEN_551; // @[NV_NVDLA_CSC_wl.scala 499:46:@17009.4]
  wire [46:0] _T_1427; // @[NV_NVDLA_CSC_wl.scala 499:46:@17009.4]
  wire [46:0] _GEN_552; // @[NV_NVDLA_CSC_wl.scala 499:46:@17010.4]
  wire [47:0] _T_1428; // @[NV_NVDLA_CSC_wl.scala 499:46:@17010.4]
  wire [47:0] _GEN_553; // @[NV_NVDLA_CSC_wl.scala 499:46:@17011.4]
  wire [48:0] _T_1429; // @[NV_NVDLA_CSC_wl.scala 499:46:@17011.4]
  wire [48:0] _GEN_554; // @[NV_NVDLA_CSC_wl.scala 499:46:@17012.4]
  wire [49:0] _T_1430; // @[NV_NVDLA_CSC_wl.scala 499:46:@17012.4]
  wire [49:0] _GEN_555; // @[NV_NVDLA_CSC_wl.scala 499:46:@17013.4]
  wire [50:0] _T_1431; // @[NV_NVDLA_CSC_wl.scala 499:46:@17013.4]
  wire [50:0] _GEN_556; // @[NV_NVDLA_CSC_wl.scala 499:46:@17014.4]
  wire [51:0] _T_1432; // @[NV_NVDLA_CSC_wl.scala 499:46:@17014.4]
  wire [51:0] _GEN_557; // @[NV_NVDLA_CSC_wl.scala 499:46:@17015.4]
  wire [52:0] _T_1433; // @[NV_NVDLA_CSC_wl.scala 499:46:@17015.4]
  wire [52:0] _GEN_558; // @[NV_NVDLA_CSC_wl.scala 499:46:@17016.4]
  wire [53:0] _T_1434; // @[NV_NVDLA_CSC_wl.scala 499:46:@17016.4]
  wire [53:0] _GEN_559; // @[NV_NVDLA_CSC_wl.scala 499:46:@17017.4]
  wire [54:0] _T_1435; // @[NV_NVDLA_CSC_wl.scala 499:46:@17017.4]
  wire [54:0] _GEN_560; // @[NV_NVDLA_CSC_wl.scala 499:46:@17018.4]
  wire [55:0] _T_1436; // @[NV_NVDLA_CSC_wl.scala 499:46:@17018.4]
  wire [55:0] _GEN_561; // @[NV_NVDLA_CSC_wl.scala 499:46:@17019.4]
  wire [56:0] _T_1437; // @[NV_NVDLA_CSC_wl.scala 499:46:@17019.4]
  wire [56:0] _GEN_562; // @[NV_NVDLA_CSC_wl.scala 499:46:@17020.4]
  wire [57:0] _T_1438; // @[NV_NVDLA_CSC_wl.scala 499:46:@17020.4]
  wire [57:0] _GEN_563; // @[NV_NVDLA_CSC_wl.scala 499:46:@17021.4]
  wire [58:0] _T_1439; // @[NV_NVDLA_CSC_wl.scala 499:46:@17021.4]
  wire [58:0] _GEN_564; // @[NV_NVDLA_CSC_wl.scala 499:46:@17022.4]
  wire [59:0] _T_1440; // @[NV_NVDLA_CSC_wl.scala 499:46:@17022.4]
  wire [59:0] _GEN_565; // @[NV_NVDLA_CSC_wl.scala 499:46:@17023.4]
  wire [60:0] _T_1441; // @[NV_NVDLA_CSC_wl.scala 499:46:@17023.4]
  wire [60:0] _GEN_566; // @[NV_NVDLA_CSC_wl.scala 499:46:@17024.4]
  wire [61:0] _T_1442; // @[NV_NVDLA_CSC_wl.scala 499:46:@17024.4]
  wire [61:0] _GEN_567; // @[NV_NVDLA_CSC_wl.scala 499:46:@17025.4]
  wire [62:0] _T_1443; // @[NV_NVDLA_CSC_wl.scala 499:46:@17025.4]
  wire [62:0] _GEN_568; // @[NV_NVDLA_CSC_wl.scala 499:46:@17026.4]
  wire [63:0] _T_1444; // @[NV_NVDLA_CSC_wl.scala 499:46:@17026.4]
  reg [63:0] _T_1447; // @[NV_NVDLA_CSC_wl.scala 502:33:@17027.4]
  reg [63:0] _RAND_53;
  wire [190:0] _T_1453; // @[NV_NVDLA_CSC_wl.scala 505:57:@17029.4]
  wire [190:0] _T_1454; // @[NV_NVDLA_CSC_wl.scala 505:26:@17030.4]
  wire  _T_1456; // @[NV_NVDLA_CSC_wl.scala 508:45:@17031.4]
  wire [63:0] _T_1467; // @[NV_NVDLA_CSC_wl.scala 508:27:@17034.4]
  wire  _T_1469; // @[NV_NVDLA_CSC_wl.scala 509:45:@17035.4]
  wire [63:0] _T_1480; // @[NV_NVDLA_CSC_wl.scala 509:27:@17038.4]
  wire  _T_1482; // @[NV_NVDLA_CSC_wl.scala 510:45:@17039.4]
  wire [63:0] _T_1493; // @[NV_NVDLA_CSC_wl.scala 510:27:@17042.4]
  wire [5:0] _T_1494; // @[NV_NVDLA_CSC_wl.scala 514:50:@17043.4]
  wire [6:0] _T_1496; // @[Cat.scala 30:58:@17044.4]
  wire [63:0] _T_1497; // @[NV_NVDLA_CSC_wl.scala 515:39:@17045.4]
  wire [190:0] _GEN_569; // @[NV_NVDLA_CSC_wl.scala 515:61:@17046.4]
  wire [190:0] _T_1498; // @[NV_NVDLA_CSC_wl.scala 515:61:@17046.4]
  wire [63:0] _T_1500; // @[NV_NVDLA_CSC_wl.scala 516:62:@17048.4]
  wire [190:0] _GEN_570; // @[NV_NVDLA_CSC_wl.scala 516:83:@17049.4]
  wire [190:0] _T_1501; // @[NV_NVDLA_CSC_wl.scala 516:83:@17049.4]
  wire [190:0] _GEN_571; // @[NV_NVDLA_CSC_wl.scala 516:100:@17050.4]
  wire [190:0] _T_1502; // @[NV_NVDLA_CSC_wl.scala 516:100:@17050.4]
  wire [63:0] _T_1504; // @[NV_NVDLA_CSC_wl.scala 517:62:@17052.4]
  wire [190:0] _GEN_572; // @[NV_NVDLA_CSC_wl.scala 517:83:@17053.4]
  wire [190:0] _T_1505; // @[NV_NVDLA_CSC_wl.scala 517:83:@17053.4]
  wire [190:0] _GEN_573; // @[NV_NVDLA_CSC_wl.scala 517:100:@17054.4]
  wire [190:0] _T_1506; // @[NV_NVDLA_CSC_wl.scala 517:100:@17054.4]
  wire [63:0] _T_1508; // @[NV_NVDLA_CSC_wl.scala 518:62:@17056.4]
  wire [190:0] _GEN_574; // @[NV_NVDLA_CSC_wl.scala 518:83:@17057.4]
  wire [190:0] _T_1509; // @[NV_NVDLA_CSC_wl.scala 518:83:@17057.4]
  wire [190:0] _GEN_575; // @[NV_NVDLA_CSC_wl.scala 518:100:@17058.4]
  wire [190:0] _T_1510; // @[NV_NVDLA_CSC_wl.scala 518:100:@17058.4]
  wire  _T_1517; // @[NV_NVDLA_CSC_wl.scala 523:41:@17060.4]
  wire  _T_1519; // @[NV_NVDLA_CSC_wl.scala 524:41:@17061.4]
  wire [31:0] _T_1520; // @[NV_NVDLA_CSC_wl.scala 524:82:@17062.4]
  wire [31:0] _T_1521; // @[NV_NVDLA_CSC_wl.scala 524:122:@17063.4]
  wire [63:0] _T_1522; // @[Cat.scala 30:58:@17064.4]
  wire [15:0] _T_1523; // @[NV_NVDLA_CSC_wl.scala 525:44:@17065.4]
  wire [15:0] _T_1524; // @[NV_NVDLA_CSC_wl.scala 525:84:@17066.4]
  wire [15:0] _T_1525; // @[NV_NVDLA_CSC_wl.scala 525:124:@17067.4]
  wire [15:0] _T_1526; // @[NV_NVDLA_CSC_wl.scala 525:164:@17068.4]
  wire [63:0] _T_1529; // @[Cat.scala 30:58:@17071.4]
  wire [63:0] _T_1530; // @[NV_NVDLA_CSC_wl.scala 524:28:@17072.4]
  wire [190:0] _T_1531; // @[NV_NVDLA_CSC_wl.scala 523:28:@17073.4]
  wire [190:0] _T_1532; // @[NV_NVDLA_CSC_wl.scala 522:28:@17074.4]
  wire [190:0] _GEN_576; // @[NV_NVDLA_CSC_wl.scala 528:61:@17075.4]
  wire  _T_1533; // @[NV_NVDLA_CSC_wl.scala 528:61:@17075.4]
  wire  _T_1534; // @[NV_NVDLA_CSC_wl.scala 528:44:@17076.4]
  reg [7:0] _T_1537; // @[NV_NVDLA_CSC_wl.scala 531:30:@17077.4]
  reg [31:0] _RAND_54;
  reg [7:0] _T_1540; // @[NV_NVDLA_CSC_wl.scala 532:35:@17078.4]
  reg [31:0] _RAND_55;
  wire [63:0] _GEN_577; // @[NV_NVDLA_CSC_wl.scala 534:57:@17079.4]
  wire  _T_1541; // @[NV_NVDLA_CSC_wl.scala 534:57:@17079.4]
  wire  _T_1542; // @[NV_NVDLA_CSC_wl.scala 534:42:@17080.4]
  wire  _T_1543; // @[NV_NVDLA_CSC_wl.scala 536:31:@17081.4]
  wire [7:0] _T_1546; // @[NV_NVDLA_CSC_wl.scala 536:30:@17082.4]
  wire [8:0] _T_1547; // @[NV_NVDLA_CSC_wl.scala 538:39:@17083.4]
  wire [7:0] _T_1548; // @[NV_NVDLA_CSC_wl.scala 538:39:@17084.4]
  wire [63:0] _GEN_578; // @[NV_NVDLA_CSC_wl.scala 538:57:@17085.4]
  wire [64:0] _T_1549; // @[NV_NVDLA_CSC_wl.scala 538:57:@17085.4]
  wire [64:0] _T_1550; // @[NV_NVDLA_CSC_wl.scala 538:57:@17086.4]
  wire [63:0] _T_1551; // @[NV_NVDLA_CSC_wl.scala 538:57:@17087.4]
  wire  _T_1553; // @[NV_NVDLA_CSC_wl.scala 540:29:@17088.4]
  wire  _T_1554; // @[NV_NVDLA_CSC_wl.scala 540:47:@17089.4]
  wire [63:0] _T_1555; // @[NV_NVDLA_CSC_wl.scala 540:28:@17090.4]
  wire [63:0] _T_1556; // @[NV_NVDLA_CSC_wl.scala 539:28:@17091.4]
  wire  _T_1557; // @[NV_NVDLA_CSC_wl.scala 543:61:@17092.4]
  wire  _T_1558; // @[NV_NVDLA_CSC_wl.scala 543:81:@17093.4]
  wire  _T_1559; // @[NV_NVDLA_CSC_wl.scala 543:40:@17094.4]
  wire  _T_1560; // @[NV_NVDLA_CSC_wl.scala 545:19:@17095.4]
  wire [63:0] _GEN_49; // @[NV_NVDLA_CSC_wl.scala 545:39:@17096.4]
  wire [63:0] _GEN_50; // @[NV_NVDLA_CSC_wl.scala 548:30:@17099.4]
  reg [12:0] _T_1563; // @[NV_NVDLA_CSC_wl.scala 553:30:@17102.4]
  reg [31:0] _RAND_56;
  reg [12:0] _T_1566; // @[NV_NVDLA_CSC_wl.scala 554:35:@17103.4]
  reg [31:0] _RAND_57;
  wire [13:0] _T_1568; // @[NV_NVDLA_CSC_wl.scala 556:39:@17104.4]
  wire [12:0] _T_1569; // @[NV_NVDLA_CSC_wl.scala 556:39:@17105.4]
  wire [13:0] _GEN_579; // @[NV_NVDLA_CSC_wl.scala 557:48:@17108.4]
  wire  _T_1576; // @[NV_NVDLA_CSC_wl.scala 557:48:@17108.4]
  wire [12:0] _T_1582; // @[NV_NVDLA_CSC_wl.scala 558:35:@17110.4]
  wire [12:0] _T_1583; // @[NV_NVDLA_CSC_wl.scala 560:53:@17111.4]
  wire [12:0] _T_1586; // @[NV_NVDLA_CSC_wl.scala 562:28:@17114.4]
  wire [12:0] _T_1587; // @[NV_NVDLA_CSC_wl.scala 561:28:@17115.4]
  wire [12:0] _T_1588; // @[NV_NVDLA_CSC_wl.scala 560:28:@17116.4]
  wire  _T_1589; // @[NV_NVDLA_CSC_wl.scala 566:40:@17117.4]
  wire  _T_1590; // @[NV_NVDLA_CSC_wl.scala 566:76:@17118.4]
  wire  _T_1591; // @[NV_NVDLA_CSC_wl.scala 566:55:@17119.4]
  wire  _T_1592; // @[NV_NVDLA_CSC_wl.scala 567:66:@17120.4]
  wire  _T_1593; // @[NV_NVDLA_CSC_wl.scala 567:86:@17121.4]
  wire  _T_1594; // @[NV_NVDLA_CSC_wl.scala 567:45:@17122.4]
  wire [13:0] _T_1600; // @[Cat.scala 30:58:@17124.4]
  wire [13:0] _GEN_580; // @[NV_NVDLA_CSC_wl.scala 568:39:@17125.4]
  wire [14:0] _T_1601; // @[NV_NVDLA_CSC_wl.scala 568:39:@17125.4]
  wire [13:0] _T_1602; // @[NV_NVDLA_CSC_wl.scala 568:39:@17126.4]
  wire [12:0] _GEN_51; // @[NV_NVDLA_CSC_wl.scala 570:29:@17127.4]
  wire [12:0] _GEN_52; // @[NV_NVDLA_CSC_wl.scala 573:34:@17130.4]
  reg  _T_1605; // @[NV_NVDLA_CSC_wl.scala 578:33:@17133.4]
  reg [31:0] _RAND_58;
  reg [14:0] _T_1608; // @[NV_NVDLA_CSC_wl.scala 579:29:@17134.4]
  reg [31:0] _RAND_59;
  wire  _T_1609; // @[NV_NVDLA_CSC_wl.scala 581:42:@17135.4]
  wire  _T_1612; // @[NV_NVDLA_CSC_wl.scala 581:76:@17136.4]
  wire  _T_1613; // @[NV_NVDLA_CSC_wl.scala 581:31:@17137.4]
  wire [15:0] _T_1615; // @[NV_NVDLA_CSC_wl.scala 582:37:@17138.4]
  wire [14:0] _T_1616; // @[NV_NVDLA_CSC_wl.scala 582:37:@17139.4]
  wire [14:0] _T_1619; // @[NV_NVDLA_CSC_wl.scala 583:84:@17140.4]
  wire [14:0] _T_1620; // @[NV_NVDLA_CSC_wl.scala 583:27:@17141.4]
  wire  _T_1621; // @[NV_NVDLA_CSC_wl.scala 584:59:@17142.4]
  wire  _T_1622; // @[NV_NVDLA_CSC_wl.scala 584:38:@17143.4]
  wire  _T_1623; // @[NV_NVDLA_CSC_wl.scala 584:82:@17144.4]
  wire  _T_1624; // @[NV_NVDLA_CSC_wl.scala 584:98:@17145.4]
  wire  _T_1625; // @[NV_NVDLA_CSC_wl.scala 584:79:@17146.4]
  wire  _T_1627; // @[NV_NVDLA_CSC_wl.scala 585:45:@17148.4]
  wire [14:0] _T_1628; // @[NV_NVDLA_CSC_wl.scala 585:29:@17149.4]
  wire [14:0] _GEN_53; // @[NV_NVDLA_CSC_wl.scala 588:28:@17151.4]
  reg  _T_1631; // @[NV_NVDLA_CSC_wl.scala 593:38:@17154.4]
  reg [31:0] _RAND_60;
  reg [12:0] _T_1634; // @[NV_NVDLA_CSC_wl.scala 594:40:@17155.4]
  reg [31:0] _RAND_61;
  reg  _T_1637; // @[NV_NVDLA_CSC_wl.scala 596:39:@17156.4]
  reg [31:0] _RAND_62;
  reg  _T_1640; // @[NV_NVDLA_CSC_wl.scala 597:39:@17157.4]
  reg [31:0] _RAND_63;
  reg  _T_1643; // @[NV_NVDLA_CSC_wl.scala 598:40:@17158.4]
  reg [31:0] _RAND_64;
  reg  _T_1646; // @[NV_NVDLA_CSC_wl.scala 599:38:@17159.4]
  reg [31:0] _RAND_65;
  reg  _T_1649; // @[NV_NVDLA_CSC_wl.scala 600:32:@17160.4]
  reg [31:0] _RAND_66;
  reg [7:0] _T_1652; // @[NV_NVDLA_CSC_wl.scala 601:34:@17161.4]
  reg [31:0] _RAND_67;
  reg  _T_1655; // @[NV_NVDLA_CSC_wl.scala 603:36:@17162.4]
  reg [31:0] _RAND_68;
  reg [8:0] _T_1658; // @[NV_NVDLA_CSC_wl.scala 604:44:@17163.4]
  reg [31:0] _RAND_69;
  reg [14:0] _T_1661; // @[NV_NVDLA_CSC_wl.scala 605:43:@17164.4]
  reg [31:0] _RAND_70;
  wire [13:0] _GEN_54; // @[NV_NVDLA_CSC_wl.scala 609:23:@17166.4]
  wire  _GEN_55; // @[NV_NVDLA_CSC_wl.scala 613:28:@17170.4]
  wire  _GEN_56; // @[NV_NVDLA_CSC_wl.scala 613:28:@17170.4]
  wire  _GEN_57; // @[NV_NVDLA_CSC_wl.scala 613:28:@17170.4]
  wire  _GEN_58; // @[NV_NVDLA_CSC_wl.scala 613:28:@17170.4]
  wire [63:0] _GEN_59; // @[NV_NVDLA_CSC_wl.scala 613:28:@17170.4]
  wire [190:0] _GEN_60; // @[NV_NVDLA_CSC_wl.scala 621:39:@17178.4]
  wire [8:0] _GEN_61; // @[NV_NVDLA_CSC_wl.scala 625:28:@17182.4]
  wire  _T_1663; // @[NV_NVDLA_CSC_wl.scala 628:28:@17185.4]
  wire [14:0] _GEN_62; // @[NV_NVDLA_CSC_wl.scala 628:41:@17186.4]
  wire [35:0] _T_1672; // @[Cat.scala 30:58:@17199.4]
  reg  _T_1677; // @[NV_NVDLA_CSC_wl.scala 654:76:@17201.4]
  reg [31:0] _RAND_71;
  reg  _T_1680; // @[NV_NVDLA_CSC_wl.scala 654:76:@17202.4]
  reg [31:0] _RAND_72;
  reg  _T_1683; // @[NV_NVDLA_CSC_wl.scala 654:76:@17203.4]
  reg [31:0] _RAND_73;
  reg  _T_1686; // @[NV_NVDLA_CSC_wl.scala 654:76:@17204.4]
  reg [31:0] _RAND_74;
  reg  _T_1689; // @[NV_NVDLA_CSC_wl.scala 654:76:@17205.4]
  reg [31:0] _RAND_75;
  reg [35:0] _T_1697; // @[NV_NVDLA_CSC_wl.scala 656:75:@17208.4]
  reg [63:0] _RAND_76;
  reg [35:0] _T_1700; // @[NV_NVDLA_CSC_wl.scala 656:75:@17209.4]
  reg [63:0] _RAND_77;
  reg [35:0] _T_1703; // @[NV_NVDLA_CSC_wl.scala 656:75:@17210.4]
  reg [63:0] _RAND_78;
  reg [35:0] _T_1706; // @[NV_NVDLA_CSC_wl.scala 656:75:@17211.4]
  reg [63:0] _RAND_79;
  reg [35:0] _T_1709; // @[NV_NVDLA_CSC_wl.scala 656:75:@17212.4]
  reg [63:0] _RAND_80;
  reg  _T_1717; // @[NV_NVDLA_CSC_wl.scala 658:74:@17215.4]
  reg [31:0] _RAND_81;
  reg  _T_1720; // @[NV_NVDLA_CSC_wl.scala 658:74:@17216.4]
  reg [31:0] _RAND_82;
  reg  _T_1723; // @[NV_NVDLA_CSC_wl.scala 658:74:@17217.4]
  reg [31:0] _RAND_83;
  reg  _T_1726; // @[NV_NVDLA_CSC_wl.scala 658:74:@17218.4]
  reg [31:0] _RAND_84;
  reg  _T_1729; // @[NV_NVDLA_CSC_wl.scala 658:74:@17219.4]
  reg [31:0] _RAND_85;
  reg  _T_1732; // @[NV_NVDLA_CSC_wl.scala 658:74:@17220.4]
  reg [31:0] _RAND_86;
  reg [63:0] _T_1737; // @[NV_NVDLA_CSC_wl.scala 660:75:@17222.4]
  reg [63:0] _RAND_87;
  reg [63:0] _T_1740; // @[NV_NVDLA_CSC_wl.scala 660:75:@17223.4]
  reg [63:0] _RAND_88;
  reg [63:0] _T_1743; // @[NV_NVDLA_CSC_wl.scala 660:75:@17224.4]
  reg [63:0] _RAND_89;
  reg [63:0] _T_1746; // @[NV_NVDLA_CSC_wl.scala 660:75:@17225.4]
  reg [63:0] _RAND_90;
  reg [63:0] _T_1749; // @[NV_NVDLA_CSC_wl.scala 660:75:@17226.4]
  reg [63:0] _RAND_91;
  reg [63:0] _T_1752; // @[NV_NVDLA_CSC_wl.scala 660:75:@17227.4]
  reg [63:0] _RAND_92;
  wire [35:0] _GEN_63; // @[NV_NVDLA_CSC_wl.scala 669:36:@17233.4]
  wire [63:0] _GEN_64; // @[NV_NVDLA_CSC_wl.scala 673:34:@17237.4]
  wire [35:0] _GEN_65; // @[NV_NVDLA_CSC_wl.scala 669:36:@17241.4]
  wire [63:0] _GEN_66; // @[NV_NVDLA_CSC_wl.scala 673:34:@17245.4]
  wire [35:0] _GEN_67; // @[NV_NVDLA_CSC_wl.scala 669:36:@17249.4]
  wire [63:0] _GEN_68; // @[NV_NVDLA_CSC_wl.scala 673:34:@17253.4]
  wire [35:0] _GEN_69; // @[NV_NVDLA_CSC_wl.scala 669:36:@17257.4]
  wire [63:0] _GEN_70; // @[NV_NVDLA_CSC_wl.scala 673:34:@17261.4]
  wire [35:0] _GEN_71; // @[NV_NVDLA_CSC_wl.scala 669:36:@17265.4]
  wire [63:0] _GEN_72; // @[NV_NVDLA_CSC_wl.scala 673:34:@17269.4]
  wire [35:0] _GEN_73; // @[NV_NVDLA_CSC_wl.scala 669:36:@17273.4]
  wire [63:0] _GEN_74; // @[NV_NVDLA_CSC_wl.scala 673:34:@17277.4]
  wire [7:0] _T_1753; // @[NV_NVDLA_CSC_wl.scala 687:38:@17281.4]
  wire  _T_1756; // @[NV_NVDLA_CSC_wl.scala 690:44:@17286.4]
  wire  _T_1757; // @[NV_NVDLA_CSC_wl.scala 691:45:@17287.4]
  wire  _T_1758; // @[NV_NVDLA_CSC_wl.scala 692:43:@17288.4]
  reg [6:0] _T_1762; // @[NV_NVDLA_CSC_wl.scala 699:37:@17291.4]
  reg [31:0] _RAND_93;
  reg [6:0] _T_1765; // @[NV_NVDLA_CSC_wl.scala 700:42:@17292.4]
  reg [31:0] _RAND_94;
  wire [7:0] _T_1768; // @[NV_NVDLA_CSC_wl.scala 702:37:@17293.4]
  wire  _T_1770; // @[NV_NVDLA_CSC_wl.scala 704:55:@17294.4]
  wire  _T_1771; // @[NV_NVDLA_CSC_wl.scala 704:53:@17295.4]
  wire [8:0] _T_1773; // @[Cat.scala 30:58:@17296.4]
  wire [7:0] _GEN_581; // @[NV_NVDLA_CSC_wl.scala 704:141:@17297.4]
  wire [8:0] _T_1774; // @[NV_NVDLA_CSC_wl.scala 704:141:@17297.4]
  wire [7:0] _T_1775; // @[NV_NVDLA_CSC_wl.scala 704:141:@17298.4]
  wire [8:0] _T_1776; // @[NV_NVDLA_CSC_wl.scala 704:166:@17299.4]
  wire [8:0] _T_1777; // @[NV_NVDLA_CSC_wl.scala 704:166:@17300.4]
  wire [7:0] _T_1778; // @[NV_NVDLA_CSC_wl.scala 704:166:@17301.4]
  wire [8:0] _T_1779; // @[NV_NVDLA_CSC_wl.scala 704:33:@17302.4]
  wire [8:0] _T_1780; // @[NV_NVDLA_CSC_wl.scala 703:35:@17303.4]
  wire [6:0] _T_1781; // @[NV_NVDLA_CSC_wl.scala 704:182:@17304.4]
  wire  _T_1782; // @[NV_NVDLA_CSC_wl.scala 705:42:@17305.4]
  wire  _T_1783; // @[NV_NVDLA_CSC_wl.scala 706:67:@17306.4]
  wire  _T_1784; // @[NV_NVDLA_CSC_wl.scala 706:47:@17307.4]
  wire [6:0] _GEN_75; // @[NV_NVDLA_CSC_wl.scala 708:32:@17308.4]
  wire [6:0] _GEN_76; // @[NV_NVDLA_CSC_wl.scala 711:37:@17311.4]
  reg [511:0] _T_1786; // @[NV_NVDLA_CSC_wl.scala 716:29:@17314.4]
  reg [511:0] _RAND_95;
  reg [511:0] _T_1788; // @[NV_NVDLA_CSC_wl.scala 717:34:@17315.4]
  reg [511:0] _RAND_96;
  wire [8:0] _T_1790; // @[NV_NVDLA_CSC_wl.scala 719:40:@17317.4]
  wire [8:0] _T_1791; // @[NV_NVDLA_CSC_wl.scala 719:40:@17318.4]
  wire [7:0] _T_1792; // @[NV_NVDLA_CSC_wl.scala 719:40:@17319.4]
  wire [10:0] _T_1795; // @[Cat.scala 30:58:@17321.4]
  wire [511:0] _T_1796; // @[NV_NVDLA_CSC_wl.scala 720:82:@17322.4]
  wire  _T_1798; // @[NV_NVDLA_CSC_wl.scala 721:58:@17323.4]
  wire  _T_1799; // @[NV_NVDLA_CSC_wl.scala 721:38:@17324.4]
  wire [511:0] _T_1801; // @[NV_NVDLA_CSC_wl.scala 721:36:@17325.4]
  wire [10:0] _T_1803; // @[Cat.scala 30:58:@17326.4]
  wire [511:0] _T_1804; // @[NV_NVDLA_CSC_wl.scala 722:45:@17327.4]
  wire  _T_1809; // @[NV_NVDLA_CSC_wl.scala 725:98:@17330.4]
  wire  _T_1810; // @[NV_NVDLA_CSC_wl.scala 725:71:@17331.4]
  wire [511:0] _T_1811; // @[NV_NVDLA_CSC_wl.scala 726:31:@17332.4]
  wire [511:0] _T_1812; // @[NV_NVDLA_CSC_wl.scala 725:31:@17333.4]
  wire [511:0] _T_1813; // @[NV_NVDLA_CSC_wl.scala 724:31:@17334.4]
  wire  _T_1815; // @[NV_NVDLA_CSC_wl.scala 729:86:@17335.4]
  wire  _T_1816; // @[NV_NVDLA_CSC_wl.scala 729:62:@17336.4]
  wire  _T_1817; // @[NV_NVDLA_CSC_wl.scala 729:42:@17337.4]
  wire  _T_1821; // @[NV_NVDLA_CSC_wl.scala 730:86:@17340.4]
  wire  _T_1822; // @[NV_NVDLA_CSC_wl.scala 730:47:@17341.4]
  wire [9:0] _T_1825; // @[Cat.scala 30:58:@17343.4]
  wire [1534:0] _GEN_583; // @[NV_NVDLA_CSC_wl.scala 731:55:@17344.4]
  wire [1534:0] _T_1826; // @[NV_NVDLA_CSC_wl.scala 731:55:@17344.4]
  wire [1534:0] _T_1828; // @[NV_NVDLA_CSC_wl.scala 732:32:@17345.4]
  reg [7:0] _T_2095_0; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_97;
  reg [7:0] _T_2095_1; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_98;
  reg [7:0] _T_2095_2; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_99;
  reg [7:0] _T_2095_3; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_100;
  reg [7:0] _T_2095_4; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_101;
  reg [7:0] _T_2095_5; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_102;
  reg [7:0] _T_2095_6; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_103;
  reg [7:0] _T_2095_7; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_104;
  reg [7:0] _T_2095_8; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_105;
  reg [7:0] _T_2095_9; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_106;
  reg [7:0] _T_2095_10; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_107;
  reg [7:0] _T_2095_11; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_108;
  reg [7:0] _T_2095_12; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_109;
  reg [7:0] _T_2095_13; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_110;
  reg [7:0] _T_2095_14; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_111;
  reg [7:0] _T_2095_15; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_112;
  reg [7:0] _T_2095_16; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_113;
  reg [7:0] _T_2095_17; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_114;
  reg [7:0] _T_2095_18; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_115;
  reg [7:0] _T_2095_19; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_116;
  reg [7:0] _T_2095_20; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_117;
  reg [7:0] _T_2095_21; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_118;
  reg [7:0] _T_2095_22; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_119;
  reg [7:0] _T_2095_23; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_120;
  reg [7:0] _T_2095_24; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_121;
  reg [7:0] _T_2095_25; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_122;
  reg [7:0] _T_2095_26; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_123;
  reg [7:0] _T_2095_27; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_124;
  reg [7:0] _T_2095_28; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_125;
  reg [7:0] _T_2095_29; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_126;
  reg [7:0] _T_2095_30; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_127;
  reg [7:0] _T_2095_31; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_128;
  reg [7:0] _T_2095_32; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_129;
  reg [7:0] _T_2095_33; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_130;
  reg [7:0] _T_2095_34; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_131;
  reg [7:0] _T_2095_35; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_132;
  reg [7:0] _T_2095_36; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_133;
  reg [7:0] _T_2095_37; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_134;
  reg [7:0] _T_2095_38; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_135;
  reg [7:0] _T_2095_39; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_136;
  reg [7:0] _T_2095_40; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_137;
  reg [7:0] _T_2095_41; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_138;
  reg [7:0] _T_2095_42; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_139;
  reg [7:0] _T_2095_43; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_140;
  reg [7:0] _T_2095_44; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_141;
  reg [7:0] _T_2095_45; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_142;
  reg [7:0] _T_2095_46; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_143;
  reg [7:0] _T_2095_47; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_144;
  reg [7:0] _T_2095_48; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_145;
  reg [7:0] _T_2095_49; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_146;
  reg [7:0] _T_2095_50; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_147;
  reg [7:0] _T_2095_51; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_148;
  reg [7:0] _T_2095_52; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_149;
  reg [7:0] _T_2095_53; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_150;
  reg [7:0] _T_2095_54; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_151;
  reg [7:0] _T_2095_55; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_152;
  reg [7:0] _T_2095_56; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_153;
  reg [7:0] _T_2095_57; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_154;
  reg [7:0] _T_2095_58; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_155;
  reg [7:0] _T_2095_59; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_156;
  reg [7:0] _T_2095_60; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_157;
  reg [7:0] _T_2095_61; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_158;
  reg [7:0] _T_2095_62; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_159;
  reg [7:0] _T_2095_63; // @[NV_NVDLA_CSC_wl.scala 742:33:@17417.4]
  reg [31:0] _RAND_160;
  wire [1534:0] _GEN_584; // @[NV_NVDLA_CSC_wl.scala 744:42:@17418.4]
  wire [1534:0] _T_2292; // @[NV_NVDLA_CSC_wl.scala 744:42:@17418.4]
  wire [7:0] _T_2293; // @[NV_NVDLA_CSC_wl.scala 747:45:@17420.6]
  wire [7:0] _T_2294; // @[NV_NVDLA_CSC_wl.scala 747:45:@17422.6]
  wire [7:0] _T_2295; // @[NV_NVDLA_CSC_wl.scala 747:45:@17424.6]
  wire [7:0] _T_2296; // @[NV_NVDLA_CSC_wl.scala 747:45:@17426.6]
  wire [7:0] _T_2297; // @[NV_NVDLA_CSC_wl.scala 747:45:@17428.6]
  wire [7:0] _T_2298; // @[NV_NVDLA_CSC_wl.scala 747:45:@17430.6]
  wire [7:0] _T_2299; // @[NV_NVDLA_CSC_wl.scala 747:45:@17432.6]
  wire [7:0] _T_2300; // @[NV_NVDLA_CSC_wl.scala 747:45:@17434.6]
  wire [7:0] _T_2301; // @[NV_NVDLA_CSC_wl.scala 747:45:@17436.6]
  wire [7:0] _T_2302; // @[NV_NVDLA_CSC_wl.scala 747:45:@17438.6]
  wire [7:0] _T_2303; // @[NV_NVDLA_CSC_wl.scala 747:45:@17440.6]
  wire [7:0] _T_2304; // @[NV_NVDLA_CSC_wl.scala 747:45:@17442.6]
  wire [7:0] _T_2305; // @[NV_NVDLA_CSC_wl.scala 747:45:@17444.6]
  wire [7:0] _T_2306; // @[NV_NVDLA_CSC_wl.scala 747:45:@17446.6]
  wire [7:0] _T_2307; // @[NV_NVDLA_CSC_wl.scala 747:45:@17448.6]
  wire [7:0] _T_2308; // @[NV_NVDLA_CSC_wl.scala 747:45:@17450.6]
  wire [7:0] _T_2309; // @[NV_NVDLA_CSC_wl.scala 747:45:@17452.6]
  wire [7:0] _T_2310; // @[NV_NVDLA_CSC_wl.scala 747:45:@17454.6]
  wire [7:0] _T_2311; // @[NV_NVDLA_CSC_wl.scala 747:45:@17456.6]
  wire [7:0] _T_2312; // @[NV_NVDLA_CSC_wl.scala 747:45:@17458.6]
  wire [7:0] _T_2313; // @[NV_NVDLA_CSC_wl.scala 747:45:@17460.6]
  wire [7:0] _T_2314; // @[NV_NVDLA_CSC_wl.scala 747:45:@17462.6]
  wire [7:0] _T_2315; // @[NV_NVDLA_CSC_wl.scala 747:45:@17464.6]
  wire [7:0] _T_2316; // @[NV_NVDLA_CSC_wl.scala 747:45:@17466.6]
  wire [7:0] _T_2317; // @[NV_NVDLA_CSC_wl.scala 747:45:@17468.6]
  wire [7:0] _T_2318; // @[NV_NVDLA_CSC_wl.scala 747:45:@17470.6]
  wire [7:0] _T_2319; // @[NV_NVDLA_CSC_wl.scala 747:45:@17472.6]
  wire [7:0] _T_2320; // @[NV_NVDLA_CSC_wl.scala 747:45:@17474.6]
  wire [7:0] _T_2321; // @[NV_NVDLA_CSC_wl.scala 747:45:@17476.6]
  wire [7:0] _T_2322; // @[NV_NVDLA_CSC_wl.scala 747:45:@17478.6]
  wire [7:0] _T_2323; // @[NV_NVDLA_CSC_wl.scala 747:45:@17480.6]
  wire [7:0] _T_2324; // @[NV_NVDLA_CSC_wl.scala 747:45:@17482.6]
  wire [7:0] _T_2325; // @[NV_NVDLA_CSC_wl.scala 747:45:@17484.6]
  wire [7:0] _T_2326; // @[NV_NVDLA_CSC_wl.scala 747:45:@17486.6]
  wire [7:0] _T_2327; // @[NV_NVDLA_CSC_wl.scala 747:45:@17488.6]
  wire [7:0] _T_2328; // @[NV_NVDLA_CSC_wl.scala 747:45:@17490.6]
  wire [7:0] _T_2329; // @[NV_NVDLA_CSC_wl.scala 747:45:@17492.6]
  wire [7:0] _T_2330; // @[NV_NVDLA_CSC_wl.scala 747:45:@17494.6]
  wire [7:0] _T_2331; // @[NV_NVDLA_CSC_wl.scala 747:45:@17496.6]
  wire [7:0] _T_2332; // @[NV_NVDLA_CSC_wl.scala 747:45:@17498.6]
  wire [7:0] _T_2333; // @[NV_NVDLA_CSC_wl.scala 747:45:@17500.6]
  wire [7:0] _T_2334; // @[NV_NVDLA_CSC_wl.scala 747:45:@17502.6]
  wire [7:0] _T_2335; // @[NV_NVDLA_CSC_wl.scala 747:45:@17504.6]
  wire [7:0] _T_2336; // @[NV_NVDLA_CSC_wl.scala 747:45:@17506.6]
  wire [7:0] _T_2337; // @[NV_NVDLA_CSC_wl.scala 747:45:@17508.6]
  wire [7:0] _T_2338; // @[NV_NVDLA_CSC_wl.scala 747:45:@17510.6]
  wire [7:0] _T_2339; // @[NV_NVDLA_CSC_wl.scala 747:45:@17512.6]
  wire [7:0] _T_2340; // @[NV_NVDLA_CSC_wl.scala 747:45:@17514.6]
  wire [7:0] _T_2341; // @[NV_NVDLA_CSC_wl.scala 747:45:@17516.6]
  wire [7:0] _T_2342; // @[NV_NVDLA_CSC_wl.scala 747:45:@17518.6]
  wire [7:0] _T_2343; // @[NV_NVDLA_CSC_wl.scala 747:45:@17520.6]
  wire [7:0] _T_2344; // @[NV_NVDLA_CSC_wl.scala 747:45:@17522.6]
  wire [7:0] _T_2345; // @[NV_NVDLA_CSC_wl.scala 747:45:@17524.6]
  wire [7:0] _T_2346; // @[NV_NVDLA_CSC_wl.scala 747:45:@17526.6]
  wire [7:0] _T_2347; // @[NV_NVDLA_CSC_wl.scala 747:45:@17528.6]
  wire [7:0] _T_2348; // @[NV_NVDLA_CSC_wl.scala 747:45:@17530.6]
  wire [7:0] _T_2349; // @[NV_NVDLA_CSC_wl.scala 747:45:@17532.6]
  wire [7:0] _T_2350; // @[NV_NVDLA_CSC_wl.scala 747:45:@17534.6]
  wire [7:0] _T_2351; // @[NV_NVDLA_CSC_wl.scala 747:45:@17536.6]
  wire [7:0] _T_2352; // @[NV_NVDLA_CSC_wl.scala 747:45:@17538.6]
  wire [7:0] _T_2353; // @[NV_NVDLA_CSC_wl.scala 747:45:@17540.6]
  wire [7:0] _T_2354; // @[NV_NVDLA_CSC_wl.scala 747:45:@17542.6]
  wire [7:0] _T_2355; // @[NV_NVDLA_CSC_wl.scala 747:45:@17544.6]
  wire [7:0] _T_2356; // @[NV_NVDLA_CSC_wl.scala 747:45:@17546.6]
  wire [7:0] _GEN_79; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_80; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_81; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_82; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_83; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_84; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_85; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_86; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_87; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_88; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_89; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_90; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_91; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_92; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_93; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_94; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_95; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_96; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_97; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_98; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_99; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_100; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_101; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_102; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_103; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_104; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_105; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_106; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_107; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_108; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_109; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_110; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_111; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_112; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_113; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_114; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_115; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_116; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_117; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_118; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_119; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_120; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_121; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_122; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_123; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_124; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_125; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_126; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_127; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_128; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_129; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_130; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_131; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_132; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_133; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_134; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_135; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_136; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_137; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_138; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_139; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_140; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_141; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  wire [7:0] _GEN_142; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  reg  _T_2359; // @[NV_NVDLA_CSC_wl.scala 753:41:@17549.4]
  reg [31:0] _RAND_161;
  reg [31:0] _T_2362; // @[NV_NVDLA_CSC_wl.scala 754:32:@17550.4]
  reg [31:0] _RAND_162;
  wire [30:0] _T_2364; // @[NV_NVDLA_CSC_wl.scala 757:41:@17551.4]
  wire  _T_2365; // @[NV_NVDLA_CSC_wl.scala 757:77:@17552.4]
  wire [31:0] _T_2366; // @[Cat.scala 30:58:@17553.4]
  wire [31:0] _T_2367; // @[NV_NVDLA_CSC_wl.scala 756:27:@17554.4]
  wire  _GEN_143; // @[NV_NVDLA_CSC_wl.scala 759:27:@17555.4]
  wire [31:0] _GEN_144; // @[NV_NVDLA_CSC_wl.scala 759:27:@17555.4]
  reg  _T_2472; // @[NV_NVDLA_CSC_wl.scala 767:39:@17656.4]
  reg [31:0] _RAND_163;
  reg  _T_2739_0; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_164;
  reg  _T_2739_1; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_165;
  reg  _T_2739_2; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_166;
  reg  _T_2739_3; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_167;
  reg  _T_2739_4; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_168;
  reg  _T_2739_5; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_169;
  reg  _T_2739_6; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_170;
  reg  _T_2739_7; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_171;
  reg  _T_2739_8; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_172;
  reg  _T_2739_9; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_173;
  reg  _T_2739_10; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_174;
  reg  _T_2739_11; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_175;
  reg  _T_2739_12; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_176;
  reg  _T_2739_13; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_177;
  reg  _T_2739_14; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_178;
  reg  _T_2739_15; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_179;
  reg  _T_2739_16; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_180;
  reg  _T_2739_17; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_181;
  reg  _T_2739_18; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_182;
  reg  _T_2739_19; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_183;
  reg  _T_2739_20; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_184;
  reg  _T_2739_21; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_185;
  reg  _T_2739_22; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_186;
  reg  _T_2739_23; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_187;
  reg  _T_2739_24; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_188;
  reg  _T_2739_25; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_189;
  reg  _T_2739_26; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_190;
  reg  _T_2739_27; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_191;
  reg  _T_2739_28; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_192;
  reg  _T_2739_29; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_193;
  reg  _T_2739_30; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_194;
  reg  _T_2739_31; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_195;
  reg  _T_2739_32; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_196;
  reg  _T_2739_33; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_197;
  reg  _T_2739_34; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_198;
  reg  _T_2739_35; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_199;
  reg  _T_2739_36; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_200;
  reg  _T_2739_37; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_201;
  reg  _T_2739_38; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_202;
  reg  _T_2739_39; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_203;
  reg  _T_2739_40; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_204;
  reg  _T_2739_41; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_205;
  reg  _T_2739_42; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_206;
  reg  _T_2739_43; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_207;
  reg  _T_2739_44; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_208;
  reg  _T_2739_45; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_209;
  reg  _T_2739_46; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_210;
  reg  _T_2739_47; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_211;
  reg  _T_2739_48; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_212;
  reg  _T_2739_49; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_213;
  reg  _T_2739_50; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_214;
  reg  _T_2739_51; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_215;
  reg  _T_2739_52; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_216;
  reg  _T_2739_53; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_217;
  reg  _T_2739_54; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_218;
  reg  _T_2739_55; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_219;
  reg  _T_2739_56; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_220;
  reg  _T_2739_57; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_221;
  reg  _T_2739_58; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_222;
  reg  _T_2739_59; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_223;
  reg  _T_2739_60; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_224;
  reg  _T_2739_61; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_225;
  reg  _T_2739_62; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_226;
  reg  _T_2739_63; // @[NV_NVDLA_CSC_wl.scala 768:33:@17722.4]
  reg [31:0] _RAND_227;
  reg [9:0] _T_2938; // @[NV_NVDLA_CSC_wl.scala 769:36:@17723.4]
  reg [31:0] _RAND_228;
  wire  _T_2939; // @[NV_NVDLA_CSC_wl.scala 773:86:@17726.6]
  wire  _T_2940; // @[NV_NVDLA_CSC_wl.scala 773:86:@17727.6]
  wire  _T_2941; // @[NV_NVDLA_CSC_wl.scala 773:86:@17728.6]
  wire  _T_2942; // @[NV_NVDLA_CSC_wl.scala 773:86:@17729.6]
  wire  _T_2943; // @[NV_NVDLA_CSC_wl.scala 773:86:@17730.6]
  wire  _T_2944; // @[NV_NVDLA_CSC_wl.scala 773:86:@17731.6]
  wire  _T_2945; // @[NV_NVDLA_CSC_wl.scala 773:86:@17732.6]
  wire  _T_2946; // @[NV_NVDLA_CSC_wl.scala 773:86:@17733.6]
  wire  _T_2947; // @[NV_NVDLA_CSC_wl.scala 773:86:@17734.6]
  wire  _T_2948; // @[NV_NVDLA_CSC_wl.scala 773:86:@17735.6]
  wire  _T_2949; // @[NV_NVDLA_CSC_wl.scala 773:86:@17736.6]
  wire  _T_2950; // @[NV_NVDLA_CSC_wl.scala 773:86:@17737.6]
  wire  _T_2951; // @[NV_NVDLA_CSC_wl.scala 773:86:@17738.6]
  wire  _T_2952; // @[NV_NVDLA_CSC_wl.scala 773:86:@17739.6]
  wire  _T_2953; // @[NV_NVDLA_CSC_wl.scala 773:86:@17740.6]
  wire  _T_2954; // @[NV_NVDLA_CSC_wl.scala 773:86:@17741.6]
  wire  _T_2955; // @[NV_NVDLA_CSC_wl.scala 773:86:@17742.6]
  wire  _T_2956; // @[NV_NVDLA_CSC_wl.scala 773:86:@17743.6]
  wire  _T_2957; // @[NV_NVDLA_CSC_wl.scala 773:86:@17744.6]
  wire  _T_2958; // @[NV_NVDLA_CSC_wl.scala 773:86:@17745.6]
  wire  _T_2959; // @[NV_NVDLA_CSC_wl.scala 773:86:@17746.6]
  wire  _T_2960; // @[NV_NVDLA_CSC_wl.scala 773:86:@17747.6]
  wire  _T_2961; // @[NV_NVDLA_CSC_wl.scala 773:86:@17748.6]
  wire  _T_2962; // @[NV_NVDLA_CSC_wl.scala 773:86:@17749.6]
  wire  _T_2963; // @[NV_NVDLA_CSC_wl.scala 773:86:@17750.6]
  wire  _T_2964; // @[NV_NVDLA_CSC_wl.scala 773:86:@17751.6]
  wire  _T_2965; // @[NV_NVDLA_CSC_wl.scala 773:86:@17752.6]
  wire  _T_2966; // @[NV_NVDLA_CSC_wl.scala 773:86:@17753.6]
  wire  _T_2967; // @[NV_NVDLA_CSC_wl.scala 773:86:@17754.6]
  wire  _T_2968; // @[NV_NVDLA_CSC_wl.scala 773:86:@17755.6]
  wire  _T_2969; // @[NV_NVDLA_CSC_wl.scala 773:86:@17756.6]
  wire  _T_2970; // @[NV_NVDLA_CSC_wl.scala 773:86:@17757.6]
  wire  _T_2971; // @[NV_NVDLA_CSC_wl.scala 773:86:@17758.6]
  wire  _T_2972; // @[NV_NVDLA_CSC_wl.scala 773:86:@17759.6]
  wire  _T_2973; // @[NV_NVDLA_CSC_wl.scala 773:86:@17760.6]
  wire  _T_2974; // @[NV_NVDLA_CSC_wl.scala 773:86:@17761.6]
  wire  _T_2975; // @[NV_NVDLA_CSC_wl.scala 773:86:@17762.6]
  wire  _T_2976; // @[NV_NVDLA_CSC_wl.scala 773:86:@17763.6]
  wire  _T_2977; // @[NV_NVDLA_CSC_wl.scala 773:86:@17764.6]
  wire  _T_2978; // @[NV_NVDLA_CSC_wl.scala 773:86:@17765.6]
  wire  _T_2979; // @[NV_NVDLA_CSC_wl.scala 773:86:@17766.6]
  wire  _T_2980; // @[NV_NVDLA_CSC_wl.scala 773:86:@17767.6]
  wire  _T_2981; // @[NV_NVDLA_CSC_wl.scala 773:86:@17768.6]
  wire  _T_2982; // @[NV_NVDLA_CSC_wl.scala 773:86:@17769.6]
  wire  _T_2983; // @[NV_NVDLA_CSC_wl.scala 773:86:@17770.6]
  wire  _T_2984; // @[NV_NVDLA_CSC_wl.scala 773:86:@17771.6]
  wire  _T_2985; // @[NV_NVDLA_CSC_wl.scala 773:86:@17772.6]
  wire  _T_2986; // @[NV_NVDLA_CSC_wl.scala 773:86:@17773.6]
  wire  _T_2987; // @[NV_NVDLA_CSC_wl.scala 773:86:@17774.6]
  wire  _T_2988; // @[NV_NVDLA_CSC_wl.scala 773:86:@17775.6]
  wire  _T_2989; // @[NV_NVDLA_CSC_wl.scala 773:86:@17776.6]
  wire  _T_2990; // @[NV_NVDLA_CSC_wl.scala 773:86:@17777.6]
  wire  _T_2991; // @[NV_NVDLA_CSC_wl.scala 773:86:@17778.6]
  wire  _T_2992; // @[NV_NVDLA_CSC_wl.scala 773:86:@17779.6]
  wire  _T_2993; // @[NV_NVDLA_CSC_wl.scala 773:86:@17780.6]
  wire  _T_2994; // @[NV_NVDLA_CSC_wl.scala 773:86:@17781.6]
  wire  _T_2995; // @[NV_NVDLA_CSC_wl.scala 773:86:@17782.6]
  wire  _T_2996; // @[NV_NVDLA_CSC_wl.scala 773:86:@17783.6]
  wire  _T_2997; // @[NV_NVDLA_CSC_wl.scala 773:86:@17784.6]
  wire  _T_2998; // @[NV_NVDLA_CSC_wl.scala 773:86:@17785.6]
  wire  _T_2999; // @[NV_NVDLA_CSC_wl.scala 773:86:@17786.6]
  wire  _T_3000; // @[NV_NVDLA_CSC_wl.scala 773:86:@17787.6]
  wire  _T_3001; // @[NV_NVDLA_CSC_wl.scala 773:86:@17788.6]
  wire  _T_3002; // @[NV_NVDLA_CSC_wl.scala 773:86:@17789.6]
  wire  _GEN_145; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_146; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_147; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_148; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_149; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_150; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_151; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_152; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_153; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_154; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_155; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_156; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_157; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_158; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_159; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_160; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_161; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_162; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_163; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_164; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_165; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_166; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_167; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_168; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_169; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_170; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_171; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_172; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_173; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_174; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_175; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_176; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_177; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_178; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_179; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_180; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_181; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_182; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_183; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_184; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_185; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_186; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_187; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_188; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_189; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_190; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_191; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_192; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_193; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_194; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_195; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_196; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_197; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_198; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_199; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_200; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_201; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_202; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_203; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_204; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_205; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_206; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_207; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire  _GEN_208; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  wire [9:0] _T_3076; // @[Bitwise.scala 72:12:@17921.4]
  wire  _T_3077; // @[Bitwise.scala 72:15:@18089.4]
  wire [15:0] _T_3080; // @[Bitwise.scala 72:12:@18090.4]
  wire [7:0] _T_3087; // @[NV_NVDLA_CSC_wl.scala 794:92:@18097.4]
  wire [15:0] _T_3095; // @[NV_NVDLA_CSC_wl.scala 794:92:@18105.4]
  wire [7:0] _T_3102; // @[NV_NVDLA_CSC_wl.scala 794:92:@18112.4]
  wire [31:0] _T_3111; // @[NV_NVDLA_CSC_wl.scala 794:92:@18121.4]
  wire [15:0] _T_3112; // @[NV_NVDLA_CSC_wl.scala 794:99:@18122.4]
  wire [15:0] _T_3113; // @[NV_NVDLA_CSC_wl.scala 794:71:@18123.4]
  wire [15:0] _T_3149; // @[NV_NVDLA_CSC_wl.scala 795:99:@18157.4]
  wire [15:0] _T_3150; // @[NV_NVDLA_CSC_wl.scala 795:71:@18158.4]
  wire  _T_3152; // @[NV_NVDLA_CSC_wl.scala 796:49:@18159.4]
  wire  _T_3154; // @[NV_NVDLA_CSC_wl.scala 797:49:@18160.4]
  reg  _T_3157; // @[NV_NVDLA_CSC_wl.scala 799:39:@18161.4]
  reg [31:0] _RAND_229;
  reg  _T_3160; // @[NV_NVDLA_CSC_wl.scala 800:39:@18162.4]
  reg [31:0] _RAND_230;
  reg  _T_3427_0; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_231;
  reg  _T_3427_1; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_232;
  reg  _T_3427_2; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_233;
  reg  _T_3427_3; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_234;
  reg  _T_3427_4; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_235;
  reg  _T_3427_5; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_236;
  reg  _T_3427_6; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_237;
  reg  _T_3427_7; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_238;
  reg  _T_3427_8; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_239;
  reg  _T_3427_9; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_240;
  reg  _T_3427_10; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_241;
  reg  _T_3427_11; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_242;
  reg  _T_3427_12; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_243;
  reg  _T_3427_13; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_244;
  reg  _T_3427_14; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_245;
  reg  _T_3427_15; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_246;
  reg  _T_3427_16; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_247;
  reg  _T_3427_17; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_248;
  reg  _T_3427_18; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_249;
  reg  _T_3427_19; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_250;
  reg  _T_3427_20; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_251;
  reg  _T_3427_21; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_252;
  reg  _T_3427_22; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_253;
  reg  _T_3427_23; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_254;
  reg  _T_3427_24; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_255;
  reg  _T_3427_25; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_256;
  reg  _T_3427_26; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_257;
  reg  _T_3427_27; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_258;
  reg  _T_3427_28; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_259;
  reg  _T_3427_29; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_260;
  reg  _T_3427_30; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_261;
  reg  _T_3427_31; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_262;
  reg  _T_3427_32; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_263;
  reg  _T_3427_33; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_264;
  reg  _T_3427_34; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_265;
  reg  _T_3427_35; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_266;
  reg  _T_3427_36; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_267;
  reg  _T_3427_37; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_268;
  reg  _T_3427_38; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_269;
  reg  _T_3427_39; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_270;
  reg  _T_3427_40; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_271;
  reg  _T_3427_41; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_272;
  reg  _T_3427_42; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_273;
  reg  _T_3427_43; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_274;
  reg  _T_3427_44; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_275;
  reg  _T_3427_45; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_276;
  reg  _T_3427_46; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_277;
  reg  _T_3427_47; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_278;
  reg  _T_3427_48; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_279;
  reg  _T_3427_49; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_280;
  reg  _T_3427_50; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_281;
  reg  _T_3427_51; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_282;
  reg  _T_3427_52; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_283;
  reg  _T_3427_53; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_284;
  reg  _T_3427_54; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_285;
  reg  _T_3427_55; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_286;
  reg  _T_3427_56; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_287;
  reg  _T_3427_57; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_288;
  reg  _T_3427_58; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_289;
  reg  _T_3427_59; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_290;
  reg  _T_3427_60; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_291;
  reg  _T_3427_61; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_292;
  reg  _T_3427_62; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_293;
  reg  _T_3427_63; // @[NV_NVDLA_CSC_wl.scala 801:39:@18228.4]
  reg [31:0] _RAND_294;
  reg  _T_3890_0; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_295;
  reg  _T_3890_1; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_296;
  reg  _T_3890_2; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_297;
  reg  _T_3890_3; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_298;
  reg  _T_3890_4; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_299;
  reg  _T_3890_5; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_300;
  reg  _T_3890_6; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_301;
  reg  _T_3890_7; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_302;
  reg  _T_3890_8; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_303;
  reg  _T_3890_9; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_304;
  reg  _T_3890_10; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_305;
  reg  _T_3890_11; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_306;
  reg  _T_3890_12; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_307;
  reg  _T_3890_13; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_308;
  reg  _T_3890_14; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_309;
  reg  _T_3890_15; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_310;
  reg  _T_3890_16; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_311;
  reg  _T_3890_17; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_312;
  reg  _T_3890_18; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_313;
  reg  _T_3890_19; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_314;
  reg  _T_3890_20; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_315;
  reg  _T_3890_21; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_316;
  reg  _T_3890_22; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_317;
  reg  _T_3890_23; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_318;
  reg  _T_3890_24; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_319;
  reg  _T_3890_25; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_320;
  reg  _T_3890_26; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_321;
  reg  _T_3890_27; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_322;
  reg  _T_3890_28; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_323;
  reg  _T_3890_29; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_324;
  reg  _T_3890_30; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_325;
  reg  _T_3890_31; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_326;
  reg  _T_3890_32; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_327;
  reg  _T_3890_33; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_328;
  reg  _T_3890_34; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_329;
  reg  _T_3890_35; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_330;
  reg  _T_3890_36; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_331;
  reg  _T_3890_37; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_332;
  reg  _T_3890_38; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_333;
  reg  _T_3890_39; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_334;
  reg  _T_3890_40; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_335;
  reg  _T_3890_41; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_336;
  reg  _T_3890_42; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_337;
  reg  _T_3890_43; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_338;
  reg  _T_3890_44; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_339;
  reg  _T_3890_45; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_340;
  reg  _T_3890_46; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_341;
  reg  _T_3890_47; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_342;
  reg  _T_3890_48; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_343;
  reg  _T_3890_49; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_344;
  reg  _T_3890_50; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_345;
  reg  _T_3890_51; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_346;
  reg  _T_3890_52; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_347;
  reg  _T_3890_53; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_348;
  reg  _T_3890_54; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_349;
  reg  _T_3890_55; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_350;
  reg  _T_3890_56; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_351;
  reg  _T_3890_57; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_352;
  reg  _T_3890_58; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_353;
  reg  _T_3890_59; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_354;
  reg  _T_3890_60; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_355;
  reg  _T_3890_61; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_356;
  reg  _T_3890_62; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_357;
  reg  _T_3890_63; // @[NV_NVDLA_CSC_wl.scala 802:39:@18294.4]
  reg [31:0] _RAND_358;
  reg  _T_4161_0; // @[NV_NVDLA_CSC_wl.scala 803:38:@18312.4]
  reg [31:0] _RAND_359;
  reg  _T_4161_1; // @[NV_NVDLA_CSC_wl.scala 803:38:@18312.4]
  reg [31:0] _RAND_360;
  reg  _T_4161_2; // @[NV_NVDLA_CSC_wl.scala 803:38:@18312.4]
  reg [31:0] _RAND_361;
  reg  _T_4161_3; // @[NV_NVDLA_CSC_wl.scala 803:38:@18312.4]
  reg [31:0] _RAND_362;
  reg  _T_4161_4; // @[NV_NVDLA_CSC_wl.scala 803:38:@18312.4]
  reg [31:0] _RAND_363;
  reg  _T_4161_5; // @[NV_NVDLA_CSC_wl.scala 803:38:@18312.4]
  reg [31:0] _RAND_364;
  reg  _T_4161_6; // @[NV_NVDLA_CSC_wl.scala 803:38:@18312.4]
  reg [31:0] _RAND_365;
  reg  _T_4161_7; // @[NV_NVDLA_CSC_wl.scala 803:38:@18312.4]
  reg [31:0] _RAND_366;
  reg  _T_4161_8; // @[NV_NVDLA_CSC_wl.scala 803:38:@18312.4]
  reg [31:0] _RAND_367;
  reg  _T_4161_9; // @[NV_NVDLA_CSC_wl.scala 803:38:@18312.4]
  reg [31:0] _RAND_368;
  reg  _T_4161_10; // @[NV_NVDLA_CSC_wl.scala 803:38:@18312.4]
  reg [31:0] _RAND_369;
  reg  _T_4161_11; // @[NV_NVDLA_CSC_wl.scala 803:38:@18312.4]
  reg [31:0] _RAND_370;
  reg  _T_4161_12; // @[NV_NVDLA_CSC_wl.scala 803:38:@18312.4]
  reg [31:0] _RAND_371;
  reg  _T_4161_13; // @[NV_NVDLA_CSC_wl.scala 803:38:@18312.4]
  reg [31:0] _RAND_372;
  reg  _T_4161_14; // @[NV_NVDLA_CSC_wl.scala 803:38:@18312.4]
  reg [31:0] _RAND_373;
  reg  _T_4161_15; // @[NV_NVDLA_CSC_wl.scala 803:38:@18312.4]
  reg [31:0] _RAND_374;
  reg  _T_4288_0; // @[NV_NVDLA_CSC_wl.scala 804:38:@18330.4]
  reg [31:0] _RAND_375;
  reg  _T_4288_1; // @[NV_NVDLA_CSC_wl.scala 804:38:@18330.4]
  reg [31:0] _RAND_376;
  reg  _T_4288_2; // @[NV_NVDLA_CSC_wl.scala 804:38:@18330.4]
  reg [31:0] _RAND_377;
  reg  _T_4288_3; // @[NV_NVDLA_CSC_wl.scala 804:38:@18330.4]
  reg [31:0] _RAND_378;
  reg  _T_4288_4; // @[NV_NVDLA_CSC_wl.scala 804:38:@18330.4]
  reg [31:0] _RAND_379;
  reg  _T_4288_5; // @[NV_NVDLA_CSC_wl.scala 804:38:@18330.4]
  reg [31:0] _RAND_380;
  reg  _T_4288_6; // @[NV_NVDLA_CSC_wl.scala 804:38:@18330.4]
  reg [31:0] _RAND_381;
  reg  _T_4288_7; // @[NV_NVDLA_CSC_wl.scala 804:38:@18330.4]
  reg [31:0] _RAND_382;
  reg  _T_4288_8; // @[NV_NVDLA_CSC_wl.scala 804:38:@18330.4]
  reg [31:0] _RAND_383;
  reg  _T_4288_9; // @[NV_NVDLA_CSC_wl.scala 804:38:@18330.4]
  reg [31:0] _RAND_384;
  reg  _T_4288_10; // @[NV_NVDLA_CSC_wl.scala 804:38:@18330.4]
  reg [31:0] _RAND_385;
  reg  _T_4288_11; // @[NV_NVDLA_CSC_wl.scala 804:38:@18330.4]
  reg [31:0] _RAND_386;
  reg  _T_4288_12; // @[NV_NVDLA_CSC_wl.scala 804:38:@18330.4]
  reg [31:0] _RAND_387;
  reg  _T_4288_13; // @[NV_NVDLA_CSC_wl.scala 804:38:@18330.4]
  reg [31:0] _RAND_388;
  reg  _T_4288_14; // @[NV_NVDLA_CSC_wl.scala 804:38:@18330.4]
  reg [31:0] _RAND_389;
  reg  _T_4288_15; // @[NV_NVDLA_CSC_wl.scala 804:38:@18330.4]
  reg [31:0] _RAND_390;
  reg [7:0] _T_4344_0; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_391;
  reg [7:0] _T_4344_1; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_392;
  reg [7:0] _T_4344_2; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_393;
  reg [7:0] _T_4344_3; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_394;
  reg [7:0] _T_4344_4; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_395;
  reg [7:0] _T_4344_5; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_396;
  reg [7:0] _T_4344_6; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_397;
  reg [7:0] _T_4344_7; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_398;
  reg [7:0] _T_4344_8; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_399;
  reg [7:0] _T_4344_9; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_400;
  reg [7:0] _T_4344_10; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_401;
  reg [7:0] _T_4344_11; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_402;
  reg [7:0] _T_4344_12; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_403;
  reg [7:0] _T_4344_13; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_404;
  reg [7:0] _T_4344_14; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_405;
  reg [7:0] _T_4344_15; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_406;
  reg [7:0] _T_4344_16; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_407;
  reg [7:0] _T_4344_17; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_408;
  reg [7:0] _T_4344_18; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_409;
  reg [7:0] _T_4344_19; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_410;
  reg [7:0] _T_4344_20; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_411;
  reg [7:0] _T_4344_21; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_412;
  reg [7:0] _T_4344_22; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_413;
  reg [7:0] _T_4344_23; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_414;
  reg [7:0] _T_4344_24; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_415;
  reg [7:0] _T_4344_25; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_416;
  reg [7:0] _T_4344_26; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_417;
  reg [7:0] _T_4344_27; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_418;
  reg [7:0] _T_4344_28; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_419;
  reg [7:0] _T_4344_29; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_420;
  reg [7:0] _T_4344_30; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_421;
  reg [7:0] _T_4344_31; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_422;
  reg [7:0] _T_4344_32; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_423;
  reg [7:0] _T_4344_33; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_424;
  reg [7:0] _T_4344_34; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_425;
  reg [7:0] _T_4344_35; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_426;
  reg [7:0] _T_4344_36; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_427;
  reg [7:0] _T_4344_37; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_428;
  reg [7:0] _T_4344_38; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_429;
  reg [7:0] _T_4344_39; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_430;
  reg [7:0] _T_4344_40; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_431;
  reg [7:0] _T_4344_41; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_432;
  reg [7:0] _T_4344_42; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_433;
  reg [7:0] _T_4344_43; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_434;
  reg [7:0] _T_4344_44; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_435;
  reg [7:0] _T_4344_45; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_436;
  reg [7:0] _T_4344_46; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_437;
  reg [7:0] _T_4344_47; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_438;
  reg [7:0] _T_4344_48; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_439;
  reg [7:0] _T_4344_49; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_440;
  reg [7:0] _T_4344_50; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_441;
  reg [7:0] _T_4344_51; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_442;
  reg [7:0] _T_4344_52; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_443;
  reg [7:0] _T_4344_53; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_444;
  reg [7:0] _T_4344_54; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_445;
  reg [7:0] _T_4344_55; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_446;
  reg [7:0] _T_4344_56; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_447;
  reg [7:0] _T_4344_57; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_448;
  reg [7:0] _T_4344_58; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_449;
  reg [7:0] _T_4344_59; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_450;
  reg [7:0] _T_4344_60; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_451;
  reg [7:0] _T_4344_61; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_452;
  reg [7:0] _T_4344_62; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_453;
  reg [7:0] _T_4344_63; // @[NV_NVDLA_CSC_wl.scala 805:35:@18331.4]
  reg [31:0] _RAND_454;
  reg [7:0] _T_4414_0; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_455;
  reg [7:0] _T_4414_1; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_456;
  reg [7:0] _T_4414_2; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_457;
  reg [7:0] _T_4414_3; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_458;
  reg [7:0] _T_4414_4; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_459;
  reg [7:0] _T_4414_5; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_460;
  reg [7:0] _T_4414_6; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_461;
  reg [7:0] _T_4414_7; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_462;
  reg [7:0] _T_4414_8; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_463;
  reg [7:0] _T_4414_9; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_464;
  reg [7:0] _T_4414_10; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_465;
  reg [7:0] _T_4414_11; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_466;
  reg [7:0] _T_4414_12; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_467;
  reg [7:0] _T_4414_13; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_468;
  reg [7:0] _T_4414_14; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_469;
  reg [7:0] _T_4414_15; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_470;
  reg [7:0] _T_4414_16; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_471;
  reg [7:0] _T_4414_17; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_472;
  reg [7:0] _T_4414_18; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_473;
  reg [7:0] _T_4414_19; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_474;
  reg [7:0] _T_4414_20; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_475;
  reg [7:0] _T_4414_21; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_476;
  reg [7:0] _T_4414_22; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_477;
  reg [7:0] _T_4414_23; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_478;
  reg [7:0] _T_4414_24; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_479;
  reg [7:0] _T_4414_25; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_480;
  reg [7:0] _T_4414_26; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_481;
  reg [7:0] _T_4414_27; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_482;
  reg [7:0] _T_4414_28; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_483;
  reg [7:0] _T_4414_29; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_484;
  reg [7:0] _T_4414_30; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_485;
  reg [7:0] _T_4414_31; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_486;
  reg [7:0] _T_4414_32; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_487;
  reg [7:0] _T_4414_33; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_488;
  reg [7:0] _T_4414_34; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_489;
  reg [7:0] _T_4414_35; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_490;
  reg [7:0] _T_4414_36; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_491;
  reg [7:0] _T_4414_37; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_492;
  reg [7:0] _T_4414_38; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_493;
  reg [7:0] _T_4414_39; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_494;
  reg [7:0] _T_4414_40; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_495;
  reg [7:0] _T_4414_41; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_496;
  reg [7:0] _T_4414_42; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_497;
  reg [7:0] _T_4414_43; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_498;
  reg [7:0] _T_4414_44; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_499;
  reg [7:0] _T_4414_45; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_500;
  reg [7:0] _T_4414_46; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_501;
  reg [7:0] _T_4414_47; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_502;
  reg [7:0] _T_4414_48; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_503;
  reg [7:0] _T_4414_49; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_504;
  reg [7:0] _T_4414_50; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_505;
  reg [7:0] _T_4414_51; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_506;
  reg [7:0] _T_4414_52; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_507;
  reg [7:0] _T_4414_53; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_508;
  reg [7:0] _T_4414_54; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_509;
  reg [7:0] _T_4414_55; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_510;
  reg [7:0] _T_4414_56; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_511;
  reg [7:0] _T_4414_57; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_512;
  reg [7:0] _T_4414_58; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_513;
  reg [7:0] _T_4414_59; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_514;
  reg [7:0] _T_4414_60; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_515;
  reg [7:0] _T_4414_61; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_516;
  reg [7:0] _T_4414_62; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_517;
  reg [7:0] _T_4414_63; // @[NV_NVDLA_CSC_wl.scala 806:35:@18332.4]
  reg [31:0] _RAND_518;
  wire  _T_4481; // @[NV_NVDLA_CSC_wl.scala 807:91:@18333.4]
  wire  _T_4482; // @[NV_NVDLA_CSC_wl.scala 807:97:@18334.4]
  wire  _T_4483; // @[NV_NVDLA_CSC_wl.scala 807:91:@18335.4]
  wire  _T_4484; // @[NV_NVDLA_CSC_wl.scala 807:97:@18336.4]
  wire  _T_4485; // @[NV_NVDLA_CSC_wl.scala 807:91:@18337.4]
  wire  _T_4486; // @[NV_NVDLA_CSC_wl.scala 807:97:@18338.4]
  wire  _T_4487; // @[NV_NVDLA_CSC_wl.scala 807:91:@18339.4]
  wire  _T_4488; // @[NV_NVDLA_CSC_wl.scala 807:97:@18340.4]
  wire  _T_4489; // @[NV_NVDLA_CSC_wl.scala 807:91:@18341.4]
  wire  _T_4490; // @[NV_NVDLA_CSC_wl.scala 807:97:@18342.4]
  wire  _T_4491; // @[NV_NVDLA_CSC_wl.scala 807:91:@18343.4]
  wire  _T_4492; // @[NV_NVDLA_CSC_wl.scala 807:97:@18344.4]
  wire  _T_4493; // @[NV_NVDLA_CSC_wl.scala 807:91:@18345.4]
  wire  _T_4494; // @[NV_NVDLA_CSC_wl.scala 807:97:@18346.4]
  wire  _T_4495; // @[NV_NVDLA_CSC_wl.scala 807:91:@18347.4]
  wire  _T_4496; // @[NV_NVDLA_CSC_wl.scala 807:97:@18348.4]
  wire  _T_4497; // @[NV_NVDLA_CSC_wl.scala 807:91:@18349.4]
  wire  _T_4498; // @[NV_NVDLA_CSC_wl.scala 807:97:@18350.4]
  wire  _T_4499; // @[NV_NVDLA_CSC_wl.scala 807:91:@18351.4]
  wire  _T_4500; // @[NV_NVDLA_CSC_wl.scala 807:97:@18352.4]
  wire  _T_4501; // @[NV_NVDLA_CSC_wl.scala 807:91:@18353.4]
  wire  _T_4502; // @[NV_NVDLA_CSC_wl.scala 807:97:@18354.4]
  wire  _T_4503; // @[NV_NVDLA_CSC_wl.scala 807:91:@18355.4]
  wire  _T_4504; // @[NV_NVDLA_CSC_wl.scala 807:97:@18356.4]
  wire  _T_4505; // @[NV_NVDLA_CSC_wl.scala 807:91:@18357.4]
  wire  _T_4506; // @[NV_NVDLA_CSC_wl.scala 807:97:@18358.4]
  wire  _T_4507; // @[NV_NVDLA_CSC_wl.scala 807:91:@18359.4]
  wire  _T_4508; // @[NV_NVDLA_CSC_wl.scala 807:97:@18360.4]
  wire  _T_4509; // @[NV_NVDLA_CSC_wl.scala 807:91:@18361.4]
  wire  _T_4510; // @[NV_NVDLA_CSC_wl.scala 807:97:@18362.4]
  wire  _T_4511; // @[NV_NVDLA_CSC_wl.scala 807:91:@18363.4]
  wire  _T_4512; // @[NV_NVDLA_CSC_wl.scala 807:97:@18364.4]
  wire  _T_4513; // @[NV_NVDLA_CSC_wl.scala 807:91:@18365.4]
  wire  _T_4514; // @[NV_NVDLA_CSC_wl.scala 807:97:@18366.4]
  wire  _T_4515; // @[NV_NVDLA_CSC_wl.scala 807:91:@18367.4]
  wire  _T_4516; // @[NV_NVDLA_CSC_wl.scala 807:97:@18368.4]
  wire  _T_4517; // @[NV_NVDLA_CSC_wl.scala 807:91:@18369.4]
  wire  _T_4518; // @[NV_NVDLA_CSC_wl.scala 807:97:@18370.4]
  wire  _T_4519; // @[NV_NVDLA_CSC_wl.scala 807:91:@18371.4]
  wire  _T_4520; // @[NV_NVDLA_CSC_wl.scala 807:97:@18372.4]
  wire  _T_4521; // @[NV_NVDLA_CSC_wl.scala 807:91:@18373.4]
  wire  _T_4522; // @[NV_NVDLA_CSC_wl.scala 807:97:@18374.4]
  wire  _T_4523; // @[NV_NVDLA_CSC_wl.scala 807:91:@18375.4]
  wire  _T_4524; // @[NV_NVDLA_CSC_wl.scala 807:97:@18376.4]
  wire  _T_4525; // @[NV_NVDLA_CSC_wl.scala 807:91:@18377.4]
  wire  _T_4526; // @[NV_NVDLA_CSC_wl.scala 807:97:@18378.4]
  wire  _T_4527; // @[NV_NVDLA_CSC_wl.scala 807:91:@18379.4]
  wire  _T_4528; // @[NV_NVDLA_CSC_wl.scala 807:97:@18380.4]
  wire  _T_4529; // @[NV_NVDLA_CSC_wl.scala 807:91:@18381.4]
  wire  _T_4530; // @[NV_NVDLA_CSC_wl.scala 807:97:@18382.4]
  wire  _T_4531; // @[NV_NVDLA_CSC_wl.scala 807:91:@18383.4]
  wire  _T_4532; // @[NV_NVDLA_CSC_wl.scala 807:97:@18384.4]
  wire  _T_4533; // @[NV_NVDLA_CSC_wl.scala 807:91:@18385.4]
  wire  _T_4534; // @[NV_NVDLA_CSC_wl.scala 807:97:@18386.4]
  wire  _T_4535; // @[NV_NVDLA_CSC_wl.scala 807:91:@18387.4]
  wire  _T_4536; // @[NV_NVDLA_CSC_wl.scala 807:97:@18388.4]
  wire  _T_4537; // @[NV_NVDLA_CSC_wl.scala 807:91:@18389.4]
  wire  _T_4538; // @[NV_NVDLA_CSC_wl.scala 807:97:@18390.4]
  wire  _T_4539; // @[NV_NVDLA_CSC_wl.scala 807:91:@18391.4]
  wire  _T_4540; // @[NV_NVDLA_CSC_wl.scala 807:97:@18392.4]
  wire  _T_4541; // @[NV_NVDLA_CSC_wl.scala 807:91:@18393.4]
  wire  _T_4542; // @[NV_NVDLA_CSC_wl.scala 807:97:@18394.4]
  wire  _T_4543; // @[NV_NVDLA_CSC_wl.scala 807:91:@18395.4]
  wire  _T_4544; // @[NV_NVDLA_CSC_wl.scala 807:97:@18396.4]
  wire  _T_4545; // @[NV_NVDLA_CSC_wl.scala 807:91:@18397.4]
  wire  _T_4546; // @[NV_NVDLA_CSC_wl.scala 807:97:@18398.4]
  wire  _T_4547; // @[NV_NVDLA_CSC_wl.scala 807:91:@18399.4]
  wire  _T_4548; // @[NV_NVDLA_CSC_wl.scala 807:97:@18400.4]
  wire  _T_4549; // @[NV_NVDLA_CSC_wl.scala 807:91:@18401.4]
  wire  _T_4550; // @[NV_NVDLA_CSC_wl.scala 807:97:@18402.4]
  wire  _T_4551; // @[NV_NVDLA_CSC_wl.scala 807:91:@18403.4]
  wire  _T_4552; // @[NV_NVDLA_CSC_wl.scala 807:97:@18404.4]
  wire  _T_4553; // @[NV_NVDLA_CSC_wl.scala 807:91:@18405.4]
  wire  _T_4554; // @[NV_NVDLA_CSC_wl.scala 807:97:@18406.4]
  wire  _T_4555; // @[NV_NVDLA_CSC_wl.scala 807:91:@18407.4]
  wire  _T_4556; // @[NV_NVDLA_CSC_wl.scala 807:97:@18408.4]
  wire  _T_4557; // @[NV_NVDLA_CSC_wl.scala 807:91:@18409.4]
  wire  _T_4558; // @[NV_NVDLA_CSC_wl.scala 807:97:@18410.4]
  wire  _T_4559; // @[NV_NVDLA_CSC_wl.scala 807:91:@18411.4]
  wire  _T_4560; // @[NV_NVDLA_CSC_wl.scala 807:97:@18412.4]
  wire  _T_4561; // @[NV_NVDLA_CSC_wl.scala 807:91:@18413.4]
  wire  _T_4562; // @[NV_NVDLA_CSC_wl.scala 807:97:@18414.4]
  wire  _T_4563; // @[NV_NVDLA_CSC_wl.scala 807:91:@18415.4]
  wire  _T_4564; // @[NV_NVDLA_CSC_wl.scala 807:97:@18416.4]
  wire  _T_4565; // @[NV_NVDLA_CSC_wl.scala 807:91:@18417.4]
  wire  _T_4566; // @[NV_NVDLA_CSC_wl.scala 807:97:@18418.4]
  wire  _T_4567; // @[NV_NVDLA_CSC_wl.scala 807:91:@18419.4]
  wire  _T_4568; // @[NV_NVDLA_CSC_wl.scala 807:97:@18420.4]
  wire  _T_4569; // @[NV_NVDLA_CSC_wl.scala 807:91:@18421.4]
  wire  _T_4570; // @[NV_NVDLA_CSC_wl.scala 807:97:@18422.4]
  wire  _T_4571; // @[NV_NVDLA_CSC_wl.scala 807:91:@18423.4]
  wire  _T_4572; // @[NV_NVDLA_CSC_wl.scala 807:97:@18424.4]
  wire  _T_4573; // @[NV_NVDLA_CSC_wl.scala 807:91:@18425.4]
  wire  _T_4574; // @[NV_NVDLA_CSC_wl.scala 807:97:@18426.4]
  wire  _T_4575; // @[NV_NVDLA_CSC_wl.scala 807:91:@18427.4]
  wire  _T_4576; // @[NV_NVDLA_CSC_wl.scala 807:97:@18428.4]
  wire  _T_4577; // @[NV_NVDLA_CSC_wl.scala 807:91:@18429.4]
  wire  _T_4578; // @[NV_NVDLA_CSC_wl.scala 807:97:@18430.4]
  wire  _T_4579; // @[NV_NVDLA_CSC_wl.scala 807:91:@18431.4]
  wire  _T_4580; // @[NV_NVDLA_CSC_wl.scala 807:97:@18432.4]
  wire  _T_4581; // @[NV_NVDLA_CSC_wl.scala 807:91:@18433.4]
  wire  _T_4582; // @[NV_NVDLA_CSC_wl.scala 807:97:@18434.4]
  wire  _T_4583; // @[NV_NVDLA_CSC_wl.scala 807:91:@18435.4]
  wire  _T_4584; // @[NV_NVDLA_CSC_wl.scala 807:97:@18436.4]
  wire  _T_4585; // @[NV_NVDLA_CSC_wl.scala 807:91:@18437.4]
  wire  _T_4586; // @[NV_NVDLA_CSC_wl.scala 807:97:@18438.4]
  wire  _T_4587; // @[NV_NVDLA_CSC_wl.scala 807:91:@18439.4]
  wire  _T_4588; // @[NV_NVDLA_CSC_wl.scala 807:97:@18440.4]
  wire  _T_4589; // @[NV_NVDLA_CSC_wl.scala 807:91:@18441.4]
  wire  _T_4590; // @[NV_NVDLA_CSC_wl.scala 807:97:@18442.4]
  wire  _T_4591; // @[NV_NVDLA_CSC_wl.scala 807:91:@18443.4]
  wire  _T_4592; // @[NV_NVDLA_CSC_wl.scala 807:97:@18444.4]
  wire  _T_4593; // @[NV_NVDLA_CSC_wl.scala 807:91:@18445.4]
  wire  _T_4594; // @[NV_NVDLA_CSC_wl.scala 807:97:@18446.4]
  wire  _T_4595; // @[NV_NVDLA_CSC_wl.scala 807:91:@18447.4]
  wire  _T_4596; // @[NV_NVDLA_CSC_wl.scala 807:97:@18448.4]
  wire  _T_4597; // @[NV_NVDLA_CSC_wl.scala 807:91:@18449.4]
  wire  _T_4598; // @[NV_NVDLA_CSC_wl.scala 807:97:@18450.4]
  wire  _T_4599; // @[NV_NVDLA_CSC_wl.scala 807:91:@18451.4]
  wire  _T_4600; // @[NV_NVDLA_CSC_wl.scala 807:97:@18452.4]
  wire  _T_4601; // @[NV_NVDLA_CSC_wl.scala 807:91:@18453.4]
  wire  _T_4602; // @[NV_NVDLA_CSC_wl.scala 807:97:@18454.4]
  wire  _T_4603; // @[NV_NVDLA_CSC_wl.scala 807:91:@18455.4]
  wire  _T_4604; // @[NV_NVDLA_CSC_wl.scala 807:97:@18456.4]
  wire  _T_4605; // @[NV_NVDLA_CSC_wl.scala 807:91:@18457.4]
  wire  _T_4606; // @[NV_NVDLA_CSC_wl.scala 807:97:@18458.4]
  wire  _T_4607; // @[NV_NVDLA_CSC_wl.scala 807:91:@18459.4]
  wire  _T_4608; // @[NV_NVDLA_CSC_wl.scala 807:97:@18460.4]
  wire  _T_4680; // @[NV_NVDLA_CSC_wl.scala 808:97:@18527.4]
  wire  _T_4682; // @[NV_NVDLA_CSC_wl.scala 808:97:@18529.4]
  wire  _T_4684; // @[NV_NVDLA_CSC_wl.scala 808:97:@18531.4]
  wire  _T_4686; // @[NV_NVDLA_CSC_wl.scala 808:97:@18533.4]
  wire  _T_4688; // @[NV_NVDLA_CSC_wl.scala 808:97:@18535.4]
  wire  _T_4690; // @[NV_NVDLA_CSC_wl.scala 808:97:@18537.4]
  wire  _T_4692; // @[NV_NVDLA_CSC_wl.scala 808:97:@18539.4]
  wire  _T_4694; // @[NV_NVDLA_CSC_wl.scala 808:97:@18541.4]
  wire  _T_4696; // @[NV_NVDLA_CSC_wl.scala 808:97:@18543.4]
  wire  _T_4698; // @[NV_NVDLA_CSC_wl.scala 808:97:@18545.4]
  wire  _T_4700; // @[NV_NVDLA_CSC_wl.scala 808:97:@18547.4]
  wire  _T_4702; // @[NV_NVDLA_CSC_wl.scala 808:97:@18549.4]
  wire  _T_4704; // @[NV_NVDLA_CSC_wl.scala 808:97:@18551.4]
  wire  _T_4706; // @[NV_NVDLA_CSC_wl.scala 808:97:@18553.4]
  wire  _T_4708; // @[NV_NVDLA_CSC_wl.scala 808:97:@18555.4]
  wire  _T_4710; // @[NV_NVDLA_CSC_wl.scala 808:97:@18557.4]
  wire  _T_4712; // @[NV_NVDLA_CSC_wl.scala 808:97:@18559.4]
  wire  _T_4714; // @[NV_NVDLA_CSC_wl.scala 808:97:@18561.4]
  wire  _T_4716; // @[NV_NVDLA_CSC_wl.scala 808:97:@18563.4]
  wire  _T_4718; // @[NV_NVDLA_CSC_wl.scala 808:97:@18565.4]
  wire  _T_4720; // @[NV_NVDLA_CSC_wl.scala 808:97:@18567.4]
  wire  _T_4722; // @[NV_NVDLA_CSC_wl.scala 808:97:@18569.4]
  wire  _T_4724; // @[NV_NVDLA_CSC_wl.scala 808:97:@18571.4]
  wire  _T_4726; // @[NV_NVDLA_CSC_wl.scala 808:97:@18573.4]
  wire  _T_4728; // @[NV_NVDLA_CSC_wl.scala 808:97:@18575.4]
  wire  _T_4730; // @[NV_NVDLA_CSC_wl.scala 808:97:@18577.4]
  wire  _T_4732; // @[NV_NVDLA_CSC_wl.scala 808:97:@18579.4]
  wire  _T_4734; // @[NV_NVDLA_CSC_wl.scala 808:97:@18581.4]
  wire  _T_4736; // @[NV_NVDLA_CSC_wl.scala 808:97:@18583.4]
  wire  _T_4738; // @[NV_NVDLA_CSC_wl.scala 808:97:@18585.4]
  wire  _T_4740; // @[NV_NVDLA_CSC_wl.scala 808:97:@18587.4]
  wire  _T_4742; // @[NV_NVDLA_CSC_wl.scala 808:97:@18589.4]
  wire  _T_4744; // @[NV_NVDLA_CSC_wl.scala 808:97:@18591.4]
  wire  _T_4746; // @[NV_NVDLA_CSC_wl.scala 808:97:@18593.4]
  wire  _T_4748; // @[NV_NVDLA_CSC_wl.scala 808:97:@18595.4]
  wire  _T_4750; // @[NV_NVDLA_CSC_wl.scala 808:97:@18597.4]
  wire  _T_4752; // @[NV_NVDLA_CSC_wl.scala 808:97:@18599.4]
  wire  _T_4754; // @[NV_NVDLA_CSC_wl.scala 808:97:@18601.4]
  wire  _T_4756; // @[NV_NVDLA_CSC_wl.scala 808:97:@18603.4]
  wire  _T_4758; // @[NV_NVDLA_CSC_wl.scala 808:97:@18605.4]
  wire  _T_4760; // @[NV_NVDLA_CSC_wl.scala 808:97:@18607.4]
  wire  _T_4762; // @[NV_NVDLA_CSC_wl.scala 808:97:@18609.4]
  wire  _T_4764; // @[NV_NVDLA_CSC_wl.scala 808:97:@18611.4]
  wire  _T_4766; // @[NV_NVDLA_CSC_wl.scala 808:97:@18613.4]
  wire  _T_4768; // @[NV_NVDLA_CSC_wl.scala 808:97:@18615.4]
  wire  _T_4770; // @[NV_NVDLA_CSC_wl.scala 808:97:@18617.4]
  wire  _T_4772; // @[NV_NVDLA_CSC_wl.scala 808:97:@18619.4]
  wire  _T_4774; // @[NV_NVDLA_CSC_wl.scala 808:97:@18621.4]
  wire  _T_4776; // @[NV_NVDLA_CSC_wl.scala 808:97:@18623.4]
  wire  _T_4778; // @[NV_NVDLA_CSC_wl.scala 808:97:@18625.4]
  wire  _T_4780; // @[NV_NVDLA_CSC_wl.scala 808:97:@18627.4]
  wire  _T_4782; // @[NV_NVDLA_CSC_wl.scala 808:97:@18629.4]
  wire  _T_4784; // @[NV_NVDLA_CSC_wl.scala 808:97:@18631.4]
  wire  _T_4786; // @[NV_NVDLA_CSC_wl.scala 808:97:@18633.4]
  wire  _T_4788; // @[NV_NVDLA_CSC_wl.scala 808:97:@18635.4]
  wire  _T_4790; // @[NV_NVDLA_CSC_wl.scala 808:97:@18637.4]
  wire  _T_4792; // @[NV_NVDLA_CSC_wl.scala 808:97:@18639.4]
  wire  _T_4794; // @[NV_NVDLA_CSC_wl.scala 808:97:@18641.4]
  wire  _T_4796; // @[NV_NVDLA_CSC_wl.scala 808:97:@18643.4]
  wire  _T_4798; // @[NV_NVDLA_CSC_wl.scala 808:97:@18645.4]
  wire  _T_4800; // @[NV_NVDLA_CSC_wl.scala 808:97:@18647.4]
  wire  _T_4802; // @[NV_NVDLA_CSC_wl.scala 808:97:@18649.4]
  wire  _T_4804; // @[NV_NVDLA_CSC_wl.scala 808:97:@18651.4]
  wire  _T_4806; // @[NV_NVDLA_CSC_wl.scala 808:97:@18653.4]
  wire  _T_4877; // @[NV_NVDLA_CSC_wl.scala 812:29:@18721.4]
  wire  _T_4878; // @[NV_NVDLA_CSC_wl.scala 814:96:@18787.6]
  wire  _T_4879; // @[NV_NVDLA_CSC_wl.scala 814:96:@18788.6]
  wire  _T_4880; // @[NV_NVDLA_CSC_wl.scala 814:96:@18789.6]
  wire  _T_4881; // @[NV_NVDLA_CSC_wl.scala 814:96:@18790.6]
  wire  _T_4882; // @[NV_NVDLA_CSC_wl.scala 814:96:@18791.6]
  wire  _T_4883; // @[NV_NVDLA_CSC_wl.scala 814:96:@18792.6]
  wire  _T_4884; // @[NV_NVDLA_CSC_wl.scala 814:96:@18793.6]
  wire  _T_4885; // @[NV_NVDLA_CSC_wl.scala 814:96:@18794.6]
  wire  _T_4886; // @[NV_NVDLA_CSC_wl.scala 814:96:@18795.6]
  wire  _T_4887; // @[NV_NVDLA_CSC_wl.scala 814:96:@18796.6]
  wire  _T_4888; // @[NV_NVDLA_CSC_wl.scala 814:96:@18797.6]
  wire  _T_4889; // @[NV_NVDLA_CSC_wl.scala 814:96:@18798.6]
  wire  _T_4890; // @[NV_NVDLA_CSC_wl.scala 814:96:@18799.6]
  wire  _T_4891; // @[NV_NVDLA_CSC_wl.scala 814:96:@18800.6]
  wire  _T_4892; // @[NV_NVDLA_CSC_wl.scala 814:96:@18801.6]
  wire  _T_4893; // @[NV_NVDLA_CSC_wl.scala 814:96:@18802.6]
  wire  _GEN_209; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_210; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_211; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_212; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_213; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_214; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_215; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_216; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_217; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_218; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_219; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_220; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_221; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_222; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_223; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_224; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_225; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_226; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_227; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_228; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_229; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_230; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_231; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_232; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_233; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_234; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_235; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_236; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_237; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_238; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_239; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_240; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_241; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_242; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_243; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_244; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_245; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_246; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_247; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_248; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_249; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_250; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_251; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_252; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_253; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_254; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_255; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_256; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_257; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_258; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_259; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_260; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_261; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_262; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_263; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_264; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_265; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_266; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_267; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_268; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_269; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_270; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_271; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_272; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_273; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_274; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_275; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_276; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_277; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_278; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_279; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_280; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_281; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_282; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_283; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_284; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_285; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_286; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_287; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _GEN_288; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  wire  _T_4916; // @[NV_NVDLA_CSC_wl.scala 816:29:@18837.4]
  wire  _T_4917; // @[NV_NVDLA_CSC_wl.scala 818:96:@18903.6]
  wire  _T_4918; // @[NV_NVDLA_CSC_wl.scala 818:96:@18904.6]
  wire  _T_4919; // @[NV_NVDLA_CSC_wl.scala 818:96:@18905.6]
  wire  _T_4920; // @[NV_NVDLA_CSC_wl.scala 818:96:@18906.6]
  wire  _T_4921; // @[NV_NVDLA_CSC_wl.scala 818:96:@18907.6]
  wire  _T_4922; // @[NV_NVDLA_CSC_wl.scala 818:96:@18908.6]
  wire  _T_4923; // @[NV_NVDLA_CSC_wl.scala 818:96:@18909.6]
  wire  _T_4924; // @[NV_NVDLA_CSC_wl.scala 818:96:@18910.6]
  wire  _T_4925; // @[NV_NVDLA_CSC_wl.scala 818:96:@18911.6]
  wire  _T_4926; // @[NV_NVDLA_CSC_wl.scala 818:96:@18912.6]
  wire  _T_4927; // @[NV_NVDLA_CSC_wl.scala 818:96:@18913.6]
  wire  _T_4928; // @[NV_NVDLA_CSC_wl.scala 818:96:@18914.6]
  wire  _T_4929; // @[NV_NVDLA_CSC_wl.scala 818:96:@18915.6]
  wire  _T_4930; // @[NV_NVDLA_CSC_wl.scala 818:96:@18916.6]
  wire  _T_4931; // @[NV_NVDLA_CSC_wl.scala 818:96:@18917.6]
  wire  _T_4932; // @[NV_NVDLA_CSC_wl.scala 818:96:@18918.6]
  wire  _GEN_289; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_290; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_291; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_292; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_293; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_294; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_295; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_296; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_297; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_298; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_299; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_300; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_301; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_302; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_303; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_304; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_305; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_306; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_307; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_308; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_309; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_310; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_311; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_312; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_313; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_314; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_315; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_316; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_317; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_318; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_319; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_320; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_321; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_322; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_323; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_324; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_325; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_326; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_327; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_328; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_329; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_330; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_331; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_332; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_333; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_334; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_335; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_336; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_337; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_338; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_339; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_340; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_341; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_342; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_343; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_344; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_345; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_346; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_347; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_348; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_349; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_350; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_351; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_352; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_353; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_354; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_355; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_356; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_357; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_358; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_359; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_360; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_361; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_362; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_363; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_364; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_365; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_366; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_367; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  wire  _GEN_368; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  NV_NVDLA_CSC_WL_dec NV_NVDLA_CSC_WL_dec ( // @[NV_NVDLA_CSC_wl.scala 778:23:@17923.4]
    .reset(NV_NVDLA_CSC_WL_dec_reset),
    .io_nvdla_core_clk(NV_NVDLA_CSC_WL_dec_io_nvdla_core_clk),
    .io_input_valid(NV_NVDLA_CSC_WL_dec_io_input_valid),
    .io_input_bits_mask_0(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_0),
    .io_input_bits_mask_1(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_1),
    .io_input_bits_mask_2(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_2),
    .io_input_bits_mask_3(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_3),
    .io_input_bits_mask_4(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_4),
    .io_input_bits_mask_5(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_5),
    .io_input_bits_mask_6(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_6),
    .io_input_bits_mask_7(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_7),
    .io_input_bits_mask_8(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_8),
    .io_input_bits_mask_9(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_9),
    .io_input_bits_mask_10(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_10),
    .io_input_bits_mask_11(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_11),
    .io_input_bits_mask_12(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_12),
    .io_input_bits_mask_13(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_13),
    .io_input_bits_mask_14(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_14),
    .io_input_bits_mask_15(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_15),
    .io_input_bits_mask_16(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_16),
    .io_input_bits_mask_17(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_17),
    .io_input_bits_mask_18(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_18),
    .io_input_bits_mask_19(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_19),
    .io_input_bits_mask_20(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_20),
    .io_input_bits_mask_21(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_21),
    .io_input_bits_mask_22(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_22),
    .io_input_bits_mask_23(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_23),
    .io_input_bits_mask_24(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_24),
    .io_input_bits_mask_25(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_25),
    .io_input_bits_mask_26(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_26),
    .io_input_bits_mask_27(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_27),
    .io_input_bits_mask_28(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_28),
    .io_input_bits_mask_29(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_29),
    .io_input_bits_mask_30(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_30),
    .io_input_bits_mask_31(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_31),
    .io_input_bits_mask_32(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_32),
    .io_input_bits_mask_33(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_33),
    .io_input_bits_mask_34(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_34),
    .io_input_bits_mask_35(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_35),
    .io_input_bits_mask_36(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_36),
    .io_input_bits_mask_37(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_37),
    .io_input_bits_mask_38(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_38),
    .io_input_bits_mask_39(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_39),
    .io_input_bits_mask_40(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_40),
    .io_input_bits_mask_41(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_41),
    .io_input_bits_mask_42(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_42),
    .io_input_bits_mask_43(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_43),
    .io_input_bits_mask_44(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_44),
    .io_input_bits_mask_45(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_45),
    .io_input_bits_mask_46(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_46),
    .io_input_bits_mask_47(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_47),
    .io_input_bits_mask_48(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_48),
    .io_input_bits_mask_49(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_49),
    .io_input_bits_mask_50(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_50),
    .io_input_bits_mask_51(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_51),
    .io_input_bits_mask_52(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_52),
    .io_input_bits_mask_53(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_53),
    .io_input_bits_mask_54(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_54),
    .io_input_bits_mask_55(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_55),
    .io_input_bits_mask_56(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_56),
    .io_input_bits_mask_57(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_57),
    .io_input_bits_mask_58(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_58),
    .io_input_bits_mask_59(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_59),
    .io_input_bits_mask_60(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_60),
    .io_input_bits_mask_61(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_61),
    .io_input_bits_mask_62(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_62),
    .io_input_bits_mask_63(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_63),
    .io_input_bits_data_0(NV_NVDLA_CSC_WL_dec_io_input_bits_data_0),
    .io_input_bits_data_1(NV_NVDLA_CSC_WL_dec_io_input_bits_data_1),
    .io_input_bits_data_2(NV_NVDLA_CSC_WL_dec_io_input_bits_data_2),
    .io_input_bits_data_3(NV_NVDLA_CSC_WL_dec_io_input_bits_data_3),
    .io_input_bits_data_4(NV_NVDLA_CSC_WL_dec_io_input_bits_data_4),
    .io_input_bits_data_5(NV_NVDLA_CSC_WL_dec_io_input_bits_data_5),
    .io_input_bits_data_6(NV_NVDLA_CSC_WL_dec_io_input_bits_data_6),
    .io_input_bits_data_7(NV_NVDLA_CSC_WL_dec_io_input_bits_data_7),
    .io_input_bits_data_8(NV_NVDLA_CSC_WL_dec_io_input_bits_data_8),
    .io_input_bits_data_9(NV_NVDLA_CSC_WL_dec_io_input_bits_data_9),
    .io_input_bits_data_10(NV_NVDLA_CSC_WL_dec_io_input_bits_data_10),
    .io_input_bits_data_11(NV_NVDLA_CSC_WL_dec_io_input_bits_data_11),
    .io_input_bits_data_12(NV_NVDLA_CSC_WL_dec_io_input_bits_data_12),
    .io_input_bits_data_13(NV_NVDLA_CSC_WL_dec_io_input_bits_data_13),
    .io_input_bits_data_14(NV_NVDLA_CSC_WL_dec_io_input_bits_data_14),
    .io_input_bits_data_15(NV_NVDLA_CSC_WL_dec_io_input_bits_data_15),
    .io_input_bits_data_16(NV_NVDLA_CSC_WL_dec_io_input_bits_data_16),
    .io_input_bits_data_17(NV_NVDLA_CSC_WL_dec_io_input_bits_data_17),
    .io_input_bits_data_18(NV_NVDLA_CSC_WL_dec_io_input_bits_data_18),
    .io_input_bits_data_19(NV_NVDLA_CSC_WL_dec_io_input_bits_data_19),
    .io_input_bits_data_20(NV_NVDLA_CSC_WL_dec_io_input_bits_data_20),
    .io_input_bits_data_21(NV_NVDLA_CSC_WL_dec_io_input_bits_data_21),
    .io_input_bits_data_22(NV_NVDLA_CSC_WL_dec_io_input_bits_data_22),
    .io_input_bits_data_23(NV_NVDLA_CSC_WL_dec_io_input_bits_data_23),
    .io_input_bits_data_24(NV_NVDLA_CSC_WL_dec_io_input_bits_data_24),
    .io_input_bits_data_25(NV_NVDLA_CSC_WL_dec_io_input_bits_data_25),
    .io_input_bits_data_26(NV_NVDLA_CSC_WL_dec_io_input_bits_data_26),
    .io_input_bits_data_27(NV_NVDLA_CSC_WL_dec_io_input_bits_data_27),
    .io_input_bits_data_28(NV_NVDLA_CSC_WL_dec_io_input_bits_data_28),
    .io_input_bits_data_29(NV_NVDLA_CSC_WL_dec_io_input_bits_data_29),
    .io_input_bits_data_30(NV_NVDLA_CSC_WL_dec_io_input_bits_data_30),
    .io_input_bits_data_31(NV_NVDLA_CSC_WL_dec_io_input_bits_data_31),
    .io_input_bits_data_32(NV_NVDLA_CSC_WL_dec_io_input_bits_data_32),
    .io_input_bits_data_33(NV_NVDLA_CSC_WL_dec_io_input_bits_data_33),
    .io_input_bits_data_34(NV_NVDLA_CSC_WL_dec_io_input_bits_data_34),
    .io_input_bits_data_35(NV_NVDLA_CSC_WL_dec_io_input_bits_data_35),
    .io_input_bits_data_36(NV_NVDLA_CSC_WL_dec_io_input_bits_data_36),
    .io_input_bits_data_37(NV_NVDLA_CSC_WL_dec_io_input_bits_data_37),
    .io_input_bits_data_38(NV_NVDLA_CSC_WL_dec_io_input_bits_data_38),
    .io_input_bits_data_39(NV_NVDLA_CSC_WL_dec_io_input_bits_data_39),
    .io_input_bits_data_40(NV_NVDLA_CSC_WL_dec_io_input_bits_data_40),
    .io_input_bits_data_41(NV_NVDLA_CSC_WL_dec_io_input_bits_data_41),
    .io_input_bits_data_42(NV_NVDLA_CSC_WL_dec_io_input_bits_data_42),
    .io_input_bits_data_43(NV_NVDLA_CSC_WL_dec_io_input_bits_data_43),
    .io_input_bits_data_44(NV_NVDLA_CSC_WL_dec_io_input_bits_data_44),
    .io_input_bits_data_45(NV_NVDLA_CSC_WL_dec_io_input_bits_data_45),
    .io_input_bits_data_46(NV_NVDLA_CSC_WL_dec_io_input_bits_data_46),
    .io_input_bits_data_47(NV_NVDLA_CSC_WL_dec_io_input_bits_data_47),
    .io_input_bits_data_48(NV_NVDLA_CSC_WL_dec_io_input_bits_data_48),
    .io_input_bits_data_49(NV_NVDLA_CSC_WL_dec_io_input_bits_data_49),
    .io_input_bits_data_50(NV_NVDLA_CSC_WL_dec_io_input_bits_data_50),
    .io_input_bits_data_51(NV_NVDLA_CSC_WL_dec_io_input_bits_data_51),
    .io_input_bits_data_52(NV_NVDLA_CSC_WL_dec_io_input_bits_data_52),
    .io_input_bits_data_53(NV_NVDLA_CSC_WL_dec_io_input_bits_data_53),
    .io_input_bits_data_54(NV_NVDLA_CSC_WL_dec_io_input_bits_data_54),
    .io_input_bits_data_55(NV_NVDLA_CSC_WL_dec_io_input_bits_data_55),
    .io_input_bits_data_56(NV_NVDLA_CSC_WL_dec_io_input_bits_data_56),
    .io_input_bits_data_57(NV_NVDLA_CSC_WL_dec_io_input_bits_data_57),
    .io_input_bits_data_58(NV_NVDLA_CSC_WL_dec_io_input_bits_data_58),
    .io_input_bits_data_59(NV_NVDLA_CSC_WL_dec_io_input_bits_data_59),
    .io_input_bits_data_60(NV_NVDLA_CSC_WL_dec_io_input_bits_data_60),
    .io_input_bits_data_61(NV_NVDLA_CSC_WL_dec_io_input_bits_data_61),
    .io_input_bits_data_62(NV_NVDLA_CSC_WL_dec_io_input_bits_data_62),
    .io_input_bits_data_63(NV_NVDLA_CSC_WL_dec_io_input_bits_data_63),
    .io_input_bits_sel_0(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_0),
    .io_input_bits_sel_1(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_1),
    .io_input_bits_sel_2(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_2),
    .io_input_bits_sel_3(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_3),
    .io_input_bits_sel_4(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_4),
    .io_input_bits_sel_5(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_5),
    .io_input_bits_sel_6(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_6),
    .io_input_bits_sel_7(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_7),
    .io_input_bits_sel_8(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_8),
    .io_input_bits_sel_9(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_9),
    .io_input_bits_sel_10(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_10),
    .io_input_bits_sel_11(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_11),
    .io_input_bits_sel_12(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_12),
    .io_input_bits_sel_13(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_13),
    .io_input_bits_sel_14(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_14),
    .io_input_bits_sel_15(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_15),
    .io_input_bits_sel_16(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_16),
    .io_input_bits_sel_17(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_17),
    .io_input_bits_sel_18(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_18),
    .io_input_bits_sel_19(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_19),
    .io_input_bits_sel_20(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_20),
    .io_input_bits_sel_21(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_21),
    .io_input_bits_sel_22(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_22),
    .io_input_bits_sel_23(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_23),
    .io_input_bits_sel_24(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_24),
    .io_input_bits_sel_25(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_25),
    .io_input_bits_sel_26(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_26),
    .io_input_bits_sel_27(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_27),
    .io_input_bits_sel_28(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_28),
    .io_input_bits_sel_29(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_29),
    .io_input_bits_sel_30(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_30),
    .io_input_bits_sel_31(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_31),
    .io_input_mask_en(NV_NVDLA_CSC_WL_dec_io_input_mask_en),
    .io_output_valid(NV_NVDLA_CSC_WL_dec_io_output_valid),
    .io_output_bits_mask_0(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_0),
    .io_output_bits_mask_1(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_1),
    .io_output_bits_mask_2(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_2),
    .io_output_bits_mask_3(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_3),
    .io_output_bits_mask_4(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_4),
    .io_output_bits_mask_5(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_5),
    .io_output_bits_mask_6(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_6),
    .io_output_bits_mask_7(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_7),
    .io_output_bits_mask_8(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_8),
    .io_output_bits_mask_9(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_9),
    .io_output_bits_mask_10(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_10),
    .io_output_bits_mask_11(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_11),
    .io_output_bits_mask_12(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_12),
    .io_output_bits_mask_13(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_13),
    .io_output_bits_mask_14(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_14),
    .io_output_bits_mask_15(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_15),
    .io_output_bits_mask_16(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_16),
    .io_output_bits_mask_17(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_17),
    .io_output_bits_mask_18(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_18),
    .io_output_bits_mask_19(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_19),
    .io_output_bits_mask_20(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_20),
    .io_output_bits_mask_21(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_21),
    .io_output_bits_mask_22(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_22),
    .io_output_bits_mask_23(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_23),
    .io_output_bits_mask_24(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_24),
    .io_output_bits_mask_25(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_25),
    .io_output_bits_mask_26(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_26),
    .io_output_bits_mask_27(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_27),
    .io_output_bits_mask_28(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_28),
    .io_output_bits_mask_29(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_29),
    .io_output_bits_mask_30(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_30),
    .io_output_bits_mask_31(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_31),
    .io_output_bits_mask_32(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_32),
    .io_output_bits_mask_33(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_33),
    .io_output_bits_mask_34(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_34),
    .io_output_bits_mask_35(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_35),
    .io_output_bits_mask_36(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_36),
    .io_output_bits_mask_37(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_37),
    .io_output_bits_mask_38(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_38),
    .io_output_bits_mask_39(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_39),
    .io_output_bits_mask_40(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_40),
    .io_output_bits_mask_41(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_41),
    .io_output_bits_mask_42(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_42),
    .io_output_bits_mask_43(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_43),
    .io_output_bits_mask_44(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_44),
    .io_output_bits_mask_45(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_45),
    .io_output_bits_mask_46(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_46),
    .io_output_bits_mask_47(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_47),
    .io_output_bits_mask_48(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_48),
    .io_output_bits_mask_49(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_49),
    .io_output_bits_mask_50(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_50),
    .io_output_bits_mask_51(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_51),
    .io_output_bits_mask_52(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_52),
    .io_output_bits_mask_53(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_53),
    .io_output_bits_mask_54(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_54),
    .io_output_bits_mask_55(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_55),
    .io_output_bits_mask_56(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_56),
    .io_output_bits_mask_57(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_57),
    .io_output_bits_mask_58(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_58),
    .io_output_bits_mask_59(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_59),
    .io_output_bits_mask_60(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_60),
    .io_output_bits_mask_61(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_61),
    .io_output_bits_mask_62(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_62),
    .io_output_bits_mask_63(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_63),
    .io_output_bits_data_0(NV_NVDLA_CSC_WL_dec_io_output_bits_data_0),
    .io_output_bits_data_1(NV_NVDLA_CSC_WL_dec_io_output_bits_data_1),
    .io_output_bits_data_2(NV_NVDLA_CSC_WL_dec_io_output_bits_data_2),
    .io_output_bits_data_3(NV_NVDLA_CSC_WL_dec_io_output_bits_data_3),
    .io_output_bits_data_4(NV_NVDLA_CSC_WL_dec_io_output_bits_data_4),
    .io_output_bits_data_5(NV_NVDLA_CSC_WL_dec_io_output_bits_data_5),
    .io_output_bits_data_6(NV_NVDLA_CSC_WL_dec_io_output_bits_data_6),
    .io_output_bits_data_7(NV_NVDLA_CSC_WL_dec_io_output_bits_data_7),
    .io_output_bits_data_8(NV_NVDLA_CSC_WL_dec_io_output_bits_data_8),
    .io_output_bits_data_9(NV_NVDLA_CSC_WL_dec_io_output_bits_data_9),
    .io_output_bits_data_10(NV_NVDLA_CSC_WL_dec_io_output_bits_data_10),
    .io_output_bits_data_11(NV_NVDLA_CSC_WL_dec_io_output_bits_data_11),
    .io_output_bits_data_12(NV_NVDLA_CSC_WL_dec_io_output_bits_data_12),
    .io_output_bits_data_13(NV_NVDLA_CSC_WL_dec_io_output_bits_data_13),
    .io_output_bits_data_14(NV_NVDLA_CSC_WL_dec_io_output_bits_data_14),
    .io_output_bits_data_15(NV_NVDLA_CSC_WL_dec_io_output_bits_data_15),
    .io_output_bits_data_16(NV_NVDLA_CSC_WL_dec_io_output_bits_data_16),
    .io_output_bits_data_17(NV_NVDLA_CSC_WL_dec_io_output_bits_data_17),
    .io_output_bits_data_18(NV_NVDLA_CSC_WL_dec_io_output_bits_data_18),
    .io_output_bits_data_19(NV_NVDLA_CSC_WL_dec_io_output_bits_data_19),
    .io_output_bits_data_20(NV_NVDLA_CSC_WL_dec_io_output_bits_data_20),
    .io_output_bits_data_21(NV_NVDLA_CSC_WL_dec_io_output_bits_data_21),
    .io_output_bits_data_22(NV_NVDLA_CSC_WL_dec_io_output_bits_data_22),
    .io_output_bits_data_23(NV_NVDLA_CSC_WL_dec_io_output_bits_data_23),
    .io_output_bits_data_24(NV_NVDLA_CSC_WL_dec_io_output_bits_data_24),
    .io_output_bits_data_25(NV_NVDLA_CSC_WL_dec_io_output_bits_data_25),
    .io_output_bits_data_26(NV_NVDLA_CSC_WL_dec_io_output_bits_data_26),
    .io_output_bits_data_27(NV_NVDLA_CSC_WL_dec_io_output_bits_data_27),
    .io_output_bits_data_28(NV_NVDLA_CSC_WL_dec_io_output_bits_data_28),
    .io_output_bits_data_29(NV_NVDLA_CSC_WL_dec_io_output_bits_data_29),
    .io_output_bits_data_30(NV_NVDLA_CSC_WL_dec_io_output_bits_data_30),
    .io_output_bits_data_31(NV_NVDLA_CSC_WL_dec_io_output_bits_data_31),
    .io_output_bits_data_32(NV_NVDLA_CSC_WL_dec_io_output_bits_data_32),
    .io_output_bits_data_33(NV_NVDLA_CSC_WL_dec_io_output_bits_data_33),
    .io_output_bits_data_34(NV_NVDLA_CSC_WL_dec_io_output_bits_data_34),
    .io_output_bits_data_35(NV_NVDLA_CSC_WL_dec_io_output_bits_data_35),
    .io_output_bits_data_36(NV_NVDLA_CSC_WL_dec_io_output_bits_data_36),
    .io_output_bits_data_37(NV_NVDLA_CSC_WL_dec_io_output_bits_data_37),
    .io_output_bits_data_38(NV_NVDLA_CSC_WL_dec_io_output_bits_data_38),
    .io_output_bits_data_39(NV_NVDLA_CSC_WL_dec_io_output_bits_data_39),
    .io_output_bits_data_40(NV_NVDLA_CSC_WL_dec_io_output_bits_data_40),
    .io_output_bits_data_41(NV_NVDLA_CSC_WL_dec_io_output_bits_data_41),
    .io_output_bits_data_42(NV_NVDLA_CSC_WL_dec_io_output_bits_data_42),
    .io_output_bits_data_43(NV_NVDLA_CSC_WL_dec_io_output_bits_data_43),
    .io_output_bits_data_44(NV_NVDLA_CSC_WL_dec_io_output_bits_data_44),
    .io_output_bits_data_45(NV_NVDLA_CSC_WL_dec_io_output_bits_data_45),
    .io_output_bits_data_46(NV_NVDLA_CSC_WL_dec_io_output_bits_data_46),
    .io_output_bits_data_47(NV_NVDLA_CSC_WL_dec_io_output_bits_data_47),
    .io_output_bits_data_48(NV_NVDLA_CSC_WL_dec_io_output_bits_data_48),
    .io_output_bits_data_49(NV_NVDLA_CSC_WL_dec_io_output_bits_data_49),
    .io_output_bits_data_50(NV_NVDLA_CSC_WL_dec_io_output_bits_data_50),
    .io_output_bits_data_51(NV_NVDLA_CSC_WL_dec_io_output_bits_data_51),
    .io_output_bits_data_52(NV_NVDLA_CSC_WL_dec_io_output_bits_data_52),
    .io_output_bits_data_53(NV_NVDLA_CSC_WL_dec_io_output_bits_data_53),
    .io_output_bits_data_54(NV_NVDLA_CSC_WL_dec_io_output_bits_data_54),
    .io_output_bits_data_55(NV_NVDLA_CSC_WL_dec_io_output_bits_data_55),
    .io_output_bits_data_56(NV_NVDLA_CSC_WL_dec_io_output_bits_data_56),
    .io_output_bits_data_57(NV_NVDLA_CSC_WL_dec_io_output_bits_data_57),
    .io_output_bits_data_58(NV_NVDLA_CSC_WL_dec_io_output_bits_data_58),
    .io_output_bits_data_59(NV_NVDLA_CSC_WL_dec_io_output_bits_data_59),
    .io_output_bits_data_60(NV_NVDLA_CSC_WL_dec_io_output_bits_data_60),
    .io_output_bits_data_61(NV_NVDLA_CSC_WL_dec_io_output_bits_data_61),
    .io_output_bits_data_62(NV_NVDLA_CSC_WL_dec_io_output_bits_data_62),
    .io_output_bits_data_63(NV_NVDLA_CSC_WL_dec_io_output_bits_data_63),
    .io_output_bits_sel_0(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_0),
    .io_output_bits_sel_1(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_1),
    .io_output_bits_sel_2(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_2),
    .io_output_bits_sel_3(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_3),
    .io_output_bits_sel_4(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_4),
    .io_output_bits_sel_5(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_5),
    .io_output_bits_sel_6(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_6),
    .io_output_bits_sel_7(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_7),
    .io_output_bits_sel_8(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_8),
    .io_output_bits_sel_9(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_9),
    .io_output_bits_sel_10(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_10),
    .io_output_bits_sel_11(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_11),
    .io_output_bits_sel_12(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_12),
    .io_output_bits_sel_13(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_13),
    .io_output_bits_sel_14(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_14),
    .io_output_bits_sel_15(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_15),
    .io_output_bits_sel_16(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_16),
    .io_output_bits_sel_17(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_17),
    .io_output_bits_sel_18(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_18),
    .io_output_bits_sel_19(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_19),
    .io_output_bits_sel_20(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_20),
    .io_output_bits_sel_21(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_21),
    .io_output_bits_sel_22(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_22),
    .io_output_bits_sel_23(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_23),
    .io_output_bits_sel_24(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_24),
    .io_output_bits_sel_25(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_25),
    .io_output_bits_sel_26(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_26),
    .io_output_bits_sel_27(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_27),
    .io_output_bits_sel_28(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_28),
    .io_output_bits_sel_29(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_29),
    .io_output_bits_sel_30(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_30),
    .io_output_bits_sel_31(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_31)
  );
  assign _T_700 = io_sc_state == 2'h0; // @[NV_NVDLA_CSC_wl.scala 97:35:@16374.4]
  assign _T_704 = io_sc_state == 2'h2; // @[NV_NVDLA_CSC_wl.scala 99:38:@16376.4]
  assign _T_706 = io_sc_state == 2'h3; // @[NV_NVDLA_CSC_wl.scala 100:35:@16377.4]
  assign _T_707 = ~ _T_698; // @[NV_NVDLA_CSC_wl.scala 101:37:@16378.4]
  assign _T_708 = _T_704 & _T_707; // @[NV_NVDLA_CSC_wl.scala 101:35:@16379.4]
  assign _T_743 = io_reg2dp_op_en & _T_700; // @[NV_NVDLA_CSC_wl.scala 115:36:@16391.4]
  assign _T_749 = io_reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CSC_wl.scala 120:42:@16395.6]
  assign _T_750 = io_reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CSC_wl.scala 120:42:@16396.6]
  assign _T_752 = io_reg2dp_weight_bank + 5'h1; // @[NV_NVDLA_CSC_wl.scala 121:46:@16398.6]
  assign _T_753 = io_reg2dp_weight_bank + 5'h1; // @[NV_NVDLA_CSC_wl.scala 121:46:@16399.6]
  assign _T_755 = 9'h9 << io_reg2dp_y_extension; // @[NV_NVDLA_CSC_wl.scala 122:42:@16401.6]
  assign _T_756 = _T_755[5:3]; // @[NV_NVDLA_CSC_wl.scala 122:67:@16402.6]
  assign _GEN_0 = _T_743 ? _T_750 : _T_715; // @[NV_NVDLA_CSC_wl.scala 119:19:@16394.4]
  assign _GEN_1 = _T_743 ? _T_753 : _T_722; // @[NV_NVDLA_CSC_wl.scala 119:19:@16394.4]
  assign _GEN_2 = _T_743 ? _T_756 : _T_739; // @[NV_NVDLA_CSC_wl.scala 119:19:@16394.4]
  assign _GEN_3 = _T_743 ? io_reg2dp_weight_format : _T_742; // @[NV_NVDLA_CSC_wl.scala 119:19:@16394.4]
  assign _T_757 = _T_706 & io_reg2dp_skip_weight_rls; // @[NV_NVDLA_CSC_wl.scala 125:21:@16406.4]
  assign _T_758 = io_reg2dp_weight_bytes[20:6]; // @[NV_NVDLA_CSC_wl.scala 126:54:@16408.6]
  assign _T_759 = io_reg2dp_wmb_bytes[14:6]; // @[NV_NVDLA_CSC_wl.scala 127:70:@16410.6]
  assign _T_761 = _T_742 ? _T_759 : 9'h0; // @[NV_NVDLA_CSC_wl.scala 127:32:@16411.6]
  assign _GEN_4 = _T_757 ? _T_758 : _T_729; // @[NV_NVDLA_CSC_wl.scala 125:49:@16407.4]
  assign _GEN_5 = _T_757 ? _T_761 : _T_736; // @[NV_NVDLA_CSC_wl.scala 125:49:@16407.4]
  assign _T_1759 = _T_1712[35]; // @[NV_NVDLA_CSC_wl.scala 693:34:@17289.4]
  assign _T_857 = _T_1692 & _T_1759; // @[NV_NVDLA_CSC_wl.scala 203:36:@16489.4]
  assign _T_858 = io_sg2wl_reuse_rls | _T_857; // @[NV_NVDLA_CSC_wl.scala 207:25:@16490.4]
  assign _T_1755 = _T_1712[31:17]; // @[NV_NVDLA_CSC_wl.scala 689:44:@17284.4]
  assign _T_859 = io_sg2wl_reuse_rls ? _T_729 : _T_1755; // @[NV_NVDLA_CSC_wl.scala 208:29:@16492.4]
  assign _T_1754 = _T_1712[16:8]; // @[NV_NVDLA_CSC_wl.scala 688:45:@17282.4]
  assign _T_860 = io_sg2wl_reuse_rls ? _T_736 : _T_1754; // @[NV_NVDLA_CSC_wl.scala 209:30:@16494.4]
  assign _T_799 = _T_798 + _T_859; // @[NV_NVDLA_CSC_wl.scala 155:39:@16436.4]
  assign _T_800 = _T_798 + _T_859; // @[NV_NVDLA_CSC_wl.scala 155:39:@16437.4]
  assign _T_802 = {_T_722,9'h0}; // @[Cat.scala 30:58:@16438.4]
  assign _GEN_497 = {{1'd0}, _T_802}; // @[NV_NVDLA_CSC_wl.scala 156:48:@16439.4]
  assign _T_803 = _T_800 - _GEN_497; // @[NV_NVDLA_CSC_wl.scala 156:48:@16439.4]
  assign _T_804 = $unsigned(_T_803); // @[NV_NVDLA_CSC_wl.scala 156:48:@16440.4]
  assign _T_805 = _T_804[14:0]; // @[NV_NVDLA_CSC_wl.scala 156:48:@16441.4]
  assign _T_808 = _T_800 >= _GEN_497; // @[NV_NVDLA_CSC_wl.scala 157:48:@16443.4]
  assign _T_810 = ~ _T_858; // @[NV_NVDLA_CSC_wl.scala 158:88:@16444.4]
  assign _T_811 = _T_808 ? _T_805 : _T_800; // @[NV_NVDLA_CSC_wl.scala 158:113:@16445.4]
  assign _T_812 = _T_810 ? _T_798 : _T_811; // @[NV_NVDLA_CSC_wl.scala 158:87:@16446.4]
  assign _T_813 = io_sc2cdma_wt_pending_req ? 15'h0 : _T_812; // @[NV_NVDLA_CSC_wl.scala 158:28:@16447.4]
  assign _T_847 = io_sc2cdma_wt_pending_req | _T_858; // @[NV_NVDLA_CSC_wl.scala 184:21:@16475.4]
  assign _GEN_8 = _T_847 ? _T_813 : _T_798; // @[NV_NVDLA_CSC_wl.scala 184:30:@16476.4]
  assign _GEN_12 = _T_858 ? _T_859 : _T_867; // @[Reg.scala 20:19:@16501.4]
  assign _GEN_13 = _T_858 ? _T_860 : _T_871; // @[Reg.scala 20:19:@16507.4]
  assign _T_879 = io_sg2wl_pd_bits[0]; // @[NV_NVDLA_CSC_wl.scala 224:26:@16514.4 NV_NVDLA_CSC_wl.scala 228:19:@16517.4]
  assign _GEN_14 = io_sg2wl_pd_valid ? {{17'd0}, _T_879} : _T_882; // @[NV_NVDLA_CSC_wl.scala 232:30:@16519.4]
  assign _T_883 = _T_882[6:0]; // @[NV_NVDLA_CSC_wl.scala 241:31:@16522.4]
  assign _T_884 = _T_882[12:7]; // @[NV_NVDLA_CSC_wl.scala 242:31:@16523.4]
  assign _T_885 = _T_882[14:13]; // @[NV_NVDLA_CSC_wl.scala 243:29:@16524.4]
  assign _T_886 = _T_882[15]; // @[NV_NVDLA_CSC_wl.scala 244:31:@16525.4]
  assign _T_887 = _T_882[16]; // @[NV_NVDLA_CSC_wl.scala 245:29:@16526.4]
  assign _T_888 = _T_882[17]; // @[NV_NVDLA_CSC_wl.scala 246:30:@16527.4]
  assign _T_898 = _T_893 + 5'h1; // @[NV_NVDLA_CSC_wl.scala 257:37:@16531.4]
  assign _T_899 = _T_893 + 5'h1; // @[NV_NVDLA_CSC_wl.scala 257:37:@16532.4]
  assign _T_904 = _T_884[4:0]; // @[NV_NVDLA_CSC_wl.scala 259:39:@16535.4]
  assign _T_905 = _T_899 == _T_904; // @[NV_NVDLA_CSC_wl.scala 260:38:@16536.4]
  assign _T_902 = _T_905 ? 5'h0 : _T_899; // @[NV_NVDLA_CSC_wl.scala 258:59:@16533.4]
  assign _T_903 = _T_743 ? 5'h0 : _T_902; // @[NV_NVDLA_CSC_wl.scala 258:27:@16534.4]
  assign _T_908 = _T_893 != 5'h0; // @[NV_NVDLA_CSC_wl.scala 262:64:@16538.4]
  assign _T_909 = ~ _T_908; // @[NV_NVDLA_CSC_wl.scala 262:51:@16539.4]
  assign _T_911 = _T_909 ? 1'h0 : _T_896; // @[NV_NVDLA_CSC_wl.scala 262:50:@16540.4]
  assign _T_912 = _T_877 ? 1'h1 : _T_911; // @[NV_NVDLA_CSC_wl.scala 262:29:@16541.4]
  assign _T_913 = _T_743 | _T_912; // @[NV_NVDLA_CSC_wl.scala 263:38:@16542.4]
  assign _GEN_15 = _T_913 ? _T_903 : _T_893; // @[NV_NVDLA_CSC_wl.scala 265:28:@16543.4]
  assign _T_966 = _T_912 & _T_742; // @[NV_NVDLA_CSC_wl.scala 289:37:@16580.4]
  assign _T_964 = 2'h0 == _T_885; // @[Mux.scala 46:19:@16577.4]
  assign _T_942 = {1'h0,_T_883}; // @[Cat.scala 30:58:@16563.4]
  assign _T_962 = 2'h1 == _T_885; // @[Mux.scala 46:19:@16575.4]
  assign _T_951 = _T_942[6:0]; // @[NV_NVDLA_CSC_wl.scala 285:101:@16567.4]
  assign _T_954 = {1'h0,_T_951,1'h0}; // @[Cat.scala 30:58:@16569.4]
  assign _T_960 = 2'h2 == _T_885; // @[Mux.scala 46:19:@16573.4]
  assign _T_958 = {_T_951,1'h0}; // @[Cat.scala 30:58:@16571.4]
  assign _T_959 = _T_958 + _T_942; // @[NV_NVDLA_CSC_wl.scala 286:109:@16572.4]
  assign _T_944 = _T_942[5:0]; // @[NV_NVDLA_CSC_wl.scala 282:92:@16564.4]
  assign _T_947 = {1'h0,_T_944,2'h0}; // @[Cat.scala 30:58:@16566.4]
  assign _T_961 = _T_960 ? _T_959 : _T_947; // @[Mux.scala 46:16:@16574.4]
  assign _T_963 = _T_962 ? _T_954 : _T_961; // @[Mux.scala 46:16:@16576.4]
  assign _T_965 = _T_964 ? {{1'd0}, _T_942} : _T_963; // @[Mux.scala 46:16:@16578.4]
  assign _T_917 = _T_965[7:0]; // @[NV_NVDLA_CSC_wl.scala 271:31:@16547.4 NV_NVDLA_CSC_wl.scala 282:21:@16579.4]
  assign _T_968 = {3'h0,_T_917}; // @[Cat.scala 30:58:@16581.4]
  assign _T_969 = _T_920 < _T_968; // @[NV_NVDLA_CSC_wl.scala 289:75:@16582.4]
  assign _T_970 = _T_966 & _T_969; // @[NV_NVDLA_CSC_wl.scala 289:56:@16583.4]
  assign _T_924 = ~ _T_970; // @[NV_NVDLA_CSC_wl.scala 275:35:@16550.4]
  assign _T_927 = _T_924 ? 11'h0 : 11'h200; // @[NV_NVDLA_CSC_wl.scala 275:34:@16551.4]
  assign _T_929 = _T_912 ? _T_917 : 8'h0; // @[NV_NVDLA_CSC_wl.scala 276:34:@16552.4]
  assign _T_930 = _T_920 + _T_927; // @[NV_NVDLA_CSC_wl.scala 277:47:@16553.4]
  assign _T_931 = _T_920 + _T_927; // @[NV_NVDLA_CSC_wl.scala 277:47:@16554.4]
  assign _GEN_501 = {{3'd0}, _T_929}; // @[NV_NVDLA_CSC_wl.scala 277:69:@16555.4]
  assign _T_932 = _T_931 - _GEN_501; // @[NV_NVDLA_CSC_wl.scala 277:69:@16555.4]
  assign _T_933 = $unsigned(_T_932); // @[NV_NVDLA_CSC_wl.scala 277:69:@16556.4]
  assign _T_934 = _T_933[10:0]; // @[NV_NVDLA_CSC_wl.scala 277:69:@16557.4]
  assign _T_936 = ~ _T_887; // @[NV_NVDLA_CSC_wl.scala 278:82:@16558.4]
  assign _T_937 = _T_905 & _T_936; // @[NV_NVDLA_CSC_wl.scala 278:80:@16559.4]
  assign _T_938 = _T_937 & _T_886; // @[NV_NVDLA_CSC_wl.scala 278:96:@16560.4]
  assign _T_939 = _T_938 ? _T_923 : _T_934; // @[NV_NVDLA_CSC_wl.scala 278:65:@16561.4]
  assign _T_940 = _T_743 ? 11'h0 : _T_939; // @[NV_NVDLA_CSC_wl.scala 278:32:@16562.4]
  assign _T_972 = _T_743 | _T_966; // @[NV_NVDLA_CSC_wl.scala 290:43:@16586.4]
  assign _T_974 = _T_966 & _T_905; // @[NV_NVDLA_CSC_wl.scala 291:85:@16588.4]
  assign _T_975 = _T_974 & _T_887; // @[NV_NVDLA_CSC_wl.scala 291:101:@16589.4]
  assign _T_976 = _T_743 | _T_975; // @[NV_NVDLA_CSC_wl.scala 291:48:@16590.4]
  assign _GEN_16 = _T_972 ? _T_940 : _T_920; // @[NV_NVDLA_CSC_wl.scala 293:33:@16591.4]
  assign _GEN_17 = _T_976 ? _T_940 : _T_923; // @[NV_NVDLA_CSC_wl.scala 296:38:@16594.4]
  assign _T_1007 = _T_887 & _T_905; // @[NV_NVDLA_CSC_wl.scala 321:58:@16624.4]
  assign _T_1008 = _T_743 | _T_1007; // @[NV_NVDLA_CSC_wl.scala 321:42:@16625.4]
  assign _T_1010 = _T_886 & _T_905; // @[NV_NVDLA_CSC_wl.scala 322:48:@16626.4]
  assign _T_1012 = _T_1010 ? 1'h1 : _T_1003; // @[NV_NVDLA_CSC_wl.scala 322:32:@16627.4]
  assign _T_1013 = _T_1008 ? 1'h0 : _T_1012; // @[NV_NVDLA_CSC_wl.scala 321:32:@16628.4]
  assign _T_1015 = _T_1006 + 9'h1; // @[NV_NVDLA_CSC_wl.scala 323:39:@16629.4]
  assign _T_1016 = _T_1006 + 9'h1; // @[NV_NVDLA_CSC_wl.scala 323:39:@16630.4]
  assign _T_1018 = _T_905 & _T_887; // @[NV_NVDLA_CSC_wl.scala 325:43:@16631.4]
  assign _T_1020 = _T_1018 ? 9'h0 : _T_1016; // @[NV_NVDLA_CSC_wl.scala 325:28:@16632.4]
  assign _T_1021 = _T_743 ? 9'h0 : _T_1020; // @[NV_NVDLA_CSC_wl.scala 324:28:@16633.4]
  assign _T_1022 = _T_742 & _T_912; // @[NV_NVDLA_CSC_wl.scala 326:58:@16634.4]
  assign _T_1023 = _T_1022 & _T_905; // @[NV_NVDLA_CSC_wl.scala 326:75:@16635.4]
  assign _T_1024 = _T_1023 & _T_887; // @[NV_NVDLA_CSC_wl.scala 326:91:@16636.4]
  assign _T_1025 = _T_743 | _T_1024; // @[NV_NVDLA_CSC_wl.scala 326:39:@16637.4]
  assign _T_1026 = _T_742 & _T_970; // @[NV_NVDLA_CSC_wl.scala 326:126:@16638.4]
  assign _T_1027 = ~ _T_1003; // @[NV_NVDLA_CSC_wl.scala 326:144:@16639.4]
  assign _T_1028 = _T_1026 & _T_1027; // @[NV_NVDLA_CSC_wl.scala 326:142:@16640.4]
  assign _T_1029 = _T_1025 | _T_1028; // @[NV_NVDLA_CSC_wl.scala 326:107:@16641.4]
  assign _T_1031 = _T_1003 | _T_924; // @[NV_NVDLA_CSC_wl.scala 327:47:@16643.4]
  assign _T_1032 = _T_1031 ? _T_1006 : _T_1016; // @[NV_NVDLA_CSC_wl.scala 327:30:@16644.4]
  assign _GEN_20 = _T_1029 ? _T_1021 : _T_1006; // @[NV_NVDLA_CSC_wl.scala 330:29:@16646.4]
  assign _GEN_22 = _T_912 ? _T_883 : _T_1041; // @[NV_NVDLA_CSC_wl.scala 351:25:@16664.4]
  assign _GEN_23 = _T_912 ? _T_917 : _T_1044; // @[NV_NVDLA_CSC_wl.scala 351:25:@16664.4]
  assign _T_1063 = _T_912 & _T_888; // @[NV_NVDLA_CSC_wl.scala 355:25:@16668.4]
  assign _T_1064 = _T_1063 & _T_905; // @[NV_NVDLA_CSC_wl.scala 355:41:@16669.4]
  assign _GEN_24 = _T_1064 ? _T_1032 : _T_1047; // @[NV_NVDLA_CSC_wl.scala 355:57:@16670.4]
  assign _T_1067 = _T_888 & _T_905; // @[NV_NVDLA_CSC_wl.scala 362:41:@16679.6]
  assign _GEN_25 = _T_912 ? _T_905 : _T_1050; // @[NV_NVDLA_CSC_wl.scala 358:25:@16673.4]
  assign _GEN_26 = _T_912 ? _T_1010 : _T_1053; // @[NV_NVDLA_CSC_wl.scala 358:25:@16673.4]
  assign _GEN_27 = _T_912 ? _T_1007 : _T_1056; // @[NV_NVDLA_CSC_wl.scala 358:25:@16673.4]
  assign _GEN_28 = _T_912 ? _T_1067 : _T_1059; // @[NV_NVDLA_CSC_wl.scala 358:25:@16673.4]
  assign _GEN_29 = _T_912 ? _T_885 : _T_1062; // @[NV_NVDLA_CSC_wl.scala 358:25:@16673.4]
  assign _T_1076 = {_T_1062,1'h0,_T_1059,_T_1056,_T_1053,_T_1050,_T_1047,_T_1044,_T_1041}; // @[Cat.scala 30:58:@16690.4]
  assign _GEN_30 = _T_896 ? _T_1076 : _T_1101; // @[NV_NVDLA_CSC_wl.scala 394:37:@16708.4]
  assign _GEN_31 = _T_1081 ? _T_1101 : _T_1104; // @[NV_NVDLA_CSC_wl.scala 394:37:@16712.4]
  assign _GEN_32 = _T_1084 ? _T_1104 : _T_1107; // @[NV_NVDLA_CSC_wl.scala 394:37:@16716.4]
  assign _GEN_33 = _T_1087 ? _T_1107 : _T_1110; // @[NV_NVDLA_CSC_wl.scala 394:37:@16720.4]
  assign _GEN_34 = _T_1090 ? _T_1110 : _T_1113; // @[NV_NVDLA_CSC_wl.scala 394:37:@16724.4]
  assign _GEN_35 = _T_1093 ? _T_1113 : _T_1116; // @[NV_NVDLA_CSC_wl.scala 394:37:@16728.4]
  assign _T_1117 = _T_1116[6:0]; // @[NV_NVDLA_CSC_wl.scala 404:46:@16731.4]
  assign _T_1118 = _T_1116[14:7]; // @[NV_NVDLA_CSC_wl.scala 405:42:@16732.4]
  assign _T_1119 = _T_1116[23:15]; // @[NV_NVDLA_CSC_wl.scala 406:46:@16733.4]
  assign _T_1120 = _T_1116[24]; // @[NV_NVDLA_CSC_wl.scala 407:45:@16734.4]
  assign _T_1121 = _T_1116[25]; // @[NV_NVDLA_CSC_wl.scala 408:46:@16735.4]
  assign _T_1122 = _T_1116[26]; // @[NV_NVDLA_CSC_wl.scala 409:44:@16736.4]
  assign _T_1123 = _T_1116[27]; // @[NV_NVDLA_CSC_wl.scala 410:38:@16737.4]
  assign _T_1124 = _T_1116[30:29]; // @[NV_NVDLA_CSC_wl.scala 411:44:@16738.4]
  assign _T_1137 = ~ _T_1122; // @[NV_NVDLA_CSC_wl.scala 421:91:@16743.4]
  assign _T_1138 = _T_1121 & _T_1137; // @[NV_NVDLA_CSC_wl.scala 421:89:@16744.4]
  assign _T_1145 = _T_1096 & _T_1122; // @[NV_NVDLA_CSC_wl.scala 422:72:@16751.4]
  assign _T_1146 = _T_1145 & _T_742; // @[NV_NVDLA_CSC_wl.scala 422:92:@16752.4]
  assign _T_1147 = _T_743 | _T_1146; // @[NV_NVDLA_CSC_wl.scala 422:51:@16753.4]
  assign _T_1148 = _T_1096 & _T_742; // @[NV_NVDLA_CSC_wl.scala 424:40:@16754.4]
  assign _T_1149 = _T_743 | _T_1148; // @[NV_NVDLA_CSC_wl.scala 424:19:@16755.4]
  assign _T_1170 = _T_1163[63:0]; // @[NV_NVDLA_CSC_wl.scala 437:63:@16771.4]
  assign _T_1171 = {{127'd0}, _T_1170}; // @[NV_NVDLA_CSC_wl.scala 437:45:@16772.4]
  assign _T_1172 = ~ _T_742; // @[NV_NVDLA_CSC_wl.scala 437:108:@16773.4]
  assign _T_1176 = _T_1172 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12:@16775.4]
  assign _GEN_503 = {{127'd0}, _T_1176}; // @[NV_NVDLA_CSC_wl.scala 437:85:@16776.4]
  assign _T_1177 = _T_1171 | _GEN_503; // @[NV_NVDLA_CSC_wl.scala 437:85:@16776.4]
  assign _T_1183 = 319'hffffffffffffffff << _T_1118; // @[NV_NVDLA_CSC_wl.scala 438:56:@16778.4]
  assign _T_1184 = ~ _T_1183; // @[NV_NVDLA_CSC_wl.scala 438:25:@16779.4]
  assign _T_1185 = _T_1177[63:0]; // @[NV_NVDLA_CSC_wl.scala 439:41:@16780.4]
  assign _GEN_504 = {{255'd0}, _T_1185}; // @[NV_NVDLA_CSC_wl.scala 439:63:@16781.4]
  assign _T_1186 = _GEN_504 & _T_1184; // @[NV_NVDLA_CSC_wl.scala 439:63:@16781.4]
  assign _GEN_38 = _T_1096 ? _T_1186 : _T_1156; // @[NV_NVDLA_CSC_wl.scala 441:28:@16782.4]
  assign _T_1199 = _T_1163 >> _T_1118; // @[NV_NVDLA_CSC_wl.scala 450:49:@16792.4]
  assign _T_1208 = _T_1138 ? _T_1193 : _T_1199; // @[NV_NVDLA_CSC_wl.scala 453:84:@16797.4]
  assign _T_1209 = _T_743 ? 512'h0 : _T_1208; // @[NV_NVDLA_CSC_wl.scala 453:33:@16798.4]
  assign _T_1215 = _T_1117[4:0]; // @[NV_NVDLA_CSC_wl.scala 456:52:@16804.4]
  assign _T_1217 = {_T_1215,1'h0}; // @[Cat.scala 30:58:@16805.4]
  assign _GEN_506 = {{1'd0}, _T_1215}; // @[NV_NVDLA_CSC_wl.scala 456:69:@16807.4]
  assign _T_1219 = _T_1217 + _GEN_506; // @[NV_NVDLA_CSC_wl.scala 456:69:@16807.4]
  assign _T_1220 = _T_1217 + _GEN_506; // @[NV_NVDLA_CSC_wl.scala 456:69:@16808.4]
  assign _GEN_39 = _T_1149 ? _T_1209 : _T_1163; // @[NV_NVDLA_CSC_wl.scala 458:34:@16809.4]
  assign _GEN_40 = _T_1147 ? _T_1209 : _T_1193; // @[NV_NVDLA_CSC_wl.scala 461:39:@16812.4]
  assign _GEN_41 = _T_1096 ? _T_1117 : _T_1226; // @[NV_NVDLA_CSC_wl.scala 477:28:@16825.4]
  assign _GEN_42 = _T_1096 ? _T_1120 : _T_1229; // @[NV_NVDLA_CSC_wl.scala 477:28:@16825.4]
  assign _GEN_43 = _T_1096 ? _T_1121 : _T_1232; // @[NV_NVDLA_CSC_wl.scala 477:28:@16825.4]
  assign _GEN_44 = _T_1096 ? _T_1122 : _T_1235; // @[NV_NVDLA_CSC_wl.scala 477:28:@16825.4]
  assign _GEN_45 = _T_1096 ? _T_1123 : _T_1238; // @[NV_NVDLA_CSC_wl.scala 477:28:@16825.4]
  assign _GEN_46 = _T_1096 ? _T_1119 : _T_1241; // @[NV_NVDLA_CSC_wl.scala 477:28:@16825.4]
  assign _GEN_47 = _T_1096 ? _T_1124 : _T_1244; // @[NV_NVDLA_CSC_wl.scala 477:28:@16825.4]
  assign _GEN_48 = _T_1096 ? {{1'd0}, _T_1220} : _T_1247; // @[NV_NVDLA_CSC_wl.scala 477:28:@16825.4]
  assign _T_1318 = _T_1156[0]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16836.4]
  assign _T_1319 = _T_1156[1]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16838.4]
  assign _T_1320 = _T_1156[2]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16840.4]
  assign _T_1321 = _T_1156[3]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16842.4]
  assign _T_1322 = _T_1156[4]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16844.4]
  assign _T_1323 = _T_1156[5]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16846.4]
  assign _T_1324 = _T_1156[6]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16848.4]
  assign _T_1325 = _T_1156[7]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16850.4]
  assign _T_1326 = _T_1156[8]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16852.4]
  assign _T_1327 = _T_1156[9]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16854.4]
  assign _T_1328 = _T_1156[10]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16856.4]
  assign _T_1329 = _T_1156[11]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16858.4]
  assign _T_1330 = _T_1156[12]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16860.4]
  assign _T_1331 = _T_1156[13]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16862.4]
  assign _T_1332 = _T_1156[14]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16864.4]
  assign _T_1333 = _T_1156[15]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16866.4]
  assign _T_1334 = _T_1156[16]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16868.4]
  assign _T_1335 = _T_1156[17]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16870.4]
  assign _T_1336 = _T_1156[18]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16872.4]
  assign _T_1337 = _T_1156[19]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16874.4]
  assign _T_1338 = _T_1156[20]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16876.4]
  assign _T_1339 = _T_1156[21]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16878.4]
  assign _T_1340 = _T_1156[22]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16880.4]
  assign _T_1341 = _T_1156[23]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16882.4]
  assign _T_1342 = _T_1156[24]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16884.4]
  assign _T_1343 = _T_1156[25]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16886.4]
  assign _T_1344 = _T_1156[26]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16888.4]
  assign _T_1345 = _T_1156[27]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16890.4]
  assign _T_1346 = _T_1156[28]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16892.4]
  assign _T_1347 = _T_1156[29]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16894.4]
  assign _T_1348 = _T_1156[30]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16896.4]
  assign _T_1349 = _T_1156[31]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16898.4]
  assign _T_1350 = _T_1156[32]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16900.4]
  assign _T_1351 = _T_1156[33]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16902.4]
  assign _T_1352 = _T_1156[34]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16904.4]
  assign _T_1353 = _T_1156[35]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16906.4]
  assign _T_1354 = _T_1156[36]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16908.4]
  assign _T_1355 = _T_1156[37]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16910.4]
  assign _T_1356 = _T_1156[38]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16912.4]
  assign _T_1357 = _T_1156[39]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16914.4]
  assign _T_1358 = _T_1156[40]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16916.4]
  assign _T_1359 = _T_1156[41]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16918.4]
  assign _T_1360 = _T_1156[42]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16920.4]
  assign _T_1361 = _T_1156[43]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16922.4]
  assign _T_1362 = _T_1156[44]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16924.4]
  assign _T_1363 = _T_1156[45]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16926.4]
  assign _T_1364 = _T_1156[46]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16928.4]
  assign _T_1365 = _T_1156[47]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16930.4]
  assign _T_1366 = _T_1156[48]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16932.4]
  assign _T_1367 = _T_1156[49]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16934.4]
  assign _T_1368 = _T_1156[50]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16936.4]
  assign _T_1369 = _T_1156[51]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16938.4]
  assign _T_1370 = _T_1156[52]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16940.4]
  assign _T_1371 = _T_1156[53]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16942.4]
  assign _T_1372 = _T_1156[54]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16944.4]
  assign _T_1373 = _T_1156[55]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16946.4]
  assign _T_1374 = _T_1156[56]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16948.4]
  assign _T_1375 = _T_1156[57]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16950.4]
  assign _T_1376 = _T_1156[58]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16952.4]
  assign _T_1377 = _T_1156[59]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16954.4]
  assign _T_1378 = _T_1156[60]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16956.4]
  assign _T_1379 = _T_1156[61]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16958.4]
  assign _T_1380 = _T_1156[62]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16960.4]
  assign _T_1381 = _T_1156[63]; // @[NV_NVDLA_CSC_wl.scala 497:40:@16962.4]
  assign _T_1382 = _T_1318 + _T_1319; // @[NV_NVDLA_CSC_wl.scala 499:46:@16964.4]
  assign _GEN_507 = {{1'd0}, _T_1320}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16965.4]
  assign _T_1383 = _T_1382 + _GEN_507; // @[NV_NVDLA_CSC_wl.scala 499:46:@16965.4]
  assign _GEN_508 = {{2'd0}, _T_1321}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16966.4]
  assign _T_1384 = _T_1383 + _GEN_508; // @[NV_NVDLA_CSC_wl.scala 499:46:@16966.4]
  assign _GEN_509 = {{3'd0}, _T_1322}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16967.4]
  assign _T_1385 = _T_1384 + _GEN_509; // @[NV_NVDLA_CSC_wl.scala 499:46:@16967.4]
  assign _GEN_510 = {{4'd0}, _T_1323}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16968.4]
  assign _T_1386 = _T_1385 + _GEN_510; // @[NV_NVDLA_CSC_wl.scala 499:46:@16968.4]
  assign _GEN_511 = {{5'd0}, _T_1324}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16969.4]
  assign _T_1387 = _T_1386 + _GEN_511; // @[NV_NVDLA_CSC_wl.scala 499:46:@16969.4]
  assign _GEN_512 = {{6'd0}, _T_1325}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16970.4]
  assign _T_1388 = _T_1387 + _GEN_512; // @[NV_NVDLA_CSC_wl.scala 499:46:@16970.4]
  assign _GEN_513 = {{7'd0}, _T_1326}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16971.4]
  assign _T_1389 = _T_1388 + _GEN_513; // @[NV_NVDLA_CSC_wl.scala 499:46:@16971.4]
  assign _GEN_514 = {{8'd0}, _T_1327}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16972.4]
  assign _T_1390 = _T_1389 + _GEN_514; // @[NV_NVDLA_CSC_wl.scala 499:46:@16972.4]
  assign _GEN_515 = {{9'd0}, _T_1328}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16973.4]
  assign _T_1391 = _T_1390 + _GEN_515; // @[NV_NVDLA_CSC_wl.scala 499:46:@16973.4]
  assign _GEN_516 = {{10'd0}, _T_1329}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16974.4]
  assign _T_1392 = _T_1391 + _GEN_516; // @[NV_NVDLA_CSC_wl.scala 499:46:@16974.4]
  assign _GEN_517 = {{11'd0}, _T_1330}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16975.4]
  assign _T_1393 = _T_1392 + _GEN_517; // @[NV_NVDLA_CSC_wl.scala 499:46:@16975.4]
  assign _GEN_518 = {{12'd0}, _T_1331}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16976.4]
  assign _T_1394 = _T_1393 + _GEN_518; // @[NV_NVDLA_CSC_wl.scala 499:46:@16976.4]
  assign _GEN_519 = {{13'd0}, _T_1332}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16977.4]
  assign _T_1395 = _T_1394 + _GEN_519; // @[NV_NVDLA_CSC_wl.scala 499:46:@16977.4]
  assign _GEN_520 = {{14'd0}, _T_1333}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16978.4]
  assign _T_1396 = _T_1395 + _GEN_520; // @[NV_NVDLA_CSC_wl.scala 499:46:@16978.4]
  assign _GEN_521 = {{15'd0}, _T_1334}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16979.4]
  assign _T_1397 = _T_1396 + _GEN_521; // @[NV_NVDLA_CSC_wl.scala 499:46:@16979.4]
  assign _GEN_522 = {{16'd0}, _T_1335}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16980.4]
  assign _T_1398 = _T_1397 + _GEN_522; // @[NV_NVDLA_CSC_wl.scala 499:46:@16980.4]
  assign _GEN_523 = {{17'd0}, _T_1336}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16981.4]
  assign _T_1399 = _T_1398 + _GEN_523; // @[NV_NVDLA_CSC_wl.scala 499:46:@16981.4]
  assign _GEN_524 = {{18'd0}, _T_1337}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16982.4]
  assign _T_1400 = _T_1399 + _GEN_524; // @[NV_NVDLA_CSC_wl.scala 499:46:@16982.4]
  assign _GEN_525 = {{19'd0}, _T_1338}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16983.4]
  assign _T_1401 = _T_1400 + _GEN_525; // @[NV_NVDLA_CSC_wl.scala 499:46:@16983.4]
  assign _GEN_526 = {{20'd0}, _T_1339}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16984.4]
  assign _T_1402 = _T_1401 + _GEN_526; // @[NV_NVDLA_CSC_wl.scala 499:46:@16984.4]
  assign _GEN_527 = {{21'd0}, _T_1340}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16985.4]
  assign _T_1403 = _T_1402 + _GEN_527; // @[NV_NVDLA_CSC_wl.scala 499:46:@16985.4]
  assign _GEN_528 = {{22'd0}, _T_1341}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16986.4]
  assign _T_1404 = _T_1403 + _GEN_528; // @[NV_NVDLA_CSC_wl.scala 499:46:@16986.4]
  assign _GEN_529 = {{23'd0}, _T_1342}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16987.4]
  assign _T_1405 = _T_1404 + _GEN_529; // @[NV_NVDLA_CSC_wl.scala 499:46:@16987.4]
  assign _GEN_530 = {{24'd0}, _T_1343}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16988.4]
  assign _T_1406 = _T_1405 + _GEN_530; // @[NV_NVDLA_CSC_wl.scala 499:46:@16988.4]
  assign _GEN_531 = {{25'd0}, _T_1344}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16989.4]
  assign _T_1407 = _T_1406 + _GEN_531; // @[NV_NVDLA_CSC_wl.scala 499:46:@16989.4]
  assign _GEN_532 = {{26'd0}, _T_1345}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16990.4]
  assign _T_1408 = _T_1407 + _GEN_532; // @[NV_NVDLA_CSC_wl.scala 499:46:@16990.4]
  assign _GEN_533 = {{27'd0}, _T_1346}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16991.4]
  assign _T_1409 = _T_1408 + _GEN_533; // @[NV_NVDLA_CSC_wl.scala 499:46:@16991.4]
  assign _GEN_534 = {{28'd0}, _T_1347}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16992.4]
  assign _T_1410 = _T_1409 + _GEN_534; // @[NV_NVDLA_CSC_wl.scala 499:46:@16992.4]
  assign _GEN_535 = {{29'd0}, _T_1348}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16993.4]
  assign _T_1411 = _T_1410 + _GEN_535; // @[NV_NVDLA_CSC_wl.scala 499:46:@16993.4]
  assign _GEN_536 = {{30'd0}, _T_1349}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16994.4]
  assign _T_1412 = _T_1411 + _GEN_536; // @[NV_NVDLA_CSC_wl.scala 499:46:@16994.4]
  assign _GEN_537 = {{31'd0}, _T_1350}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16995.4]
  assign _T_1413 = _T_1412 + _GEN_537; // @[NV_NVDLA_CSC_wl.scala 499:46:@16995.4]
  assign _GEN_538 = {{32'd0}, _T_1351}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16996.4]
  assign _T_1414 = _T_1413 + _GEN_538; // @[NV_NVDLA_CSC_wl.scala 499:46:@16996.4]
  assign _GEN_539 = {{33'd0}, _T_1352}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16997.4]
  assign _T_1415 = _T_1414 + _GEN_539; // @[NV_NVDLA_CSC_wl.scala 499:46:@16997.4]
  assign _GEN_540 = {{34'd0}, _T_1353}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16998.4]
  assign _T_1416 = _T_1415 + _GEN_540; // @[NV_NVDLA_CSC_wl.scala 499:46:@16998.4]
  assign _GEN_541 = {{35'd0}, _T_1354}; // @[NV_NVDLA_CSC_wl.scala 499:46:@16999.4]
  assign _T_1417 = _T_1416 + _GEN_541; // @[NV_NVDLA_CSC_wl.scala 499:46:@16999.4]
  assign _GEN_542 = {{36'd0}, _T_1355}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17000.4]
  assign _T_1418 = _T_1417 + _GEN_542; // @[NV_NVDLA_CSC_wl.scala 499:46:@17000.4]
  assign _GEN_543 = {{37'd0}, _T_1356}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17001.4]
  assign _T_1419 = _T_1418 + _GEN_543; // @[NV_NVDLA_CSC_wl.scala 499:46:@17001.4]
  assign _GEN_544 = {{38'd0}, _T_1357}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17002.4]
  assign _T_1420 = _T_1419 + _GEN_544; // @[NV_NVDLA_CSC_wl.scala 499:46:@17002.4]
  assign _GEN_545 = {{39'd0}, _T_1358}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17003.4]
  assign _T_1421 = _T_1420 + _GEN_545; // @[NV_NVDLA_CSC_wl.scala 499:46:@17003.4]
  assign _GEN_546 = {{40'd0}, _T_1359}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17004.4]
  assign _T_1422 = _T_1421 + _GEN_546; // @[NV_NVDLA_CSC_wl.scala 499:46:@17004.4]
  assign _GEN_547 = {{41'd0}, _T_1360}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17005.4]
  assign _T_1423 = _T_1422 + _GEN_547; // @[NV_NVDLA_CSC_wl.scala 499:46:@17005.4]
  assign _GEN_548 = {{42'd0}, _T_1361}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17006.4]
  assign _T_1424 = _T_1423 + _GEN_548; // @[NV_NVDLA_CSC_wl.scala 499:46:@17006.4]
  assign _GEN_549 = {{43'd0}, _T_1362}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17007.4]
  assign _T_1425 = _T_1424 + _GEN_549; // @[NV_NVDLA_CSC_wl.scala 499:46:@17007.4]
  assign _GEN_550 = {{44'd0}, _T_1363}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17008.4]
  assign _T_1426 = _T_1425 + _GEN_550; // @[NV_NVDLA_CSC_wl.scala 499:46:@17008.4]
  assign _GEN_551 = {{45'd0}, _T_1364}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17009.4]
  assign _T_1427 = _T_1426 + _GEN_551; // @[NV_NVDLA_CSC_wl.scala 499:46:@17009.4]
  assign _GEN_552 = {{46'd0}, _T_1365}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17010.4]
  assign _T_1428 = _T_1427 + _GEN_552; // @[NV_NVDLA_CSC_wl.scala 499:46:@17010.4]
  assign _GEN_553 = {{47'd0}, _T_1366}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17011.4]
  assign _T_1429 = _T_1428 + _GEN_553; // @[NV_NVDLA_CSC_wl.scala 499:46:@17011.4]
  assign _GEN_554 = {{48'd0}, _T_1367}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17012.4]
  assign _T_1430 = _T_1429 + _GEN_554; // @[NV_NVDLA_CSC_wl.scala 499:46:@17012.4]
  assign _GEN_555 = {{49'd0}, _T_1368}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17013.4]
  assign _T_1431 = _T_1430 + _GEN_555; // @[NV_NVDLA_CSC_wl.scala 499:46:@17013.4]
  assign _GEN_556 = {{50'd0}, _T_1369}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17014.4]
  assign _T_1432 = _T_1431 + _GEN_556; // @[NV_NVDLA_CSC_wl.scala 499:46:@17014.4]
  assign _GEN_557 = {{51'd0}, _T_1370}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17015.4]
  assign _T_1433 = _T_1432 + _GEN_557; // @[NV_NVDLA_CSC_wl.scala 499:46:@17015.4]
  assign _GEN_558 = {{52'd0}, _T_1371}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17016.4]
  assign _T_1434 = _T_1433 + _GEN_558; // @[NV_NVDLA_CSC_wl.scala 499:46:@17016.4]
  assign _GEN_559 = {{53'd0}, _T_1372}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17017.4]
  assign _T_1435 = _T_1434 + _GEN_559; // @[NV_NVDLA_CSC_wl.scala 499:46:@17017.4]
  assign _GEN_560 = {{54'd0}, _T_1373}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17018.4]
  assign _T_1436 = _T_1435 + _GEN_560; // @[NV_NVDLA_CSC_wl.scala 499:46:@17018.4]
  assign _GEN_561 = {{55'd0}, _T_1374}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17019.4]
  assign _T_1437 = _T_1436 + _GEN_561; // @[NV_NVDLA_CSC_wl.scala 499:46:@17019.4]
  assign _GEN_562 = {{56'd0}, _T_1375}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17020.4]
  assign _T_1438 = _T_1437 + _GEN_562; // @[NV_NVDLA_CSC_wl.scala 499:46:@17020.4]
  assign _GEN_563 = {{57'd0}, _T_1376}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17021.4]
  assign _T_1439 = _T_1438 + _GEN_563; // @[NV_NVDLA_CSC_wl.scala 499:46:@17021.4]
  assign _GEN_564 = {{58'd0}, _T_1377}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17022.4]
  assign _T_1440 = _T_1439 + _GEN_564; // @[NV_NVDLA_CSC_wl.scala 499:46:@17022.4]
  assign _GEN_565 = {{59'd0}, _T_1378}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17023.4]
  assign _T_1441 = _T_1440 + _GEN_565; // @[NV_NVDLA_CSC_wl.scala 499:46:@17023.4]
  assign _GEN_566 = {{60'd0}, _T_1379}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17024.4]
  assign _T_1442 = _T_1441 + _GEN_566; // @[NV_NVDLA_CSC_wl.scala 499:46:@17024.4]
  assign _GEN_567 = {{61'd0}, _T_1380}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17025.4]
  assign _T_1443 = _T_1442 + _GEN_567; // @[NV_NVDLA_CSC_wl.scala 499:46:@17025.4]
  assign _GEN_568 = {{62'd0}, _T_1381}; // @[NV_NVDLA_CSC_wl.scala 499:46:@17026.4]
  assign _T_1444 = _T_1443 + _GEN_568; // @[NV_NVDLA_CSC_wl.scala 499:46:@17026.4]
  assign _T_1453 = 191'hffffffffffffffff << _T_1226; // @[NV_NVDLA_CSC_wl.scala 505:57:@17029.4]
  assign _T_1454 = ~ _T_1453; // @[NV_NVDLA_CSC_wl.scala 505:26:@17030.4]
  assign _T_1456 = _T_1244 >= 2'h1; // @[NV_NVDLA_CSC_wl.scala 508:45:@17031.4]
  assign _T_1467 = _T_1456 ? 64'hffffffffffffffff : 64'h0; // @[NV_NVDLA_CSC_wl.scala 508:27:@17034.4]
  assign _T_1469 = _T_1244 >= 2'h2; // @[NV_NVDLA_CSC_wl.scala 509:45:@17035.4]
  assign _T_1480 = _T_1469 ? 64'hffffffffffffffff : 64'h0; // @[NV_NVDLA_CSC_wl.scala 509:27:@17038.4]
  assign _T_1482 = _T_1244 >= 2'h3; // @[NV_NVDLA_CSC_wl.scala 510:45:@17039.4]
  assign _T_1493 = _T_1482 ? 64'hffffffffffffffff : 64'h0; // @[NV_NVDLA_CSC_wl.scala 510:27:@17042.4]
  assign _T_1494 = _T_1226[5:0]; // @[NV_NVDLA_CSC_wl.scala 514:50:@17043.4]
  assign _T_1496 = {_T_1494,1'h0}; // @[Cat.scala 30:58:@17044.4]
  assign _T_1497 = _T_1156[63:0]; // @[NV_NVDLA_CSC_wl.scala 515:39:@17045.4]
  assign _GEN_569 = {{127'd0}, _T_1497}; // @[NV_NVDLA_CSC_wl.scala 515:61:@17046.4]
  assign _T_1498 = _GEN_569 & _T_1454; // @[NV_NVDLA_CSC_wl.scala 515:61:@17046.4]
  assign _T_1500 = _T_1497 >> _T_1226; // @[NV_NVDLA_CSC_wl.scala 516:62:@17048.4]
  assign _GEN_570 = {{127'd0}, _T_1500}; // @[NV_NVDLA_CSC_wl.scala 516:83:@17049.4]
  assign _T_1501 = _GEN_570 & _T_1454; // @[NV_NVDLA_CSC_wl.scala 516:83:@17049.4]
  assign _GEN_571 = {{127'd0}, _T_1467}; // @[NV_NVDLA_CSC_wl.scala 516:100:@17050.4]
  assign _T_1502 = _T_1501 & _GEN_571; // @[NV_NVDLA_CSC_wl.scala 516:100:@17050.4]
  assign _T_1504 = _T_1497 >> _T_1496; // @[NV_NVDLA_CSC_wl.scala 517:62:@17052.4]
  assign _GEN_572 = {{127'd0}, _T_1504}; // @[NV_NVDLA_CSC_wl.scala 517:83:@17053.4]
  assign _T_1505 = _GEN_572 & _T_1454; // @[NV_NVDLA_CSC_wl.scala 517:83:@17053.4]
  assign _GEN_573 = {{127'd0}, _T_1480}; // @[NV_NVDLA_CSC_wl.scala 517:100:@17054.4]
  assign _T_1506 = _T_1505 & _GEN_573; // @[NV_NVDLA_CSC_wl.scala 517:100:@17054.4]
  assign _T_1508 = _T_1497 >> _T_1247; // @[NV_NVDLA_CSC_wl.scala 518:62:@17056.4]
  assign _GEN_574 = {{127'd0}, _T_1508}; // @[NV_NVDLA_CSC_wl.scala 518:83:@17057.4]
  assign _T_1509 = _GEN_574 & _T_1454; // @[NV_NVDLA_CSC_wl.scala 518:83:@17057.4]
  assign _GEN_575 = {{127'd0}, _T_1493}; // @[NV_NVDLA_CSC_wl.scala 518:100:@17058.4]
  assign _T_1510 = _T_1509 & _GEN_575; // @[NV_NVDLA_CSC_wl.scala 518:100:@17058.4]
  assign _T_1517 = _T_739 == 3'h1; // @[NV_NVDLA_CSC_wl.scala 523:41:@17060.4]
  assign _T_1519 = _T_739 == 3'h2; // @[NV_NVDLA_CSC_wl.scala 524:41:@17061.4]
  assign _T_1520 = _T_1502[31:0]; // @[NV_NVDLA_CSC_wl.scala 524:82:@17062.4]
  assign _T_1521 = _T_1498[31:0]; // @[NV_NVDLA_CSC_wl.scala 524:122:@17063.4]
  assign _T_1522 = {_T_1520,_T_1521}; // @[Cat.scala 30:58:@17064.4]
  assign _T_1523 = _T_1510[15:0]; // @[NV_NVDLA_CSC_wl.scala 525:44:@17065.4]
  assign _T_1524 = _T_1506[15:0]; // @[NV_NVDLA_CSC_wl.scala 525:84:@17066.4]
  assign _T_1525 = _T_1502[15:0]; // @[NV_NVDLA_CSC_wl.scala 525:124:@17067.4]
  assign _T_1526 = _T_1498[15:0]; // @[NV_NVDLA_CSC_wl.scala 525:164:@17068.4]
  assign _T_1529 = {_T_1523,_T_1524,_T_1525,_T_1526}; // @[Cat.scala 30:58:@17071.4]
  assign _T_1530 = _T_1519 ? _T_1522 : _T_1529; // @[NV_NVDLA_CSC_wl.scala 524:28:@17072.4]
  assign _T_1531 = _T_1517 ? _T_1498 : {{127'd0}, _T_1530}; // @[NV_NVDLA_CSC_wl.scala 523:28:@17073.4]
  assign _T_1532 = _T_743 ? 191'h0 : _T_1531; // @[NV_NVDLA_CSC_wl.scala 522:28:@17074.4]
  assign _GEN_576 = {{127'd0}, _T_1447}; // @[NV_NVDLA_CSC_wl.scala 528:61:@17075.4]
  assign _T_1533 = _T_1532 != _GEN_576; // @[NV_NVDLA_CSC_wl.scala 528:61:@17075.4]
  assign _T_1534 = _T_1223 & _T_1533; // @[NV_NVDLA_CSC_wl.scala 528:44:@17076.4]
  assign _GEN_577 = {{56'd0}, _T_1537}; // @[NV_NVDLA_CSC_wl.scala 534:57:@17079.4]
  assign _T_1541 = _GEN_577 < _T_1444; // @[NV_NVDLA_CSC_wl.scala 534:57:@17079.4]
  assign _T_1542 = _T_1223 & _T_1541; // @[NV_NVDLA_CSC_wl.scala 534:42:@17080.4]
  assign _T_1543 = ~ _T_1542; // @[NV_NVDLA_CSC_wl.scala 536:31:@17081.4]
  assign _T_1546 = _T_1543 ? 8'h0 : 8'h40; // @[NV_NVDLA_CSC_wl.scala 536:30:@17082.4]
  assign _T_1547 = _T_1537 + _T_1546; // @[NV_NVDLA_CSC_wl.scala 538:39:@17083.4]
  assign _T_1548 = _T_1537 + _T_1546; // @[NV_NVDLA_CSC_wl.scala 538:39:@17084.4]
  assign _GEN_578 = {{56'd0}, _T_1548}; // @[NV_NVDLA_CSC_wl.scala 538:57:@17085.4]
  assign _T_1549 = _GEN_578 - _T_1444; // @[NV_NVDLA_CSC_wl.scala 538:57:@17085.4]
  assign _T_1550 = $unsigned(_T_1549); // @[NV_NVDLA_CSC_wl.scala 538:57:@17086.4]
  assign _T_1551 = _T_1550[63:0]; // @[NV_NVDLA_CSC_wl.scala 538:57:@17087.4]
  assign _T_1553 = ~ _T_1235; // @[NV_NVDLA_CSC_wl.scala 540:29:@17088.4]
  assign _T_1554 = _T_1553 & _T_1232; // @[NV_NVDLA_CSC_wl.scala 540:47:@17089.4]
  assign _T_1555 = _T_1554 ? {{56'd0}, _T_1540} : _T_1551; // @[NV_NVDLA_CSC_wl.scala 540:28:@17090.4]
  assign _T_1556 = _T_743 ? 64'h0 : _T_1555; // @[NV_NVDLA_CSC_wl.scala 539:28:@17091.4]
  assign _T_1557 = _T_1223 & _T_1229; // @[NV_NVDLA_CSC_wl.scala 543:61:@17092.4]
  assign _T_1558 = _T_1557 & _T_1235; // @[NV_NVDLA_CSC_wl.scala 543:81:@17093.4]
  assign _T_1559 = _T_743 | _T_1558; // @[NV_NVDLA_CSC_wl.scala 543:40:@17094.4]
  assign _T_1560 = _T_743 | _T_1223; // @[NV_NVDLA_CSC_wl.scala 545:19:@17095.4]
  assign _GEN_49 = _T_1560 ? _T_1556 : {{56'd0}, _T_1537}; // @[NV_NVDLA_CSC_wl.scala 545:39:@17096.4]
  assign _GEN_50 = _T_1559 ? _T_1556 : {{56'd0}, _T_1540}; // @[NV_NVDLA_CSC_wl.scala 548:30:@17099.4]
  assign _T_1568 = _T_1563 + 13'h1; // @[NV_NVDLA_CSC_wl.scala 556:39:@17104.4]
  assign _T_1569 = _T_1563 + 13'h1; // @[NV_NVDLA_CSC_wl.scala 556:39:@17105.4]
  assign _GEN_579 = {{1'd0}, _T_1569}; // @[NV_NVDLA_CSC_wl.scala 557:48:@17108.4]
  assign _T_1576 = _GEN_579 == _T_802; // @[NV_NVDLA_CSC_wl.scala 557:48:@17108.4]
  assign _T_1582 = _T_1576 ? 13'h0 : _T_1569; // @[NV_NVDLA_CSC_wl.scala 558:35:@17110.4]
  assign _T_1583 = _T_813[12:0]; // @[NV_NVDLA_CSC_wl.scala 560:53:@17111.4]
  assign _T_1586 = _T_1542 ? _T_1582 : _T_1563; // @[NV_NVDLA_CSC_wl.scala 562:28:@17114.4]
  assign _T_1587 = _T_1554 ? _T_1566 : _T_1586; // @[NV_NVDLA_CSC_wl.scala 561:28:@17115.4]
  assign _T_1588 = _T_708 ? _T_1583 : _T_1587; // @[NV_NVDLA_CSC_wl.scala 560:28:@17116.4]
  assign _T_1589 = _T_708 | _T_1542; // @[NV_NVDLA_CSC_wl.scala 566:40:@17117.4]
  assign _T_1590 = _T_1223 & _T_1232; // @[NV_NVDLA_CSC_wl.scala 566:76:@17118.4]
  assign _T_1591 = _T_1589 | _T_1590; // @[NV_NVDLA_CSC_wl.scala 566:55:@17119.4]
  assign _T_1592 = _T_1223 & _T_1223; // @[NV_NVDLA_CSC_wl.scala 567:66:@17120.4]
  assign _T_1593 = _T_1592 & _T_1235; // @[NV_NVDLA_CSC_wl.scala 567:86:@17121.4]
  assign _T_1594 = _T_708 | _T_1593; // @[NV_NVDLA_CSC_wl.scala 567:45:@17122.4]
  assign _T_1600 = {_T_715,9'h0}; // @[Cat.scala 30:58:@17124.4]
  assign _GEN_580 = {{1'd0}, _T_1563}; // @[NV_NVDLA_CSC_wl.scala 568:39:@17125.4]
  assign _T_1601 = _GEN_580 + _T_1600; // @[NV_NVDLA_CSC_wl.scala 568:39:@17125.4]
  assign _T_1602 = _GEN_580 + _T_1600; // @[NV_NVDLA_CSC_wl.scala 568:39:@17126.4]
  assign _GEN_51 = _T_1591 ? _T_1588 : _T_1563; // @[NV_NVDLA_CSC_wl.scala 570:29:@17127.4]
  assign _GEN_52 = _T_1594 ? _T_1588 : _T_1566; // @[NV_NVDLA_CSC_wl.scala 573:34:@17130.4]
  assign _T_1609 = _T_743 | _T_1235; // @[NV_NVDLA_CSC_wl.scala 581:42:@17135.4]
  assign _T_1612 = _T_1232 ? 1'h1 : _T_1605; // @[NV_NVDLA_CSC_wl.scala 581:76:@17136.4]
  assign _T_1613 = _T_1609 ? 1'h0 : _T_1612; // @[NV_NVDLA_CSC_wl.scala 581:31:@17137.4]
  assign _T_1615 = _T_1608 + 15'h1; // @[NV_NVDLA_CSC_wl.scala 582:37:@17138.4]
  assign _T_1616 = _T_1608 + 15'h1; // @[NV_NVDLA_CSC_wl.scala 582:37:@17139.4]
  assign _T_1619 = _T_1235 ? 15'h0 : _T_1616; // @[NV_NVDLA_CSC_wl.scala 583:84:@17140.4]
  assign _T_1620 = _T_743 ? 15'h0 : _T_1619; // @[NV_NVDLA_CSC_wl.scala 583:27:@17141.4]
  assign _T_1621 = _T_1223 & _T_1235; // @[NV_NVDLA_CSC_wl.scala 584:59:@17142.4]
  assign _T_1622 = _T_743 | _T_1621; // @[NV_NVDLA_CSC_wl.scala 584:38:@17143.4]
  assign _T_1623 = ~ _T_1605; // @[NV_NVDLA_CSC_wl.scala 584:82:@17144.4]
  assign _T_1624 = _T_1623 & _T_1542; // @[NV_NVDLA_CSC_wl.scala 584:98:@17145.4]
  assign _T_1625 = _T_1622 | _T_1624; // @[NV_NVDLA_CSC_wl.scala 584:79:@17146.4]
  assign _T_1627 = _T_1605 | _T_1543; // @[NV_NVDLA_CSC_wl.scala 585:45:@17148.4]
  assign _T_1628 = _T_1627 ? _T_1608 : _T_1616; // @[NV_NVDLA_CSC_wl.scala 585:29:@17149.4]
  assign _GEN_53 = _T_1625 ? _T_1620 : _T_1608; // @[NV_NVDLA_CSC_wl.scala 588:28:@17151.4]
  assign _GEN_54 = _T_1542 ? _T_1602 : {{1'd0}, _T_1634}; // @[NV_NVDLA_CSC_wl.scala 609:23:@17166.4]
  assign _GEN_55 = _T_1223 ? _T_1229 : _T_1640; // @[NV_NVDLA_CSC_wl.scala 613:28:@17170.4]
  assign _GEN_56 = _T_1223 ? _T_1232 : _T_1643; // @[NV_NVDLA_CSC_wl.scala 613:28:@17170.4]
  assign _GEN_57 = _T_1223 ? _T_1235 : _T_1646; // @[NV_NVDLA_CSC_wl.scala 613:28:@17170.4]
  assign _GEN_58 = _T_1223 ? _T_1238 : _T_1649; // @[NV_NVDLA_CSC_wl.scala 613:28:@17170.4]
  assign _GEN_59 = _T_1223 ? _T_1444 : {{56'd0}, _T_1652}; // @[NV_NVDLA_CSC_wl.scala 613:28:@17170.4]
  assign _GEN_60 = _T_1560 ? _T_1532 : {{127'd0}, _T_1447}; // @[NV_NVDLA_CSC_wl.scala 621:39:@17178.4]
  assign _GEN_61 = _T_1223 ? _T_1241 : _T_1658; // @[NV_NVDLA_CSC_wl.scala 625:28:@17182.4]
  assign _T_1663 = _T_1223 & _T_1238; // @[NV_NVDLA_CSC_wl.scala 628:28:@17185.4]
  assign _GEN_62 = _T_1663 ? _T_1628 : _T_1661; // @[NV_NVDLA_CSC_wl.scala 628:41:@17186.4]
  assign _T_1672 = {_T_1649,_T_1646,_T_1643,_T_1640,_T_1661,_T_1658,_T_1652}; // @[Cat.scala 30:58:@17199.4]
  assign _GEN_63 = _T_1637 ? _T_1672 : _T_1697; // @[NV_NVDLA_CSC_wl.scala 669:36:@17233.4]
  assign _GEN_64 = _T_1655 ? _T_1447 : _T_1737; // @[NV_NVDLA_CSC_wl.scala 673:34:@17237.4]
  assign _GEN_65 = _T_1677 ? _T_1697 : _T_1700; // @[NV_NVDLA_CSC_wl.scala 669:36:@17241.4]
  assign _GEN_66 = _T_1717 ? _T_1737 : _T_1740; // @[NV_NVDLA_CSC_wl.scala 673:34:@17245.4]
  assign _GEN_67 = _T_1680 ? _T_1700 : _T_1703; // @[NV_NVDLA_CSC_wl.scala 669:36:@17249.4]
  assign _GEN_68 = _T_1720 ? _T_1740 : _T_1743; // @[NV_NVDLA_CSC_wl.scala 673:34:@17253.4]
  assign _GEN_69 = _T_1683 ? _T_1703 : _T_1706; // @[NV_NVDLA_CSC_wl.scala 669:36:@17257.4]
  assign _GEN_70 = _T_1723 ? _T_1743 : _T_1746; // @[NV_NVDLA_CSC_wl.scala 673:34:@17261.4]
  assign _GEN_71 = _T_1686 ? _T_1706 : _T_1709; // @[NV_NVDLA_CSC_wl.scala 669:36:@17265.4]
  assign _GEN_72 = _T_1726 ? _T_1746 : _T_1749; // @[NV_NVDLA_CSC_wl.scala 673:34:@17269.4]
  assign _GEN_73 = _T_1689 ? _T_1709 : _T_1712; // @[NV_NVDLA_CSC_wl.scala 669:36:@17273.4]
  assign _GEN_74 = _T_1729 ? _T_1749 : _T_1752; // @[NV_NVDLA_CSC_wl.scala 673:34:@17277.4]
  assign _T_1753 = _T_1712[7:0]; // @[NV_NVDLA_CSC_wl.scala 687:38:@17281.4]
  assign _T_1756 = _T_1712[32]; // @[NV_NVDLA_CSC_wl.scala 690:44:@17286.4]
  assign _T_1757 = _T_1712[33]; // @[NV_NVDLA_CSC_wl.scala 691:45:@17287.4]
  assign _T_1758 = _T_1712[34]; // @[NV_NVDLA_CSC_wl.scala 692:43:@17288.4]
  assign _T_1768 = io_sc2buf_wt_rd_data_valid ? 8'h40 : 8'h0; // @[NV_NVDLA_CSC_wl.scala 702:37:@17293.4]
  assign _T_1770 = ~ _T_1758; // @[NV_NVDLA_CSC_wl.scala 704:55:@17294.4]
  assign _T_1771 = _T_1757 & _T_1770; // @[NV_NVDLA_CSC_wl.scala 704:53:@17295.4]
  assign _T_1773 = {2'h0,_T_1765}; // @[Cat.scala 30:58:@17296.4]
  assign _GEN_581 = {{1'd0}, _T_1762}; // @[NV_NVDLA_CSC_wl.scala 704:141:@17297.4]
  assign _T_1774 = _GEN_581 + _T_1768; // @[NV_NVDLA_CSC_wl.scala 704:141:@17297.4]
  assign _T_1775 = _GEN_581 + _T_1768; // @[NV_NVDLA_CSC_wl.scala 704:141:@17298.4]
  assign _T_1776 = _T_1775 - _T_1753; // @[NV_NVDLA_CSC_wl.scala 704:166:@17299.4]
  assign _T_1777 = $unsigned(_T_1776); // @[NV_NVDLA_CSC_wl.scala 704:166:@17300.4]
  assign _T_1778 = _T_1777[7:0]; // @[NV_NVDLA_CSC_wl.scala 704:166:@17301.4]
  assign _T_1779 = _T_1771 ? _T_1773 : {{1'd0}, _T_1778}; // @[NV_NVDLA_CSC_wl.scala 704:33:@17302.4]
  assign _T_1780 = _T_743 ? 9'h0 : _T_1779; // @[NV_NVDLA_CSC_wl.scala 703:35:@17303.4]
  assign _T_1781 = _T_1780[6:0]; // @[NV_NVDLA_CSC_wl.scala 704:182:@17304.4]
  assign _T_1782 = _T_743 | _T_1692; // @[NV_NVDLA_CSC_wl.scala 705:42:@17305.4]
  assign _T_1783 = _T_1692 & _T_1758; // @[NV_NVDLA_CSC_wl.scala 706:67:@17306.4]
  assign _T_1784 = _T_743 | _T_1783; // @[NV_NVDLA_CSC_wl.scala 706:47:@17307.4]
  assign _GEN_75 = _T_1782 ? _T_1781 : _T_1762; // @[NV_NVDLA_CSC_wl.scala 708:32:@17308.4]
  assign _GEN_76 = _T_1784 ? _T_1781 : _T_1765; // @[NV_NVDLA_CSC_wl.scala 711:37:@17311.4]
  assign _T_1790 = _T_1753 - _GEN_581; // @[NV_NVDLA_CSC_wl.scala 719:40:@17317.4]
  assign _T_1791 = $unsigned(_T_1790); // @[NV_NVDLA_CSC_wl.scala 719:40:@17318.4]
  assign _T_1792 = _T_1791[7:0]; // @[NV_NVDLA_CSC_wl.scala 719:40:@17319.4]
  assign _T_1795 = {_T_1792,3'h0}; // @[Cat.scala 30:58:@17321.4]
  assign _T_1796 = io_sc2buf_wt_rd_data_bits >> _T_1795; // @[NV_NVDLA_CSC_wl.scala 720:82:@17322.4]
  assign _T_1798 = _T_1762 != 7'h0; // @[NV_NVDLA_CSC_wl.scala 721:58:@17323.4]
  assign _T_1799 = ~ _T_1798; // @[NV_NVDLA_CSC_wl.scala 721:38:@17324.4]
  assign _T_1801 = _T_1799 ? 512'h0 : _T_1786; // @[NV_NVDLA_CSC_wl.scala 721:36:@17325.4]
  assign _T_1803 = {_T_1753,3'h0}; // @[Cat.scala 30:58:@17326.4]
  assign _T_1804 = _T_1786 >> _T_1803; // @[NV_NVDLA_CSC_wl.scala 722:45:@17327.4]
  assign _T_1809 = _T_1765 != 7'h0; // @[NV_NVDLA_CSC_wl.scala 725:98:@17330.4]
  assign _T_1810 = _T_1771 & _T_1809; // @[NV_NVDLA_CSC_wl.scala 725:71:@17331.4]
  assign _T_1811 = io_sc2buf_wt_rd_data_valid ? _T_1796 : _T_1804; // @[NV_NVDLA_CSC_wl.scala 726:31:@17332.4]
  assign _T_1812 = _T_1810 ? _T_1788 : _T_1811; // @[NV_NVDLA_CSC_wl.scala 725:31:@17333.4]
  assign _T_1813 = _T_743 ? 512'h0 : _T_1812; // @[NV_NVDLA_CSC_wl.scala 724:31:@17334.4]
  assign _T_1815 = _T_1781 != 7'h0; // @[NV_NVDLA_CSC_wl.scala 729:86:@17335.4]
  assign _T_1816 = _T_1692 & _T_1815; // @[NV_NVDLA_CSC_wl.scala 729:62:@17336.4]
  assign _T_1817 = _T_743 | _T_1816; // @[NV_NVDLA_CSC_wl.scala 729:42:@17337.4]
  assign _T_1821 = _T_1783 & _T_1815; // @[NV_NVDLA_CSC_wl.scala 730:86:@17340.4]
  assign _T_1822 = _T_743 | _T_1821; // @[NV_NVDLA_CSC_wl.scala 730:47:@17341.4]
  assign _T_1825 = {_T_1762,3'h0}; // @[Cat.scala 30:58:@17343.4]
  assign _GEN_583 = {{1023'd0}, io_sc2buf_wt_rd_data_bits}; // @[NV_NVDLA_CSC_wl.scala 731:55:@17344.4]
  assign _T_1826 = _GEN_583 << _T_1825; // @[NV_NVDLA_CSC_wl.scala 731:55:@17344.4]
  assign _T_1828 = io_sc2buf_wt_rd_data_valid ? _T_1826 : 1535'h0; // @[NV_NVDLA_CSC_wl.scala 732:32:@17345.4]
  assign _GEN_584 = {{1023'd0}, _T_1801}; // @[NV_NVDLA_CSC_wl.scala 744:42:@17418.4]
  assign _T_2292 = _T_1828 | _GEN_584; // @[NV_NVDLA_CSC_wl.scala 744:42:@17418.4]
  assign _T_2293 = _T_2292[7:0]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17420.6]
  assign _T_2294 = _T_2292[15:8]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17422.6]
  assign _T_2295 = _T_2292[23:16]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17424.6]
  assign _T_2296 = _T_2292[31:24]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17426.6]
  assign _T_2297 = _T_2292[39:32]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17428.6]
  assign _T_2298 = _T_2292[47:40]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17430.6]
  assign _T_2299 = _T_2292[55:48]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17432.6]
  assign _T_2300 = _T_2292[63:56]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17434.6]
  assign _T_2301 = _T_2292[71:64]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17436.6]
  assign _T_2302 = _T_2292[79:72]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17438.6]
  assign _T_2303 = _T_2292[87:80]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17440.6]
  assign _T_2304 = _T_2292[95:88]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17442.6]
  assign _T_2305 = _T_2292[103:96]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17444.6]
  assign _T_2306 = _T_2292[111:104]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17446.6]
  assign _T_2307 = _T_2292[119:112]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17448.6]
  assign _T_2308 = _T_2292[127:120]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17450.6]
  assign _T_2309 = _T_2292[135:128]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17452.6]
  assign _T_2310 = _T_2292[143:136]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17454.6]
  assign _T_2311 = _T_2292[151:144]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17456.6]
  assign _T_2312 = _T_2292[159:152]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17458.6]
  assign _T_2313 = _T_2292[167:160]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17460.6]
  assign _T_2314 = _T_2292[175:168]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17462.6]
  assign _T_2315 = _T_2292[183:176]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17464.6]
  assign _T_2316 = _T_2292[191:184]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17466.6]
  assign _T_2317 = _T_2292[199:192]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17468.6]
  assign _T_2318 = _T_2292[207:200]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17470.6]
  assign _T_2319 = _T_2292[215:208]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17472.6]
  assign _T_2320 = _T_2292[223:216]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17474.6]
  assign _T_2321 = _T_2292[231:224]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17476.6]
  assign _T_2322 = _T_2292[239:232]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17478.6]
  assign _T_2323 = _T_2292[247:240]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17480.6]
  assign _T_2324 = _T_2292[255:248]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17482.6]
  assign _T_2325 = _T_2292[263:256]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17484.6]
  assign _T_2326 = _T_2292[271:264]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17486.6]
  assign _T_2327 = _T_2292[279:272]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17488.6]
  assign _T_2328 = _T_2292[287:280]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17490.6]
  assign _T_2329 = _T_2292[295:288]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17492.6]
  assign _T_2330 = _T_2292[303:296]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17494.6]
  assign _T_2331 = _T_2292[311:304]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17496.6]
  assign _T_2332 = _T_2292[319:312]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17498.6]
  assign _T_2333 = _T_2292[327:320]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17500.6]
  assign _T_2334 = _T_2292[335:328]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17502.6]
  assign _T_2335 = _T_2292[343:336]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17504.6]
  assign _T_2336 = _T_2292[351:344]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17506.6]
  assign _T_2337 = _T_2292[359:352]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17508.6]
  assign _T_2338 = _T_2292[367:360]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17510.6]
  assign _T_2339 = _T_2292[375:368]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17512.6]
  assign _T_2340 = _T_2292[383:376]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17514.6]
  assign _T_2341 = _T_2292[391:384]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17516.6]
  assign _T_2342 = _T_2292[399:392]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17518.6]
  assign _T_2343 = _T_2292[407:400]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17520.6]
  assign _T_2344 = _T_2292[415:408]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17522.6]
  assign _T_2345 = _T_2292[423:416]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17524.6]
  assign _T_2346 = _T_2292[431:424]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17526.6]
  assign _T_2347 = _T_2292[439:432]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17528.6]
  assign _T_2348 = _T_2292[447:440]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17530.6]
  assign _T_2349 = _T_2292[455:448]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17532.6]
  assign _T_2350 = _T_2292[463:456]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17534.6]
  assign _T_2351 = _T_2292[471:464]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17536.6]
  assign _T_2352 = _T_2292[479:472]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17538.6]
  assign _T_2353 = _T_2292[487:480]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17540.6]
  assign _T_2354 = _T_2292[495:488]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17542.6]
  assign _T_2355 = _T_2292[503:496]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17544.6]
  assign _T_2356 = _T_2292[511:504]; // @[NV_NVDLA_CSC_wl.scala 747:45:@17546.6]
  assign _GEN_79 = _T_1692 ? _T_2293 : _T_2095_0; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_80 = _T_1692 ? _T_2294 : _T_2095_1; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_81 = _T_1692 ? _T_2295 : _T_2095_2; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_82 = _T_1692 ? _T_2296 : _T_2095_3; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_83 = _T_1692 ? _T_2297 : _T_2095_4; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_84 = _T_1692 ? _T_2298 : _T_2095_5; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_85 = _T_1692 ? _T_2299 : _T_2095_6; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_86 = _T_1692 ? _T_2300 : _T_2095_7; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_87 = _T_1692 ? _T_2301 : _T_2095_8; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_88 = _T_1692 ? _T_2302 : _T_2095_9; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_89 = _T_1692 ? _T_2303 : _T_2095_10; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_90 = _T_1692 ? _T_2304 : _T_2095_11; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_91 = _T_1692 ? _T_2305 : _T_2095_12; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_92 = _T_1692 ? _T_2306 : _T_2095_13; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_93 = _T_1692 ? _T_2307 : _T_2095_14; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_94 = _T_1692 ? _T_2308 : _T_2095_15; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_95 = _T_1692 ? _T_2309 : _T_2095_16; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_96 = _T_1692 ? _T_2310 : _T_2095_17; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_97 = _T_1692 ? _T_2311 : _T_2095_18; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_98 = _T_1692 ? _T_2312 : _T_2095_19; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_99 = _T_1692 ? _T_2313 : _T_2095_20; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_100 = _T_1692 ? _T_2314 : _T_2095_21; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_101 = _T_1692 ? _T_2315 : _T_2095_22; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_102 = _T_1692 ? _T_2316 : _T_2095_23; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_103 = _T_1692 ? _T_2317 : _T_2095_24; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_104 = _T_1692 ? _T_2318 : _T_2095_25; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_105 = _T_1692 ? _T_2319 : _T_2095_26; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_106 = _T_1692 ? _T_2320 : _T_2095_27; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_107 = _T_1692 ? _T_2321 : _T_2095_28; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_108 = _T_1692 ? _T_2322 : _T_2095_29; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_109 = _T_1692 ? _T_2323 : _T_2095_30; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_110 = _T_1692 ? _T_2324 : _T_2095_31; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_111 = _T_1692 ? _T_2325 : _T_2095_32; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_112 = _T_1692 ? _T_2326 : _T_2095_33; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_113 = _T_1692 ? _T_2327 : _T_2095_34; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_114 = _T_1692 ? _T_2328 : _T_2095_35; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_115 = _T_1692 ? _T_2329 : _T_2095_36; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_116 = _T_1692 ? _T_2330 : _T_2095_37; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_117 = _T_1692 ? _T_2331 : _T_2095_38; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_118 = _T_1692 ? _T_2332 : _T_2095_39; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_119 = _T_1692 ? _T_2333 : _T_2095_40; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_120 = _T_1692 ? _T_2334 : _T_2095_41; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_121 = _T_1692 ? _T_2335 : _T_2095_42; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_122 = _T_1692 ? _T_2336 : _T_2095_43; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_123 = _T_1692 ? _T_2337 : _T_2095_44; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_124 = _T_1692 ? _T_2338 : _T_2095_45; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_125 = _T_1692 ? _T_2339 : _T_2095_46; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_126 = _T_1692 ? _T_2340 : _T_2095_47; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_127 = _T_1692 ? _T_2341 : _T_2095_48; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_128 = _T_1692 ? _T_2342 : _T_2095_49; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_129 = _T_1692 ? _T_2343 : _T_2095_50; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_130 = _T_1692 ? _T_2344 : _T_2095_51; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_131 = _T_1692 ? _T_2345 : _T_2095_52; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_132 = _T_1692 ? _T_2346 : _T_2095_53; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_133 = _T_1692 ? _T_2347 : _T_2095_54; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_134 = _T_1692 ? _T_2348 : _T_2095_55; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_135 = _T_1692 ? _T_2349 : _T_2095_56; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_136 = _T_1692 ? _T_2350 : _T_2095_57; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_137 = _T_1692 ? _T_2351 : _T_2095_58; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_138 = _T_1692 ? _T_2352 : _T_2095_59; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_139 = _T_1692 ? _T_2353 : _T_2095_60; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_140 = _T_1692 ? _T_2354 : _T_2095_61; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_141 = _T_1692 ? _T_2355 : _T_2095_62; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _GEN_142 = _T_1692 ? _T_2356 : _T_2095_63; // @[NV_NVDLA_CSC_wl.scala 745:27:@17419.4]
  assign _T_2364 = _T_2362[30:0]; // @[NV_NVDLA_CSC_wl.scala 757:41:@17551.4]
  assign _T_2365 = _T_2362[31]; // @[NV_NVDLA_CSC_wl.scala 757:77:@17552.4]
  assign _T_2366 = {_T_2364,_T_2365}; // @[Cat.scala 30:58:@17553.4]
  assign _T_2367 = _T_2359 ? 32'h1 : _T_2366; // @[NV_NVDLA_CSC_wl.scala 756:27:@17554.4]
  assign _GEN_143 = _T_1692 ? _T_1756 : _T_2359; // @[NV_NVDLA_CSC_wl.scala 759:27:@17555.4]
  assign _GEN_144 = _T_1692 ? _T_2367 : _T_2362; // @[NV_NVDLA_CSC_wl.scala 759:27:@17555.4]
  assign _T_2939 = _T_1752[0]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17726.6]
  assign _T_2940 = _T_1752[1]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17727.6]
  assign _T_2941 = _T_1752[2]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17728.6]
  assign _T_2942 = _T_1752[3]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17729.6]
  assign _T_2943 = _T_1752[4]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17730.6]
  assign _T_2944 = _T_1752[5]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17731.6]
  assign _T_2945 = _T_1752[6]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17732.6]
  assign _T_2946 = _T_1752[7]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17733.6]
  assign _T_2947 = _T_1752[8]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17734.6]
  assign _T_2948 = _T_1752[9]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17735.6]
  assign _T_2949 = _T_1752[10]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17736.6]
  assign _T_2950 = _T_1752[11]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17737.6]
  assign _T_2951 = _T_1752[12]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17738.6]
  assign _T_2952 = _T_1752[13]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17739.6]
  assign _T_2953 = _T_1752[14]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17740.6]
  assign _T_2954 = _T_1752[15]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17741.6]
  assign _T_2955 = _T_1752[16]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17742.6]
  assign _T_2956 = _T_1752[17]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17743.6]
  assign _T_2957 = _T_1752[18]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17744.6]
  assign _T_2958 = _T_1752[19]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17745.6]
  assign _T_2959 = _T_1752[20]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17746.6]
  assign _T_2960 = _T_1752[21]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17747.6]
  assign _T_2961 = _T_1752[22]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17748.6]
  assign _T_2962 = _T_1752[23]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17749.6]
  assign _T_2963 = _T_1752[24]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17750.6]
  assign _T_2964 = _T_1752[25]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17751.6]
  assign _T_2965 = _T_1752[26]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17752.6]
  assign _T_2966 = _T_1752[27]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17753.6]
  assign _T_2967 = _T_1752[28]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17754.6]
  assign _T_2968 = _T_1752[29]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17755.6]
  assign _T_2969 = _T_1752[30]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17756.6]
  assign _T_2970 = _T_1752[31]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17757.6]
  assign _T_2971 = _T_1752[32]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17758.6]
  assign _T_2972 = _T_1752[33]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17759.6]
  assign _T_2973 = _T_1752[34]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17760.6]
  assign _T_2974 = _T_1752[35]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17761.6]
  assign _T_2975 = _T_1752[36]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17762.6]
  assign _T_2976 = _T_1752[37]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17763.6]
  assign _T_2977 = _T_1752[38]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17764.6]
  assign _T_2978 = _T_1752[39]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17765.6]
  assign _T_2979 = _T_1752[40]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17766.6]
  assign _T_2980 = _T_1752[41]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17767.6]
  assign _T_2981 = _T_1752[42]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17768.6]
  assign _T_2982 = _T_1752[43]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17769.6]
  assign _T_2983 = _T_1752[44]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17770.6]
  assign _T_2984 = _T_1752[45]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17771.6]
  assign _T_2985 = _T_1752[46]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17772.6]
  assign _T_2986 = _T_1752[47]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17773.6]
  assign _T_2987 = _T_1752[48]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17774.6]
  assign _T_2988 = _T_1752[49]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17775.6]
  assign _T_2989 = _T_1752[50]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17776.6]
  assign _T_2990 = _T_1752[51]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17777.6]
  assign _T_2991 = _T_1752[52]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17778.6]
  assign _T_2992 = _T_1752[53]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17779.6]
  assign _T_2993 = _T_1752[54]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17780.6]
  assign _T_2994 = _T_1752[55]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17781.6]
  assign _T_2995 = _T_1752[56]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17782.6]
  assign _T_2996 = _T_1752[57]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17783.6]
  assign _T_2997 = _T_1752[58]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17784.6]
  assign _T_2998 = _T_1752[59]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17785.6]
  assign _T_2999 = _T_1752[60]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17786.6]
  assign _T_3000 = _T_1752[61]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17787.6]
  assign _T_3001 = _T_1752[62]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17788.6]
  assign _T_3002 = _T_1752[63]; // @[NV_NVDLA_CSC_wl.scala 773:86:@17789.6]
  assign _GEN_145 = _T_1732 ? _T_2939 : _T_2739_0; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_146 = _T_1732 ? _T_2940 : _T_2739_1; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_147 = _T_1732 ? _T_2941 : _T_2739_2; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_148 = _T_1732 ? _T_2942 : _T_2739_3; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_149 = _T_1732 ? _T_2943 : _T_2739_4; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_150 = _T_1732 ? _T_2944 : _T_2739_5; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_151 = _T_1732 ? _T_2945 : _T_2739_6; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_152 = _T_1732 ? _T_2946 : _T_2739_7; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_153 = _T_1732 ? _T_2947 : _T_2739_8; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_154 = _T_1732 ? _T_2948 : _T_2739_9; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_155 = _T_1732 ? _T_2949 : _T_2739_10; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_156 = _T_1732 ? _T_2950 : _T_2739_11; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_157 = _T_1732 ? _T_2951 : _T_2739_12; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_158 = _T_1732 ? _T_2952 : _T_2739_13; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_159 = _T_1732 ? _T_2953 : _T_2739_14; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_160 = _T_1732 ? _T_2954 : _T_2739_15; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_161 = _T_1732 ? _T_2955 : _T_2739_16; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_162 = _T_1732 ? _T_2956 : _T_2739_17; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_163 = _T_1732 ? _T_2957 : _T_2739_18; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_164 = _T_1732 ? _T_2958 : _T_2739_19; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_165 = _T_1732 ? _T_2959 : _T_2739_20; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_166 = _T_1732 ? _T_2960 : _T_2739_21; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_167 = _T_1732 ? _T_2961 : _T_2739_22; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_168 = _T_1732 ? _T_2962 : _T_2739_23; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_169 = _T_1732 ? _T_2963 : _T_2739_24; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_170 = _T_1732 ? _T_2964 : _T_2739_25; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_171 = _T_1732 ? _T_2965 : _T_2739_26; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_172 = _T_1732 ? _T_2966 : _T_2739_27; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_173 = _T_1732 ? _T_2967 : _T_2739_28; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_174 = _T_1732 ? _T_2968 : _T_2739_29; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_175 = _T_1732 ? _T_2969 : _T_2739_30; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_176 = _T_1732 ? _T_2970 : _T_2739_31; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_177 = _T_1732 ? _T_2971 : _T_2739_32; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_178 = _T_1732 ? _T_2972 : _T_2739_33; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_179 = _T_1732 ? _T_2973 : _T_2739_34; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_180 = _T_1732 ? _T_2974 : _T_2739_35; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_181 = _T_1732 ? _T_2975 : _T_2739_36; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_182 = _T_1732 ? _T_2976 : _T_2739_37; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_183 = _T_1732 ? _T_2977 : _T_2739_38; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_184 = _T_1732 ? _T_2978 : _T_2739_39; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_185 = _T_1732 ? _T_2979 : _T_2739_40; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_186 = _T_1732 ? _T_2980 : _T_2739_41; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_187 = _T_1732 ? _T_2981 : _T_2739_42; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_188 = _T_1732 ? _T_2982 : _T_2739_43; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_189 = _T_1732 ? _T_2983 : _T_2739_44; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_190 = _T_1732 ? _T_2984 : _T_2739_45; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_191 = _T_1732 ? _T_2985 : _T_2739_46; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_192 = _T_1732 ? _T_2986 : _T_2739_47; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_193 = _T_1732 ? _T_2987 : _T_2739_48; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_194 = _T_1732 ? _T_2988 : _T_2739_49; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_195 = _T_1732 ? _T_2989 : _T_2739_50; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_196 = _T_1732 ? _T_2990 : _T_2739_51; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_197 = _T_1732 ? _T_2991 : _T_2739_52; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_198 = _T_1732 ? _T_2992 : _T_2739_53; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_199 = _T_1732 ? _T_2993 : _T_2739_54; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_200 = _T_1732 ? _T_2994 : _T_2739_55; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_201 = _T_1732 ? _T_2995 : _T_2739_56; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_202 = _T_1732 ? _T_2996 : _T_2739_57; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_203 = _T_1732 ? _T_2997 : _T_2739_58; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_204 = _T_1732 ? _T_2998 : _T_2739_59; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_205 = _T_1732 ? _T_2999 : _T_2739_60; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_206 = _T_1732 ? _T_3000 : _T_2739_61; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_207 = _T_1732 ? _T_3001 : _T_2739_62; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _GEN_208 = _T_1732 ? _T_3002 : _T_2739_63; // @[NV_NVDLA_CSC_wl.scala 772:25:@17725.4]
  assign _T_3076 = _T_1732 ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12:@17921.4]
  assign _T_3077 = NV_NVDLA_CSC_WL_dec_io_output_valid; // @[Bitwise.scala 72:15:@18089.4]
  assign _T_3080 = _T_3077 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@18090.4]
  assign _T_3087 = {NV_NVDLA_CSC_WL_dec_io_output_bits_sel_7,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_6,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_5,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_4,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_3,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_2,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_1,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_0}; // @[NV_NVDLA_CSC_wl.scala 794:92:@18097.4]
  assign _T_3095 = {NV_NVDLA_CSC_WL_dec_io_output_bits_sel_15,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_14,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_13,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_12,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_11,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_10,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_9,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_8,_T_3087}; // @[NV_NVDLA_CSC_wl.scala 794:92:@18105.4]
  assign _T_3102 = {NV_NVDLA_CSC_WL_dec_io_output_bits_sel_23,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_22,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_21,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_20,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_19,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_18,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_17,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_16}; // @[NV_NVDLA_CSC_wl.scala 794:92:@18112.4]
  assign _T_3111 = {NV_NVDLA_CSC_WL_dec_io_output_bits_sel_31,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_30,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_29,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_28,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_27,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_26,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_25,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_24,_T_3102,_T_3095}; // @[NV_NVDLA_CSC_wl.scala 794:92:@18121.4]
  assign _T_3112 = _T_3111[15:0]; // @[NV_NVDLA_CSC_wl.scala 794:99:@18122.4]
  assign _T_3113 = _T_3080 & _T_3112; // @[NV_NVDLA_CSC_wl.scala 794:71:@18123.4]
  assign _T_3149 = _T_3111[31:16]; // @[NV_NVDLA_CSC_wl.scala 795:99:@18157.4]
  assign _T_3150 = _T_3080 & _T_3149; // @[NV_NVDLA_CSC_wl.scala 795:71:@18158.4]
  assign _T_3152 = _T_3113 != 16'h0; // @[NV_NVDLA_CSC_wl.scala 796:49:@18159.4]
  assign _T_3154 = _T_3150 != 16'h0; // @[NV_NVDLA_CSC_wl.scala 797:49:@18160.4]
  assign _T_4481 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_0; // @[NV_NVDLA_CSC_wl.scala 807:91:@18333.4]
  assign _T_4482 = _T_4481 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18334.4]
  assign _T_4483 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_1; // @[NV_NVDLA_CSC_wl.scala 807:91:@18335.4]
  assign _T_4484 = _T_4483 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18336.4]
  assign _T_4485 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_2; // @[NV_NVDLA_CSC_wl.scala 807:91:@18337.4]
  assign _T_4486 = _T_4485 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18338.4]
  assign _T_4487 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_3; // @[NV_NVDLA_CSC_wl.scala 807:91:@18339.4]
  assign _T_4488 = _T_4487 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18340.4]
  assign _T_4489 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_4; // @[NV_NVDLA_CSC_wl.scala 807:91:@18341.4]
  assign _T_4490 = _T_4489 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18342.4]
  assign _T_4491 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_5; // @[NV_NVDLA_CSC_wl.scala 807:91:@18343.4]
  assign _T_4492 = _T_4491 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18344.4]
  assign _T_4493 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_6; // @[NV_NVDLA_CSC_wl.scala 807:91:@18345.4]
  assign _T_4494 = _T_4493 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18346.4]
  assign _T_4495 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_7; // @[NV_NVDLA_CSC_wl.scala 807:91:@18347.4]
  assign _T_4496 = _T_4495 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18348.4]
  assign _T_4497 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_8; // @[NV_NVDLA_CSC_wl.scala 807:91:@18349.4]
  assign _T_4498 = _T_4497 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18350.4]
  assign _T_4499 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_9; // @[NV_NVDLA_CSC_wl.scala 807:91:@18351.4]
  assign _T_4500 = _T_4499 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18352.4]
  assign _T_4501 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_10; // @[NV_NVDLA_CSC_wl.scala 807:91:@18353.4]
  assign _T_4502 = _T_4501 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18354.4]
  assign _T_4503 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_11; // @[NV_NVDLA_CSC_wl.scala 807:91:@18355.4]
  assign _T_4504 = _T_4503 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18356.4]
  assign _T_4505 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_12; // @[NV_NVDLA_CSC_wl.scala 807:91:@18357.4]
  assign _T_4506 = _T_4505 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18358.4]
  assign _T_4507 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_13; // @[NV_NVDLA_CSC_wl.scala 807:91:@18359.4]
  assign _T_4508 = _T_4507 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18360.4]
  assign _T_4509 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_14; // @[NV_NVDLA_CSC_wl.scala 807:91:@18361.4]
  assign _T_4510 = _T_4509 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18362.4]
  assign _T_4511 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_15; // @[NV_NVDLA_CSC_wl.scala 807:91:@18363.4]
  assign _T_4512 = _T_4511 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18364.4]
  assign _T_4513 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_16; // @[NV_NVDLA_CSC_wl.scala 807:91:@18365.4]
  assign _T_4514 = _T_4513 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18366.4]
  assign _T_4515 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_17; // @[NV_NVDLA_CSC_wl.scala 807:91:@18367.4]
  assign _T_4516 = _T_4515 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18368.4]
  assign _T_4517 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_18; // @[NV_NVDLA_CSC_wl.scala 807:91:@18369.4]
  assign _T_4518 = _T_4517 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18370.4]
  assign _T_4519 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_19; // @[NV_NVDLA_CSC_wl.scala 807:91:@18371.4]
  assign _T_4520 = _T_4519 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18372.4]
  assign _T_4521 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_20; // @[NV_NVDLA_CSC_wl.scala 807:91:@18373.4]
  assign _T_4522 = _T_4521 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18374.4]
  assign _T_4523 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_21; // @[NV_NVDLA_CSC_wl.scala 807:91:@18375.4]
  assign _T_4524 = _T_4523 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18376.4]
  assign _T_4525 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_22; // @[NV_NVDLA_CSC_wl.scala 807:91:@18377.4]
  assign _T_4526 = _T_4525 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18378.4]
  assign _T_4527 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_23; // @[NV_NVDLA_CSC_wl.scala 807:91:@18379.4]
  assign _T_4528 = _T_4527 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18380.4]
  assign _T_4529 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_24; // @[NV_NVDLA_CSC_wl.scala 807:91:@18381.4]
  assign _T_4530 = _T_4529 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18382.4]
  assign _T_4531 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_25; // @[NV_NVDLA_CSC_wl.scala 807:91:@18383.4]
  assign _T_4532 = _T_4531 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18384.4]
  assign _T_4533 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_26; // @[NV_NVDLA_CSC_wl.scala 807:91:@18385.4]
  assign _T_4534 = _T_4533 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18386.4]
  assign _T_4535 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_27; // @[NV_NVDLA_CSC_wl.scala 807:91:@18387.4]
  assign _T_4536 = _T_4535 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18388.4]
  assign _T_4537 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_28; // @[NV_NVDLA_CSC_wl.scala 807:91:@18389.4]
  assign _T_4538 = _T_4537 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18390.4]
  assign _T_4539 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_29; // @[NV_NVDLA_CSC_wl.scala 807:91:@18391.4]
  assign _T_4540 = _T_4539 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18392.4]
  assign _T_4541 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_30; // @[NV_NVDLA_CSC_wl.scala 807:91:@18393.4]
  assign _T_4542 = _T_4541 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18394.4]
  assign _T_4543 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_31; // @[NV_NVDLA_CSC_wl.scala 807:91:@18395.4]
  assign _T_4544 = _T_4543 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18396.4]
  assign _T_4545 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_32; // @[NV_NVDLA_CSC_wl.scala 807:91:@18397.4]
  assign _T_4546 = _T_4545 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18398.4]
  assign _T_4547 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_33; // @[NV_NVDLA_CSC_wl.scala 807:91:@18399.4]
  assign _T_4548 = _T_4547 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18400.4]
  assign _T_4549 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_34; // @[NV_NVDLA_CSC_wl.scala 807:91:@18401.4]
  assign _T_4550 = _T_4549 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18402.4]
  assign _T_4551 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_35; // @[NV_NVDLA_CSC_wl.scala 807:91:@18403.4]
  assign _T_4552 = _T_4551 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18404.4]
  assign _T_4553 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_36; // @[NV_NVDLA_CSC_wl.scala 807:91:@18405.4]
  assign _T_4554 = _T_4553 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18406.4]
  assign _T_4555 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_37; // @[NV_NVDLA_CSC_wl.scala 807:91:@18407.4]
  assign _T_4556 = _T_4555 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18408.4]
  assign _T_4557 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_38; // @[NV_NVDLA_CSC_wl.scala 807:91:@18409.4]
  assign _T_4558 = _T_4557 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18410.4]
  assign _T_4559 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_39; // @[NV_NVDLA_CSC_wl.scala 807:91:@18411.4]
  assign _T_4560 = _T_4559 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18412.4]
  assign _T_4561 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_40; // @[NV_NVDLA_CSC_wl.scala 807:91:@18413.4]
  assign _T_4562 = _T_4561 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18414.4]
  assign _T_4563 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_41; // @[NV_NVDLA_CSC_wl.scala 807:91:@18415.4]
  assign _T_4564 = _T_4563 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18416.4]
  assign _T_4565 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_42; // @[NV_NVDLA_CSC_wl.scala 807:91:@18417.4]
  assign _T_4566 = _T_4565 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18418.4]
  assign _T_4567 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_43; // @[NV_NVDLA_CSC_wl.scala 807:91:@18419.4]
  assign _T_4568 = _T_4567 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18420.4]
  assign _T_4569 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_44; // @[NV_NVDLA_CSC_wl.scala 807:91:@18421.4]
  assign _T_4570 = _T_4569 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18422.4]
  assign _T_4571 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_45; // @[NV_NVDLA_CSC_wl.scala 807:91:@18423.4]
  assign _T_4572 = _T_4571 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18424.4]
  assign _T_4573 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_46; // @[NV_NVDLA_CSC_wl.scala 807:91:@18425.4]
  assign _T_4574 = _T_4573 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18426.4]
  assign _T_4575 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_47; // @[NV_NVDLA_CSC_wl.scala 807:91:@18427.4]
  assign _T_4576 = _T_4575 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18428.4]
  assign _T_4577 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_48; // @[NV_NVDLA_CSC_wl.scala 807:91:@18429.4]
  assign _T_4578 = _T_4577 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18430.4]
  assign _T_4579 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_49; // @[NV_NVDLA_CSC_wl.scala 807:91:@18431.4]
  assign _T_4580 = _T_4579 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18432.4]
  assign _T_4581 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_50; // @[NV_NVDLA_CSC_wl.scala 807:91:@18433.4]
  assign _T_4582 = _T_4581 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18434.4]
  assign _T_4583 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_51; // @[NV_NVDLA_CSC_wl.scala 807:91:@18435.4]
  assign _T_4584 = _T_4583 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18436.4]
  assign _T_4585 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_52; // @[NV_NVDLA_CSC_wl.scala 807:91:@18437.4]
  assign _T_4586 = _T_4585 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18438.4]
  assign _T_4587 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_53; // @[NV_NVDLA_CSC_wl.scala 807:91:@18439.4]
  assign _T_4588 = _T_4587 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18440.4]
  assign _T_4589 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_54; // @[NV_NVDLA_CSC_wl.scala 807:91:@18441.4]
  assign _T_4590 = _T_4589 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18442.4]
  assign _T_4591 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_55; // @[NV_NVDLA_CSC_wl.scala 807:91:@18443.4]
  assign _T_4592 = _T_4591 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18444.4]
  assign _T_4593 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_56; // @[NV_NVDLA_CSC_wl.scala 807:91:@18445.4]
  assign _T_4594 = _T_4593 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18446.4]
  assign _T_4595 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_57; // @[NV_NVDLA_CSC_wl.scala 807:91:@18447.4]
  assign _T_4596 = _T_4595 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18448.4]
  assign _T_4597 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_58; // @[NV_NVDLA_CSC_wl.scala 807:91:@18449.4]
  assign _T_4598 = _T_4597 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18450.4]
  assign _T_4599 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_59; // @[NV_NVDLA_CSC_wl.scala 807:91:@18451.4]
  assign _T_4600 = _T_4599 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18452.4]
  assign _T_4601 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_60; // @[NV_NVDLA_CSC_wl.scala 807:91:@18453.4]
  assign _T_4602 = _T_4601 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18454.4]
  assign _T_4603 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_61; // @[NV_NVDLA_CSC_wl.scala 807:91:@18455.4]
  assign _T_4604 = _T_4603 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18456.4]
  assign _T_4605 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_62; // @[NV_NVDLA_CSC_wl.scala 807:91:@18457.4]
  assign _T_4606 = _T_4605 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18458.4]
  assign _T_4607 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_63; // @[NV_NVDLA_CSC_wl.scala 807:91:@18459.4]
  assign _T_4608 = _T_4607 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@18460.4]
  assign _T_4680 = _T_4481 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18527.4]
  assign _T_4682 = _T_4483 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18529.4]
  assign _T_4684 = _T_4485 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18531.4]
  assign _T_4686 = _T_4487 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18533.4]
  assign _T_4688 = _T_4489 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18535.4]
  assign _T_4690 = _T_4491 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18537.4]
  assign _T_4692 = _T_4493 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18539.4]
  assign _T_4694 = _T_4495 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18541.4]
  assign _T_4696 = _T_4497 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18543.4]
  assign _T_4698 = _T_4499 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18545.4]
  assign _T_4700 = _T_4501 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18547.4]
  assign _T_4702 = _T_4503 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18549.4]
  assign _T_4704 = _T_4505 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18551.4]
  assign _T_4706 = _T_4507 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18553.4]
  assign _T_4708 = _T_4509 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18555.4]
  assign _T_4710 = _T_4511 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18557.4]
  assign _T_4712 = _T_4513 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18559.4]
  assign _T_4714 = _T_4515 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18561.4]
  assign _T_4716 = _T_4517 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18563.4]
  assign _T_4718 = _T_4519 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18565.4]
  assign _T_4720 = _T_4521 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18567.4]
  assign _T_4722 = _T_4523 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18569.4]
  assign _T_4724 = _T_4525 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18571.4]
  assign _T_4726 = _T_4527 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18573.4]
  assign _T_4728 = _T_4529 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18575.4]
  assign _T_4730 = _T_4531 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18577.4]
  assign _T_4732 = _T_4533 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18579.4]
  assign _T_4734 = _T_4535 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18581.4]
  assign _T_4736 = _T_4537 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18583.4]
  assign _T_4738 = _T_4539 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18585.4]
  assign _T_4740 = _T_4541 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18587.4]
  assign _T_4742 = _T_4543 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18589.4]
  assign _T_4744 = _T_4545 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18591.4]
  assign _T_4746 = _T_4547 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18593.4]
  assign _T_4748 = _T_4549 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18595.4]
  assign _T_4750 = _T_4551 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18597.4]
  assign _T_4752 = _T_4553 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18599.4]
  assign _T_4754 = _T_4555 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18601.4]
  assign _T_4756 = _T_4557 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18603.4]
  assign _T_4758 = _T_4559 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18605.4]
  assign _T_4760 = _T_4561 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18607.4]
  assign _T_4762 = _T_4563 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18609.4]
  assign _T_4764 = _T_4565 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18611.4]
  assign _T_4766 = _T_4567 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18613.4]
  assign _T_4768 = _T_4569 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18615.4]
  assign _T_4770 = _T_4571 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18617.4]
  assign _T_4772 = _T_4573 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18619.4]
  assign _T_4774 = _T_4575 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18621.4]
  assign _T_4776 = _T_4577 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18623.4]
  assign _T_4778 = _T_4579 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18625.4]
  assign _T_4780 = _T_4581 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18627.4]
  assign _T_4782 = _T_4583 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18629.4]
  assign _T_4784 = _T_4585 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18631.4]
  assign _T_4786 = _T_4587 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18633.4]
  assign _T_4788 = _T_4589 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18635.4]
  assign _T_4790 = _T_4591 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18637.4]
  assign _T_4792 = _T_4593 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18639.4]
  assign _T_4794 = _T_4595 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18641.4]
  assign _T_4796 = _T_4597 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18643.4]
  assign _T_4798 = _T_4599 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18645.4]
  assign _T_4800 = _T_4601 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18647.4]
  assign _T_4802 = _T_4603 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18649.4]
  assign _T_4804 = _T_4605 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18651.4]
  assign _T_4806 = _T_4607 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@18653.4]
  assign _T_4877 = _T_3152 | _T_3157; // @[NV_NVDLA_CSC_wl.scala 812:29:@18721.4]
  assign _T_4878 = _T_3113[0]; // @[NV_NVDLA_CSC_wl.scala 814:96:@18787.6]
  assign _T_4879 = _T_3113[1]; // @[NV_NVDLA_CSC_wl.scala 814:96:@18788.6]
  assign _T_4880 = _T_3113[2]; // @[NV_NVDLA_CSC_wl.scala 814:96:@18789.6]
  assign _T_4881 = _T_3113[3]; // @[NV_NVDLA_CSC_wl.scala 814:96:@18790.6]
  assign _T_4882 = _T_3113[4]; // @[NV_NVDLA_CSC_wl.scala 814:96:@18791.6]
  assign _T_4883 = _T_3113[5]; // @[NV_NVDLA_CSC_wl.scala 814:96:@18792.6]
  assign _T_4884 = _T_3113[6]; // @[NV_NVDLA_CSC_wl.scala 814:96:@18793.6]
  assign _T_4885 = _T_3113[7]; // @[NV_NVDLA_CSC_wl.scala 814:96:@18794.6]
  assign _T_4886 = _T_3113[8]; // @[NV_NVDLA_CSC_wl.scala 814:96:@18795.6]
  assign _T_4887 = _T_3113[9]; // @[NV_NVDLA_CSC_wl.scala 814:96:@18796.6]
  assign _T_4888 = _T_3113[10]; // @[NV_NVDLA_CSC_wl.scala 814:96:@18797.6]
  assign _T_4889 = _T_3113[11]; // @[NV_NVDLA_CSC_wl.scala 814:96:@18798.6]
  assign _T_4890 = _T_3113[12]; // @[NV_NVDLA_CSC_wl.scala 814:96:@18799.6]
  assign _T_4891 = _T_3113[13]; // @[NV_NVDLA_CSC_wl.scala 814:96:@18800.6]
  assign _T_4892 = _T_3113[14]; // @[NV_NVDLA_CSC_wl.scala 814:96:@18801.6]
  assign _T_4893 = _T_3113[15]; // @[NV_NVDLA_CSC_wl.scala 814:96:@18802.6]
  assign _GEN_209 = _T_4877 ? _T_4482 : _T_3427_0; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_210 = _T_4877 ? _T_4484 : _T_3427_1; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_211 = _T_4877 ? _T_4486 : _T_3427_2; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_212 = _T_4877 ? _T_4488 : _T_3427_3; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_213 = _T_4877 ? _T_4490 : _T_3427_4; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_214 = _T_4877 ? _T_4492 : _T_3427_5; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_215 = _T_4877 ? _T_4494 : _T_3427_6; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_216 = _T_4877 ? _T_4496 : _T_3427_7; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_217 = _T_4877 ? _T_4498 : _T_3427_8; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_218 = _T_4877 ? _T_4500 : _T_3427_9; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_219 = _T_4877 ? _T_4502 : _T_3427_10; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_220 = _T_4877 ? _T_4504 : _T_3427_11; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_221 = _T_4877 ? _T_4506 : _T_3427_12; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_222 = _T_4877 ? _T_4508 : _T_3427_13; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_223 = _T_4877 ? _T_4510 : _T_3427_14; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_224 = _T_4877 ? _T_4512 : _T_3427_15; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_225 = _T_4877 ? _T_4514 : _T_3427_16; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_226 = _T_4877 ? _T_4516 : _T_3427_17; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_227 = _T_4877 ? _T_4518 : _T_3427_18; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_228 = _T_4877 ? _T_4520 : _T_3427_19; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_229 = _T_4877 ? _T_4522 : _T_3427_20; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_230 = _T_4877 ? _T_4524 : _T_3427_21; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_231 = _T_4877 ? _T_4526 : _T_3427_22; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_232 = _T_4877 ? _T_4528 : _T_3427_23; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_233 = _T_4877 ? _T_4530 : _T_3427_24; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_234 = _T_4877 ? _T_4532 : _T_3427_25; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_235 = _T_4877 ? _T_4534 : _T_3427_26; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_236 = _T_4877 ? _T_4536 : _T_3427_27; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_237 = _T_4877 ? _T_4538 : _T_3427_28; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_238 = _T_4877 ? _T_4540 : _T_3427_29; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_239 = _T_4877 ? _T_4542 : _T_3427_30; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_240 = _T_4877 ? _T_4544 : _T_3427_31; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_241 = _T_4877 ? _T_4546 : _T_3427_32; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_242 = _T_4877 ? _T_4548 : _T_3427_33; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_243 = _T_4877 ? _T_4550 : _T_3427_34; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_244 = _T_4877 ? _T_4552 : _T_3427_35; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_245 = _T_4877 ? _T_4554 : _T_3427_36; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_246 = _T_4877 ? _T_4556 : _T_3427_37; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_247 = _T_4877 ? _T_4558 : _T_3427_38; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_248 = _T_4877 ? _T_4560 : _T_3427_39; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_249 = _T_4877 ? _T_4562 : _T_3427_40; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_250 = _T_4877 ? _T_4564 : _T_3427_41; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_251 = _T_4877 ? _T_4566 : _T_3427_42; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_252 = _T_4877 ? _T_4568 : _T_3427_43; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_253 = _T_4877 ? _T_4570 : _T_3427_44; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_254 = _T_4877 ? _T_4572 : _T_3427_45; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_255 = _T_4877 ? _T_4574 : _T_3427_46; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_256 = _T_4877 ? _T_4576 : _T_3427_47; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_257 = _T_4877 ? _T_4578 : _T_3427_48; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_258 = _T_4877 ? _T_4580 : _T_3427_49; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_259 = _T_4877 ? _T_4582 : _T_3427_50; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_260 = _T_4877 ? _T_4584 : _T_3427_51; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_261 = _T_4877 ? _T_4586 : _T_3427_52; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_262 = _T_4877 ? _T_4588 : _T_3427_53; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_263 = _T_4877 ? _T_4590 : _T_3427_54; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_264 = _T_4877 ? _T_4592 : _T_3427_55; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_265 = _T_4877 ? _T_4594 : _T_3427_56; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_266 = _T_4877 ? _T_4596 : _T_3427_57; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_267 = _T_4877 ? _T_4598 : _T_3427_58; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_268 = _T_4877 ? _T_4600 : _T_3427_59; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_269 = _T_4877 ? _T_4602 : _T_3427_60; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_270 = _T_4877 ? _T_4604 : _T_3427_61; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_271 = _T_4877 ? _T_4606 : _T_3427_62; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_272 = _T_4877 ? _T_4608 : _T_3427_63; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_273 = _T_4877 ? _T_4878 : _T_4161_0; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_274 = _T_4877 ? _T_4879 : _T_4161_1; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_275 = _T_4877 ? _T_4880 : _T_4161_2; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_276 = _T_4877 ? _T_4881 : _T_4161_3; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_277 = _T_4877 ? _T_4882 : _T_4161_4; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_278 = _T_4877 ? _T_4883 : _T_4161_5; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_279 = _T_4877 ? _T_4884 : _T_4161_6; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_280 = _T_4877 ? _T_4885 : _T_4161_7; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_281 = _T_4877 ? _T_4886 : _T_4161_8; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_282 = _T_4877 ? _T_4887 : _T_4161_9; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_283 = _T_4877 ? _T_4888 : _T_4161_10; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_284 = _T_4877 ? _T_4889 : _T_4161_11; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_285 = _T_4877 ? _T_4890 : _T_4161_12; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_286 = _T_4877 ? _T_4891 : _T_4161_13; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_287 = _T_4877 ? _T_4892 : _T_4161_14; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _GEN_288 = _T_4877 ? _T_4893 : _T_4161_15; // @[NV_NVDLA_CSC_wl.scala 812:52:@18722.4]
  assign _T_4916 = _T_3154 | _T_3160; // @[NV_NVDLA_CSC_wl.scala 816:29:@18837.4]
  assign _T_4917 = _T_3150[0]; // @[NV_NVDLA_CSC_wl.scala 818:96:@18903.6]
  assign _T_4918 = _T_3150[1]; // @[NV_NVDLA_CSC_wl.scala 818:96:@18904.6]
  assign _T_4919 = _T_3150[2]; // @[NV_NVDLA_CSC_wl.scala 818:96:@18905.6]
  assign _T_4920 = _T_3150[3]; // @[NV_NVDLA_CSC_wl.scala 818:96:@18906.6]
  assign _T_4921 = _T_3150[4]; // @[NV_NVDLA_CSC_wl.scala 818:96:@18907.6]
  assign _T_4922 = _T_3150[5]; // @[NV_NVDLA_CSC_wl.scala 818:96:@18908.6]
  assign _T_4923 = _T_3150[6]; // @[NV_NVDLA_CSC_wl.scala 818:96:@18909.6]
  assign _T_4924 = _T_3150[7]; // @[NV_NVDLA_CSC_wl.scala 818:96:@18910.6]
  assign _T_4925 = _T_3150[8]; // @[NV_NVDLA_CSC_wl.scala 818:96:@18911.6]
  assign _T_4926 = _T_3150[9]; // @[NV_NVDLA_CSC_wl.scala 818:96:@18912.6]
  assign _T_4927 = _T_3150[10]; // @[NV_NVDLA_CSC_wl.scala 818:96:@18913.6]
  assign _T_4928 = _T_3150[11]; // @[NV_NVDLA_CSC_wl.scala 818:96:@18914.6]
  assign _T_4929 = _T_3150[12]; // @[NV_NVDLA_CSC_wl.scala 818:96:@18915.6]
  assign _T_4930 = _T_3150[13]; // @[NV_NVDLA_CSC_wl.scala 818:96:@18916.6]
  assign _T_4931 = _T_3150[14]; // @[NV_NVDLA_CSC_wl.scala 818:96:@18917.6]
  assign _T_4932 = _T_3150[15]; // @[NV_NVDLA_CSC_wl.scala 818:96:@18918.6]
  assign _GEN_289 = _T_4916 ? _T_4680 : _T_3890_0; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_290 = _T_4916 ? _T_4682 : _T_3890_1; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_291 = _T_4916 ? _T_4684 : _T_3890_2; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_292 = _T_4916 ? _T_4686 : _T_3890_3; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_293 = _T_4916 ? _T_4688 : _T_3890_4; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_294 = _T_4916 ? _T_4690 : _T_3890_5; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_295 = _T_4916 ? _T_4692 : _T_3890_6; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_296 = _T_4916 ? _T_4694 : _T_3890_7; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_297 = _T_4916 ? _T_4696 : _T_3890_8; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_298 = _T_4916 ? _T_4698 : _T_3890_9; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_299 = _T_4916 ? _T_4700 : _T_3890_10; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_300 = _T_4916 ? _T_4702 : _T_3890_11; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_301 = _T_4916 ? _T_4704 : _T_3890_12; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_302 = _T_4916 ? _T_4706 : _T_3890_13; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_303 = _T_4916 ? _T_4708 : _T_3890_14; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_304 = _T_4916 ? _T_4710 : _T_3890_15; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_305 = _T_4916 ? _T_4712 : _T_3890_16; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_306 = _T_4916 ? _T_4714 : _T_3890_17; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_307 = _T_4916 ? _T_4716 : _T_3890_18; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_308 = _T_4916 ? _T_4718 : _T_3890_19; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_309 = _T_4916 ? _T_4720 : _T_3890_20; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_310 = _T_4916 ? _T_4722 : _T_3890_21; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_311 = _T_4916 ? _T_4724 : _T_3890_22; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_312 = _T_4916 ? _T_4726 : _T_3890_23; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_313 = _T_4916 ? _T_4728 : _T_3890_24; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_314 = _T_4916 ? _T_4730 : _T_3890_25; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_315 = _T_4916 ? _T_4732 : _T_3890_26; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_316 = _T_4916 ? _T_4734 : _T_3890_27; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_317 = _T_4916 ? _T_4736 : _T_3890_28; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_318 = _T_4916 ? _T_4738 : _T_3890_29; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_319 = _T_4916 ? _T_4740 : _T_3890_30; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_320 = _T_4916 ? _T_4742 : _T_3890_31; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_321 = _T_4916 ? _T_4744 : _T_3890_32; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_322 = _T_4916 ? _T_4746 : _T_3890_33; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_323 = _T_4916 ? _T_4748 : _T_3890_34; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_324 = _T_4916 ? _T_4750 : _T_3890_35; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_325 = _T_4916 ? _T_4752 : _T_3890_36; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_326 = _T_4916 ? _T_4754 : _T_3890_37; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_327 = _T_4916 ? _T_4756 : _T_3890_38; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_328 = _T_4916 ? _T_4758 : _T_3890_39; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_329 = _T_4916 ? _T_4760 : _T_3890_40; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_330 = _T_4916 ? _T_4762 : _T_3890_41; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_331 = _T_4916 ? _T_4764 : _T_3890_42; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_332 = _T_4916 ? _T_4766 : _T_3890_43; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_333 = _T_4916 ? _T_4768 : _T_3890_44; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_334 = _T_4916 ? _T_4770 : _T_3890_45; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_335 = _T_4916 ? _T_4772 : _T_3890_46; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_336 = _T_4916 ? _T_4774 : _T_3890_47; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_337 = _T_4916 ? _T_4776 : _T_3890_48; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_338 = _T_4916 ? _T_4778 : _T_3890_49; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_339 = _T_4916 ? _T_4780 : _T_3890_50; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_340 = _T_4916 ? _T_4782 : _T_3890_51; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_341 = _T_4916 ? _T_4784 : _T_3890_52; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_342 = _T_4916 ? _T_4786 : _T_3890_53; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_343 = _T_4916 ? _T_4788 : _T_3890_54; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_344 = _T_4916 ? _T_4790 : _T_3890_55; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_345 = _T_4916 ? _T_4792 : _T_3890_56; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_346 = _T_4916 ? _T_4794 : _T_3890_57; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_347 = _T_4916 ? _T_4796 : _T_3890_58; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_348 = _T_4916 ? _T_4798 : _T_3890_59; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_349 = _T_4916 ? _T_4800 : _T_3890_60; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_350 = _T_4916 ? _T_4802 : _T_3890_61; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_351 = _T_4916 ? _T_4804 : _T_3890_62; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_352 = _T_4916 ? _T_4806 : _T_3890_63; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_353 = _T_4916 ? _T_4917 : _T_4288_0; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_354 = _T_4916 ? _T_4918 : _T_4288_1; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_355 = _T_4916 ? _T_4919 : _T_4288_2; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_356 = _T_4916 ? _T_4920 : _T_4288_3; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_357 = _T_4916 ? _T_4921 : _T_4288_4; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_358 = _T_4916 ? _T_4922 : _T_4288_5; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_359 = _T_4916 ? _T_4923 : _T_4288_6; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_360 = _T_4916 ? _T_4924 : _T_4288_7; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_361 = _T_4916 ? _T_4925 : _T_4288_8; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_362 = _T_4916 ? _T_4926 : _T_4288_9; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_363 = _T_4916 ? _T_4927 : _T_4288_10; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_364 = _T_4916 ? _T_4928 : _T_4288_11; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_365 = _T_4916 ? _T_4929 : _T_4288_12; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_366 = _T_4916 ? _T_4930 : _T_4288_13; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_367 = _T_4916 ? _T_4931 : _T_4288_14; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign _GEN_368 = _T_4916 ? _T_4932 : _T_4288_15; // @[NV_NVDLA_CSC_wl.scala 816:52:@18838.4]
  assign io_sc2cdma_wt_updt_valid = _T_863; // @[NV_NVDLA_CSC_wl.scala 212:30:@16498.4]
  assign io_sc2cdma_wt_updt_bits_entries = _T_867; // @[NV_NVDLA_CSC_wl.scala 213:37:@16504.4]
  assign io_sc2cdma_wmb_entries = _T_871; // @[NV_NVDLA_CSC_wl.scala 214:28:@16510.4]
  assign io_sc2buf_wt_rd_addr_valid = _T_1631; // @[NV_NVDLA_CSC_wl.scala 631:32:@17189.4]
  assign io_sc2buf_wt_rd_addr_bits = _T_1634; // @[NV_NVDLA_CSC_wl.scala 632:31:@17190.4]
  assign io_sc2mac_wt_a_valid = _T_3157; // @[NV_NVDLA_CSC_wl.scala 829:26:@19337.4]
  assign io_sc2mac_wt_a_bits_sel_0 = _T_4161_0; // @[NV_NVDLA_CSC_wl.scala 833:29:@19467.4]
  assign io_sc2mac_wt_a_bits_sel_1 = _T_4161_1; // @[NV_NVDLA_CSC_wl.scala 833:29:@19468.4]
  assign io_sc2mac_wt_a_bits_sel_2 = _T_4161_2; // @[NV_NVDLA_CSC_wl.scala 833:29:@19469.4]
  assign io_sc2mac_wt_a_bits_sel_3 = _T_4161_3; // @[NV_NVDLA_CSC_wl.scala 833:29:@19470.4]
  assign io_sc2mac_wt_a_bits_sel_4 = _T_4161_4; // @[NV_NVDLA_CSC_wl.scala 833:29:@19471.4]
  assign io_sc2mac_wt_a_bits_sel_5 = _T_4161_5; // @[NV_NVDLA_CSC_wl.scala 833:29:@19472.4]
  assign io_sc2mac_wt_a_bits_sel_6 = _T_4161_6; // @[NV_NVDLA_CSC_wl.scala 833:29:@19473.4]
  assign io_sc2mac_wt_a_bits_sel_7 = _T_4161_7; // @[NV_NVDLA_CSC_wl.scala 833:29:@19474.4]
  assign io_sc2mac_wt_a_bits_sel_8 = _T_4161_8; // @[NV_NVDLA_CSC_wl.scala 833:29:@19475.4]
  assign io_sc2mac_wt_a_bits_sel_9 = _T_4161_9; // @[NV_NVDLA_CSC_wl.scala 833:29:@19476.4]
  assign io_sc2mac_wt_a_bits_sel_10 = _T_4161_10; // @[NV_NVDLA_CSC_wl.scala 833:29:@19477.4]
  assign io_sc2mac_wt_a_bits_sel_11 = _T_4161_11; // @[NV_NVDLA_CSC_wl.scala 833:29:@19478.4]
  assign io_sc2mac_wt_a_bits_sel_12 = _T_4161_12; // @[NV_NVDLA_CSC_wl.scala 833:29:@19479.4]
  assign io_sc2mac_wt_a_bits_sel_13 = _T_4161_13; // @[NV_NVDLA_CSC_wl.scala 833:29:@19480.4]
  assign io_sc2mac_wt_a_bits_sel_14 = _T_4161_14; // @[NV_NVDLA_CSC_wl.scala 833:29:@19481.4]
  assign io_sc2mac_wt_a_bits_sel_15 = _T_4161_15; // @[NV_NVDLA_CSC_wl.scala 833:29:@19482.4]
  assign io_sc2mac_wt_a_bits_mask_0 = _T_3427_0; // @[NV_NVDLA_CSC_wl.scala 831:30:@19339.4]
  assign io_sc2mac_wt_a_bits_mask_1 = _T_3427_1; // @[NV_NVDLA_CSC_wl.scala 831:30:@19340.4]
  assign io_sc2mac_wt_a_bits_mask_2 = _T_3427_2; // @[NV_NVDLA_CSC_wl.scala 831:30:@19341.4]
  assign io_sc2mac_wt_a_bits_mask_3 = _T_3427_3; // @[NV_NVDLA_CSC_wl.scala 831:30:@19342.4]
  assign io_sc2mac_wt_a_bits_mask_4 = _T_3427_4; // @[NV_NVDLA_CSC_wl.scala 831:30:@19343.4]
  assign io_sc2mac_wt_a_bits_mask_5 = _T_3427_5; // @[NV_NVDLA_CSC_wl.scala 831:30:@19344.4]
  assign io_sc2mac_wt_a_bits_mask_6 = _T_3427_6; // @[NV_NVDLA_CSC_wl.scala 831:30:@19345.4]
  assign io_sc2mac_wt_a_bits_mask_7 = _T_3427_7; // @[NV_NVDLA_CSC_wl.scala 831:30:@19346.4]
  assign io_sc2mac_wt_a_bits_mask_8 = _T_3427_8; // @[NV_NVDLA_CSC_wl.scala 831:30:@19347.4]
  assign io_sc2mac_wt_a_bits_mask_9 = _T_3427_9; // @[NV_NVDLA_CSC_wl.scala 831:30:@19348.4]
  assign io_sc2mac_wt_a_bits_mask_10 = _T_3427_10; // @[NV_NVDLA_CSC_wl.scala 831:30:@19349.4]
  assign io_sc2mac_wt_a_bits_mask_11 = _T_3427_11; // @[NV_NVDLA_CSC_wl.scala 831:30:@19350.4]
  assign io_sc2mac_wt_a_bits_mask_12 = _T_3427_12; // @[NV_NVDLA_CSC_wl.scala 831:30:@19351.4]
  assign io_sc2mac_wt_a_bits_mask_13 = _T_3427_13; // @[NV_NVDLA_CSC_wl.scala 831:30:@19352.4]
  assign io_sc2mac_wt_a_bits_mask_14 = _T_3427_14; // @[NV_NVDLA_CSC_wl.scala 831:30:@19353.4]
  assign io_sc2mac_wt_a_bits_mask_15 = _T_3427_15; // @[NV_NVDLA_CSC_wl.scala 831:30:@19354.4]
  assign io_sc2mac_wt_a_bits_mask_16 = _T_3427_16; // @[NV_NVDLA_CSC_wl.scala 831:30:@19355.4]
  assign io_sc2mac_wt_a_bits_mask_17 = _T_3427_17; // @[NV_NVDLA_CSC_wl.scala 831:30:@19356.4]
  assign io_sc2mac_wt_a_bits_mask_18 = _T_3427_18; // @[NV_NVDLA_CSC_wl.scala 831:30:@19357.4]
  assign io_sc2mac_wt_a_bits_mask_19 = _T_3427_19; // @[NV_NVDLA_CSC_wl.scala 831:30:@19358.4]
  assign io_sc2mac_wt_a_bits_mask_20 = _T_3427_20; // @[NV_NVDLA_CSC_wl.scala 831:30:@19359.4]
  assign io_sc2mac_wt_a_bits_mask_21 = _T_3427_21; // @[NV_NVDLA_CSC_wl.scala 831:30:@19360.4]
  assign io_sc2mac_wt_a_bits_mask_22 = _T_3427_22; // @[NV_NVDLA_CSC_wl.scala 831:30:@19361.4]
  assign io_sc2mac_wt_a_bits_mask_23 = _T_3427_23; // @[NV_NVDLA_CSC_wl.scala 831:30:@19362.4]
  assign io_sc2mac_wt_a_bits_mask_24 = _T_3427_24; // @[NV_NVDLA_CSC_wl.scala 831:30:@19363.4]
  assign io_sc2mac_wt_a_bits_mask_25 = _T_3427_25; // @[NV_NVDLA_CSC_wl.scala 831:30:@19364.4]
  assign io_sc2mac_wt_a_bits_mask_26 = _T_3427_26; // @[NV_NVDLA_CSC_wl.scala 831:30:@19365.4]
  assign io_sc2mac_wt_a_bits_mask_27 = _T_3427_27; // @[NV_NVDLA_CSC_wl.scala 831:30:@19366.4]
  assign io_sc2mac_wt_a_bits_mask_28 = _T_3427_28; // @[NV_NVDLA_CSC_wl.scala 831:30:@19367.4]
  assign io_sc2mac_wt_a_bits_mask_29 = _T_3427_29; // @[NV_NVDLA_CSC_wl.scala 831:30:@19368.4]
  assign io_sc2mac_wt_a_bits_mask_30 = _T_3427_30; // @[NV_NVDLA_CSC_wl.scala 831:30:@19369.4]
  assign io_sc2mac_wt_a_bits_mask_31 = _T_3427_31; // @[NV_NVDLA_CSC_wl.scala 831:30:@19370.4]
  assign io_sc2mac_wt_a_bits_mask_32 = _T_3427_32; // @[NV_NVDLA_CSC_wl.scala 831:30:@19371.4]
  assign io_sc2mac_wt_a_bits_mask_33 = _T_3427_33; // @[NV_NVDLA_CSC_wl.scala 831:30:@19372.4]
  assign io_sc2mac_wt_a_bits_mask_34 = _T_3427_34; // @[NV_NVDLA_CSC_wl.scala 831:30:@19373.4]
  assign io_sc2mac_wt_a_bits_mask_35 = _T_3427_35; // @[NV_NVDLA_CSC_wl.scala 831:30:@19374.4]
  assign io_sc2mac_wt_a_bits_mask_36 = _T_3427_36; // @[NV_NVDLA_CSC_wl.scala 831:30:@19375.4]
  assign io_sc2mac_wt_a_bits_mask_37 = _T_3427_37; // @[NV_NVDLA_CSC_wl.scala 831:30:@19376.4]
  assign io_sc2mac_wt_a_bits_mask_38 = _T_3427_38; // @[NV_NVDLA_CSC_wl.scala 831:30:@19377.4]
  assign io_sc2mac_wt_a_bits_mask_39 = _T_3427_39; // @[NV_NVDLA_CSC_wl.scala 831:30:@19378.4]
  assign io_sc2mac_wt_a_bits_mask_40 = _T_3427_40; // @[NV_NVDLA_CSC_wl.scala 831:30:@19379.4]
  assign io_sc2mac_wt_a_bits_mask_41 = _T_3427_41; // @[NV_NVDLA_CSC_wl.scala 831:30:@19380.4]
  assign io_sc2mac_wt_a_bits_mask_42 = _T_3427_42; // @[NV_NVDLA_CSC_wl.scala 831:30:@19381.4]
  assign io_sc2mac_wt_a_bits_mask_43 = _T_3427_43; // @[NV_NVDLA_CSC_wl.scala 831:30:@19382.4]
  assign io_sc2mac_wt_a_bits_mask_44 = _T_3427_44; // @[NV_NVDLA_CSC_wl.scala 831:30:@19383.4]
  assign io_sc2mac_wt_a_bits_mask_45 = _T_3427_45; // @[NV_NVDLA_CSC_wl.scala 831:30:@19384.4]
  assign io_sc2mac_wt_a_bits_mask_46 = _T_3427_46; // @[NV_NVDLA_CSC_wl.scala 831:30:@19385.4]
  assign io_sc2mac_wt_a_bits_mask_47 = _T_3427_47; // @[NV_NVDLA_CSC_wl.scala 831:30:@19386.4]
  assign io_sc2mac_wt_a_bits_mask_48 = _T_3427_48; // @[NV_NVDLA_CSC_wl.scala 831:30:@19387.4]
  assign io_sc2mac_wt_a_bits_mask_49 = _T_3427_49; // @[NV_NVDLA_CSC_wl.scala 831:30:@19388.4]
  assign io_sc2mac_wt_a_bits_mask_50 = _T_3427_50; // @[NV_NVDLA_CSC_wl.scala 831:30:@19389.4]
  assign io_sc2mac_wt_a_bits_mask_51 = _T_3427_51; // @[NV_NVDLA_CSC_wl.scala 831:30:@19390.4]
  assign io_sc2mac_wt_a_bits_mask_52 = _T_3427_52; // @[NV_NVDLA_CSC_wl.scala 831:30:@19391.4]
  assign io_sc2mac_wt_a_bits_mask_53 = _T_3427_53; // @[NV_NVDLA_CSC_wl.scala 831:30:@19392.4]
  assign io_sc2mac_wt_a_bits_mask_54 = _T_3427_54; // @[NV_NVDLA_CSC_wl.scala 831:30:@19393.4]
  assign io_sc2mac_wt_a_bits_mask_55 = _T_3427_55; // @[NV_NVDLA_CSC_wl.scala 831:30:@19394.4]
  assign io_sc2mac_wt_a_bits_mask_56 = _T_3427_56; // @[NV_NVDLA_CSC_wl.scala 831:30:@19395.4]
  assign io_sc2mac_wt_a_bits_mask_57 = _T_3427_57; // @[NV_NVDLA_CSC_wl.scala 831:30:@19396.4]
  assign io_sc2mac_wt_a_bits_mask_58 = _T_3427_58; // @[NV_NVDLA_CSC_wl.scala 831:30:@19397.4]
  assign io_sc2mac_wt_a_bits_mask_59 = _T_3427_59; // @[NV_NVDLA_CSC_wl.scala 831:30:@19398.4]
  assign io_sc2mac_wt_a_bits_mask_60 = _T_3427_60; // @[NV_NVDLA_CSC_wl.scala 831:30:@19399.4]
  assign io_sc2mac_wt_a_bits_mask_61 = _T_3427_61; // @[NV_NVDLA_CSC_wl.scala 831:30:@19400.4]
  assign io_sc2mac_wt_a_bits_mask_62 = _T_3427_62; // @[NV_NVDLA_CSC_wl.scala 831:30:@19401.4]
  assign io_sc2mac_wt_a_bits_mask_63 = _T_3427_63; // @[NV_NVDLA_CSC_wl.scala 831:30:@19402.4]
  assign io_sc2mac_wt_a_bits_data_0 = _T_4344_0; // @[NV_NVDLA_CSC_wl.scala 835:30:@19499.4]
  assign io_sc2mac_wt_a_bits_data_1 = _T_4344_1; // @[NV_NVDLA_CSC_wl.scala 835:30:@19500.4]
  assign io_sc2mac_wt_a_bits_data_2 = _T_4344_2; // @[NV_NVDLA_CSC_wl.scala 835:30:@19501.4]
  assign io_sc2mac_wt_a_bits_data_3 = _T_4344_3; // @[NV_NVDLA_CSC_wl.scala 835:30:@19502.4]
  assign io_sc2mac_wt_a_bits_data_4 = _T_4344_4; // @[NV_NVDLA_CSC_wl.scala 835:30:@19503.4]
  assign io_sc2mac_wt_a_bits_data_5 = _T_4344_5; // @[NV_NVDLA_CSC_wl.scala 835:30:@19504.4]
  assign io_sc2mac_wt_a_bits_data_6 = _T_4344_6; // @[NV_NVDLA_CSC_wl.scala 835:30:@19505.4]
  assign io_sc2mac_wt_a_bits_data_7 = _T_4344_7; // @[NV_NVDLA_CSC_wl.scala 835:30:@19506.4]
  assign io_sc2mac_wt_a_bits_data_8 = _T_4344_8; // @[NV_NVDLA_CSC_wl.scala 835:30:@19507.4]
  assign io_sc2mac_wt_a_bits_data_9 = _T_4344_9; // @[NV_NVDLA_CSC_wl.scala 835:30:@19508.4]
  assign io_sc2mac_wt_a_bits_data_10 = _T_4344_10; // @[NV_NVDLA_CSC_wl.scala 835:30:@19509.4]
  assign io_sc2mac_wt_a_bits_data_11 = _T_4344_11; // @[NV_NVDLA_CSC_wl.scala 835:30:@19510.4]
  assign io_sc2mac_wt_a_bits_data_12 = _T_4344_12; // @[NV_NVDLA_CSC_wl.scala 835:30:@19511.4]
  assign io_sc2mac_wt_a_bits_data_13 = _T_4344_13; // @[NV_NVDLA_CSC_wl.scala 835:30:@19512.4]
  assign io_sc2mac_wt_a_bits_data_14 = _T_4344_14; // @[NV_NVDLA_CSC_wl.scala 835:30:@19513.4]
  assign io_sc2mac_wt_a_bits_data_15 = _T_4344_15; // @[NV_NVDLA_CSC_wl.scala 835:30:@19514.4]
  assign io_sc2mac_wt_a_bits_data_16 = _T_4344_16; // @[NV_NVDLA_CSC_wl.scala 835:30:@19515.4]
  assign io_sc2mac_wt_a_bits_data_17 = _T_4344_17; // @[NV_NVDLA_CSC_wl.scala 835:30:@19516.4]
  assign io_sc2mac_wt_a_bits_data_18 = _T_4344_18; // @[NV_NVDLA_CSC_wl.scala 835:30:@19517.4]
  assign io_sc2mac_wt_a_bits_data_19 = _T_4344_19; // @[NV_NVDLA_CSC_wl.scala 835:30:@19518.4]
  assign io_sc2mac_wt_a_bits_data_20 = _T_4344_20; // @[NV_NVDLA_CSC_wl.scala 835:30:@19519.4]
  assign io_sc2mac_wt_a_bits_data_21 = _T_4344_21; // @[NV_NVDLA_CSC_wl.scala 835:30:@19520.4]
  assign io_sc2mac_wt_a_bits_data_22 = _T_4344_22; // @[NV_NVDLA_CSC_wl.scala 835:30:@19521.4]
  assign io_sc2mac_wt_a_bits_data_23 = _T_4344_23; // @[NV_NVDLA_CSC_wl.scala 835:30:@19522.4]
  assign io_sc2mac_wt_a_bits_data_24 = _T_4344_24; // @[NV_NVDLA_CSC_wl.scala 835:30:@19523.4]
  assign io_sc2mac_wt_a_bits_data_25 = _T_4344_25; // @[NV_NVDLA_CSC_wl.scala 835:30:@19524.4]
  assign io_sc2mac_wt_a_bits_data_26 = _T_4344_26; // @[NV_NVDLA_CSC_wl.scala 835:30:@19525.4]
  assign io_sc2mac_wt_a_bits_data_27 = _T_4344_27; // @[NV_NVDLA_CSC_wl.scala 835:30:@19526.4]
  assign io_sc2mac_wt_a_bits_data_28 = _T_4344_28; // @[NV_NVDLA_CSC_wl.scala 835:30:@19527.4]
  assign io_sc2mac_wt_a_bits_data_29 = _T_4344_29; // @[NV_NVDLA_CSC_wl.scala 835:30:@19528.4]
  assign io_sc2mac_wt_a_bits_data_30 = _T_4344_30; // @[NV_NVDLA_CSC_wl.scala 835:30:@19529.4]
  assign io_sc2mac_wt_a_bits_data_31 = _T_4344_31; // @[NV_NVDLA_CSC_wl.scala 835:30:@19530.4]
  assign io_sc2mac_wt_a_bits_data_32 = _T_4344_32; // @[NV_NVDLA_CSC_wl.scala 835:30:@19531.4]
  assign io_sc2mac_wt_a_bits_data_33 = _T_4344_33; // @[NV_NVDLA_CSC_wl.scala 835:30:@19532.4]
  assign io_sc2mac_wt_a_bits_data_34 = _T_4344_34; // @[NV_NVDLA_CSC_wl.scala 835:30:@19533.4]
  assign io_sc2mac_wt_a_bits_data_35 = _T_4344_35; // @[NV_NVDLA_CSC_wl.scala 835:30:@19534.4]
  assign io_sc2mac_wt_a_bits_data_36 = _T_4344_36; // @[NV_NVDLA_CSC_wl.scala 835:30:@19535.4]
  assign io_sc2mac_wt_a_bits_data_37 = _T_4344_37; // @[NV_NVDLA_CSC_wl.scala 835:30:@19536.4]
  assign io_sc2mac_wt_a_bits_data_38 = _T_4344_38; // @[NV_NVDLA_CSC_wl.scala 835:30:@19537.4]
  assign io_sc2mac_wt_a_bits_data_39 = _T_4344_39; // @[NV_NVDLA_CSC_wl.scala 835:30:@19538.4]
  assign io_sc2mac_wt_a_bits_data_40 = _T_4344_40; // @[NV_NVDLA_CSC_wl.scala 835:30:@19539.4]
  assign io_sc2mac_wt_a_bits_data_41 = _T_4344_41; // @[NV_NVDLA_CSC_wl.scala 835:30:@19540.4]
  assign io_sc2mac_wt_a_bits_data_42 = _T_4344_42; // @[NV_NVDLA_CSC_wl.scala 835:30:@19541.4]
  assign io_sc2mac_wt_a_bits_data_43 = _T_4344_43; // @[NV_NVDLA_CSC_wl.scala 835:30:@19542.4]
  assign io_sc2mac_wt_a_bits_data_44 = _T_4344_44; // @[NV_NVDLA_CSC_wl.scala 835:30:@19543.4]
  assign io_sc2mac_wt_a_bits_data_45 = _T_4344_45; // @[NV_NVDLA_CSC_wl.scala 835:30:@19544.4]
  assign io_sc2mac_wt_a_bits_data_46 = _T_4344_46; // @[NV_NVDLA_CSC_wl.scala 835:30:@19545.4]
  assign io_sc2mac_wt_a_bits_data_47 = _T_4344_47; // @[NV_NVDLA_CSC_wl.scala 835:30:@19546.4]
  assign io_sc2mac_wt_a_bits_data_48 = _T_4344_48; // @[NV_NVDLA_CSC_wl.scala 835:30:@19547.4]
  assign io_sc2mac_wt_a_bits_data_49 = _T_4344_49; // @[NV_NVDLA_CSC_wl.scala 835:30:@19548.4]
  assign io_sc2mac_wt_a_bits_data_50 = _T_4344_50; // @[NV_NVDLA_CSC_wl.scala 835:30:@19549.4]
  assign io_sc2mac_wt_a_bits_data_51 = _T_4344_51; // @[NV_NVDLA_CSC_wl.scala 835:30:@19550.4]
  assign io_sc2mac_wt_a_bits_data_52 = _T_4344_52; // @[NV_NVDLA_CSC_wl.scala 835:30:@19551.4]
  assign io_sc2mac_wt_a_bits_data_53 = _T_4344_53; // @[NV_NVDLA_CSC_wl.scala 835:30:@19552.4]
  assign io_sc2mac_wt_a_bits_data_54 = _T_4344_54; // @[NV_NVDLA_CSC_wl.scala 835:30:@19553.4]
  assign io_sc2mac_wt_a_bits_data_55 = _T_4344_55; // @[NV_NVDLA_CSC_wl.scala 835:30:@19554.4]
  assign io_sc2mac_wt_a_bits_data_56 = _T_4344_56; // @[NV_NVDLA_CSC_wl.scala 835:30:@19555.4]
  assign io_sc2mac_wt_a_bits_data_57 = _T_4344_57; // @[NV_NVDLA_CSC_wl.scala 835:30:@19556.4]
  assign io_sc2mac_wt_a_bits_data_58 = _T_4344_58; // @[NV_NVDLA_CSC_wl.scala 835:30:@19557.4]
  assign io_sc2mac_wt_a_bits_data_59 = _T_4344_59; // @[NV_NVDLA_CSC_wl.scala 835:30:@19558.4]
  assign io_sc2mac_wt_a_bits_data_60 = _T_4344_60; // @[NV_NVDLA_CSC_wl.scala 835:30:@19559.4]
  assign io_sc2mac_wt_a_bits_data_61 = _T_4344_61; // @[NV_NVDLA_CSC_wl.scala 835:30:@19560.4]
  assign io_sc2mac_wt_a_bits_data_62 = _T_4344_62; // @[NV_NVDLA_CSC_wl.scala 835:30:@19561.4]
  assign io_sc2mac_wt_a_bits_data_63 = _T_4344_63; // @[NV_NVDLA_CSC_wl.scala 835:30:@19562.4]
  assign io_sc2mac_wt_b_valid = _T_3160; // @[NV_NVDLA_CSC_wl.scala 830:26:@19338.4]
  assign io_sc2mac_wt_b_bits_sel_0 = _T_4288_0; // @[NV_NVDLA_CSC_wl.scala 834:29:@19483.4]
  assign io_sc2mac_wt_b_bits_sel_1 = _T_4288_1; // @[NV_NVDLA_CSC_wl.scala 834:29:@19484.4]
  assign io_sc2mac_wt_b_bits_sel_2 = _T_4288_2; // @[NV_NVDLA_CSC_wl.scala 834:29:@19485.4]
  assign io_sc2mac_wt_b_bits_sel_3 = _T_4288_3; // @[NV_NVDLA_CSC_wl.scala 834:29:@19486.4]
  assign io_sc2mac_wt_b_bits_sel_4 = _T_4288_4; // @[NV_NVDLA_CSC_wl.scala 834:29:@19487.4]
  assign io_sc2mac_wt_b_bits_sel_5 = _T_4288_5; // @[NV_NVDLA_CSC_wl.scala 834:29:@19488.4]
  assign io_sc2mac_wt_b_bits_sel_6 = _T_4288_6; // @[NV_NVDLA_CSC_wl.scala 834:29:@19489.4]
  assign io_sc2mac_wt_b_bits_sel_7 = _T_4288_7; // @[NV_NVDLA_CSC_wl.scala 834:29:@19490.4]
  assign io_sc2mac_wt_b_bits_sel_8 = _T_4288_8; // @[NV_NVDLA_CSC_wl.scala 834:29:@19491.4]
  assign io_sc2mac_wt_b_bits_sel_9 = _T_4288_9; // @[NV_NVDLA_CSC_wl.scala 834:29:@19492.4]
  assign io_sc2mac_wt_b_bits_sel_10 = _T_4288_10; // @[NV_NVDLA_CSC_wl.scala 834:29:@19493.4]
  assign io_sc2mac_wt_b_bits_sel_11 = _T_4288_11; // @[NV_NVDLA_CSC_wl.scala 834:29:@19494.4]
  assign io_sc2mac_wt_b_bits_sel_12 = _T_4288_12; // @[NV_NVDLA_CSC_wl.scala 834:29:@19495.4]
  assign io_sc2mac_wt_b_bits_sel_13 = _T_4288_13; // @[NV_NVDLA_CSC_wl.scala 834:29:@19496.4]
  assign io_sc2mac_wt_b_bits_sel_14 = _T_4288_14; // @[NV_NVDLA_CSC_wl.scala 834:29:@19497.4]
  assign io_sc2mac_wt_b_bits_sel_15 = _T_4288_15; // @[NV_NVDLA_CSC_wl.scala 834:29:@19498.4]
  assign io_sc2mac_wt_b_bits_mask_0 = _T_3890_0; // @[NV_NVDLA_CSC_wl.scala 832:30:@19403.4]
  assign io_sc2mac_wt_b_bits_mask_1 = _T_3890_1; // @[NV_NVDLA_CSC_wl.scala 832:30:@19404.4]
  assign io_sc2mac_wt_b_bits_mask_2 = _T_3890_2; // @[NV_NVDLA_CSC_wl.scala 832:30:@19405.4]
  assign io_sc2mac_wt_b_bits_mask_3 = _T_3890_3; // @[NV_NVDLA_CSC_wl.scala 832:30:@19406.4]
  assign io_sc2mac_wt_b_bits_mask_4 = _T_3890_4; // @[NV_NVDLA_CSC_wl.scala 832:30:@19407.4]
  assign io_sc2mac_wt_b_bits_mask_5 = _T_3890_5; // @[NV_NVDLA_CSC_wl.scala 832:30:@19408.4]
  assign io_sc2mac_wt_b_bits_mask_6 = _T_3890_6; // @[NV_NVDLA_CSC_wl.scala 832:30:@19409.4]
  assign io_sc2mac_wt_b_bits_mask_7 = _T_3890_7; // @[NV_NVDLA_CSC_wl.scala 832:30:@19410.4]
  assign io_sc2mac_wt_b_bits_mask_8 = _T_3890_8; // @[NV_NVDLA_CSC_wl.scala 832:30:@19411.4]
  assign io_sc2mac_wt_b_bits_mask_9 = _T_3890_9; // @[NV_NVDLA_CSC_wl.scala 832:30:@19412.4]
  assign io_sc2mac_wt_b_bits_mask_10 = _T_3890_10; // @[NV_NVDLA_CSC_wl.scala 832:30:@19413.4]
  assign io_sc2mac_wt_b_bits_mask_11 = _T_3890_11; // @[NV_NVDLA_CSC_wl.scala 832:30:@19414.4]
  assign io_sc2mac_wt_b_bits_mask_12 = _T_3890_12; // @[NV_NVDLA_CSC_wl.scala 832:30:@19415.4]
  assign io_sc2mac_wt_b_bits_mask_13 = _T_3890_13; // @[NV_NVDLA_CSC_wl.scala 832:30:@19416.4]
  assign io_sc2mac_wt_b_bits_mask_14 = _T_3890_14; // @[NV_NVDLA_CSC_wl.scala 832:30:@19417.4]
  assign io_sc2mac_wt_b_bits_mask_15 = _T_3890_15; // @[NV_NVDLA_CSC_wl.scala 832:30:@19418.4]
  assign io_sc2mac_wt_b_bits_mask_16 = _T_3890_16; // @[NV_NVDLA_CSC_wl.scala 832:30:@19419.4]
  assign io_sc2mac_wt_b_bits_mask_17 = _T_3890_17; // @[NV_NVDLA_CSC_wl.scala 832:30:@19420.4]
  assign io_sc2mac_wt_b_bits_mask_18 = _T_3890_18; // @[NV_NVDLA_CSC_wl.scala 832:30:@19421.4]
  assign io_sc2mac_wt_b_bits_mask_19 = _T_3890_19; // @[NV_NVDLA_CSC_wl.scala 832:30:@19422.4]
  assign io_sc2mac_wt_b_bits_mask_20 = _T_3890_20; // @[NV_NVDLA_CSC_wl.scala 832:30:@19423.4]
  assign io_sc2mac_wt_b_bits_mask_21 = _T_3890_21; // @[NV_NVDLA_CSC_wl.scala 832:30:@19424.4]
  assign io_sc2mac_wt_b_bits_mask_22 = _T_3890_22; // @[NV_NVDLA_CSC_wl.scala 832:30:@19425.4]
  assign io_sc2mac_wt_b_bits_mask_23 = _T_3890_23; // @[NV_NVDLA_CSC_wl.scala 832:30:@19426.4]
  assign io_sc2mac_wt_b_bits_mask_24 = _T_3890_24; // @[NV_NVDLA_CSC_wl.scala 832:30:@19427.4]
  assign io_sc2mac_wt_b_bits_mask_25 = _T_3890_25; // @[NV_NVDLA_CSC_wl.scala 832:30:@19428.4]
  assign io_sc2mac_wt_b_bits_mask_26 = _T_3890_26; // @[NV_NVDLA_CSC_wl.scala 832:30:@19429.4]
  assign io_sc2mac_wt_b_bits_mask_27 = _T_3890_27; // @[NV_NVDLA_CSC_wl.scala 832:30:@19430.4]
  assign io_sc2mac_wt_b_bits_mask_28 = _T_3890_28; // @[NV_NVDLA_CSC_wl.scala 832:30:@19431.4]
  assign io_sc2mac_wt_b_bits_mask_29 = _T_3890_29; // @[NV_NVDLA_CSC_wl.scala 832:30:@19432.4]
  assign io_sc2mac_wt_b_bits_mask_30 = _T_3890_30; // @[NV_NVDLA_CSC_wl.scala 832:30:@19433.4]
  assign io_sc2mac_wt_b_bits_mask_31 = _T_3890_31; // @[NV_NVDLA_CSC_wl.scala 832:30:@19434.4]
  assign io_sc2mac_wt_b_bits_mask_32 = _T_3890_32; // @[NV_NVDLA_CSC_wl.scala 832:30:@19435.4]
  assign io_sc2mac_wt_b_bits_mask_33 = _T_3890_33; // @[NV_NVDLA_CSC_wl.scala 832:30:@19436.4]
  assign io_sc2mac_wt_b_bits_mask_34 = _T_3890_34; // @[NV_NVDLA_CSC_wl.scala 832:30:@19437.4]
  assign io_sc2mac_wt_b_bits_mask_35 = _T_3890_35; // @[NV_NVDLA_CSC_wl.scala 832:30:@19438.4]
  assign io_sc2mac_wt_b_bits_mask_36 = _T_3890_36; // @[NV_NVDLA_CSC_wl.scala 832:30:@19439.4]
  assign io_sc2mac_wt_b_bits_mask_37 = _T_3890_37; // @[NV_NVDLA_CSC_wl.scala 832:30:@19440.4]
  assign io_sc2mac_wt_b_bits_mask_38 = _T_3890_38; // @[NV_NVDLA_CSC_wl.scala 832:30:@19441.4]
  assign io_sc2mac_wt_b_bits_mask_39 = _T_3890_39; // @[NV_NVDLA_CSC_wl.scala 832:30:@19442.4]
  assign io_sc2mac_wt_b_bits_mask_40 = _T_3890_40; // @[NV_NVDLA_CSC_wl.scala 832:30:@19443.4]
  assign io_sc2mac_wt_b_bits_mask_41 = _T_3890_41; // @[NV_NVDLA_CSC_wl.scala 832:30:@19444.4]
  assign io_sc2mac_wt_b_bits_mask_42 = _T_3890_42; // @[NV_NVDLA_CSC_wl.scala 832:30:@19445.4]
  assign io_sc2mac_wt_b_bits_mask_43 = _T_3890_43; // @[NV_NVDLA_CSC_wl.scala 832:30:@19446.4]
  assign io_sc2mac_wt_b_bits_mask_44 = _T_3890_44; // @[NV_NVDLA_CSC_wl.scala 832:30:@19447.4]
  assign io_sc2mac_wt_b_bits_mask_45 = _T_3890_45; // @[NV_NVDLA_CSC_wl.scala 832:30:@19448.4]
  assign io_sc2mac_wt_b_bits_mask_46 = _T_3890_46; // @[NV_NVDLA_CSC_wl.scala 832:30:@19449.4]
  assign io_sc2mac_wt_b_bits_mask_47 = _T_3890_47; // @[NV_NVDLA_CSC_wl.scala 832:30:@19450.4]
  assign io_sc2mac_wt_b_bits_mask_48 = _T_3890_48; // @[NV_NVDLA_CSC_wl.scala 832:30:@19451.4]
  assign io_sc2mac_wt_b_bits_mask_49 = _T_3890_49; // @[NV_NVDLA_CSC_wl.scala 832:30:@19452.4]
  assign io_sc2mac_wt_b_bits_mask_50 = _T_3890_50; // @[NV_NVDLA_CSC_wl.scala 832:30:@19453.4]
  assign io_sc2mac_wt_b_bits_mask_51 = _T_3890_51; // @[NV_NVDLA_CSC_wl.scala 832:30:@19454.4]
  assign io_sc2mac_wt_b_bits_mask_52 = _T_3890_52; // @[NV_NVDLA_CSC_wl.scala 832:30:@19455.4]
  assign io_sc2mac_wt_b_bits_mask_53 = _T_3890_53; // @[NV_NVDLA_CSC_wl.scala 832:30:@19456.4]
  assign io_sc2mac_wt_b_bits_mask_54 = _T_3890_54; // @[NV_NVDLA_CSC_wl.scala 832:30:@19457.4]
  assign io_sc2mac_wt_b_bits_mask_55 = _T_3890_55; // @[NV_NVDLA_CSC_wl.scala 832:30:@19458.4]
  assign io_sc2mac_wt_b_bits_mask_56 = _T_3890_56; // @[NV_NVDLA_CSC_wl.scala 832:30:@19459.4]
  assign io_sc2mac_wt_b_bits_mask_57 = _T_3890_57; // @[NV_NVDLA_CSC_wl.scala 832:30:@19460.4]
  assign io_sc2mac_wt_b_bits_mask_58 = _T_3890_58; // @[NV_NVDLA_CSC_wl.scala 832:30:@19461.4]
  assign io_sc2mac_wt_b_bits_mask_59 = _T_3890_59; // @[NV_NVDLA_CSC_wl.scala 832:30:@19462.4]
  assign io_sc2mac_wt_b_bits_mask_60 = _T_3890_60; // @[NV_NVDLA_CSC_wl.scala 832:30:@19463.4]
  assign io_sc2mac_wt_b_bits_mask_61 = _T_3890_61; // @[NV_NVDLA_CSC_wl.scala 832:30:@19464.4]
  assign io_sc2mac_wt_b_bits_mask_62 = _T_3890_62; // @[NV_NVDLA_CSC_wl.scala 832:30:@19465.4]
  assign io_sc2mac_wt_b_bits_mask_63 = _T_3890_63; // @[NV_NVDLA_CSC_wl.scala 832:30:@19466.4]
  assign io_sc2mac_wt_b_bits_data_0 = _T_4414_0; // @[NV_NVDLA_CSC_wl.scala 836:30:@19563.4]
  assign io_sc2mac_wt_b_bits_data_1 = _T_4414_1; // @[NV_NVDLA_CSC_wl.scala 836:30:@19564.4]
  assign io_sc2mac_wt_b_bits_data_2 = _T_4414_2; // @[NV_NVDLA_CSC_wl.scala 836:30:@19565.4]
  assign io_sc2mac_wt_b_bits_data_3 = _T_4414_3; // @[NV_NVDLA_CSC_wl.scala 836:30:@19566.4]
  assign io_sc2mac_wt_b_bits_data_4 = _T_4414_4; // @[NV_NVDLA_CSC_wl.scala 836:30:@19567.4]
  assign io_sc2mac_wt_b_bits_data_5 = _T_4414_5; // @[NV_NVDLA_CSC_wl.scala 836:30:@19568.4]
  assign io_sc2mac_wt_b_bits_data_6 = _T_4414_6; // @[NV_NVDLA_CSC_wl.scala 836:30:@19569.4]
  assign io_sc2mac_wt_b_bits_data_7 = _T_4414_7; // @[NV_NVDLA_CSC_wl.scala 836:30:@19570.4]
  assign io_sc2mac_wt_b_bits_data_8 = _T_4414_8; // @[NV_NVDLA_CSC_wl.scala 836:30:@19571.4]
  assign io_sc2mac_wt_b_bits_data_9 = _T_4414_9; // @[NV_NVDLA_CSC_wl.scala 836:30:@19572.4]
  assign io_sc2mac_wt_b_bits_data_10 = _T_4414_10; // @[NV_NVDLA_CSC_wl.scala 836:30:@19573.4]
  assign io_sc2mac_wt_b_bits_data_11 = _T_4414_11; // @[NV_NVDLA_CSC_wl.scala 836:30:@19574.4]
  assign io_sc2mac_wt_b_bits_data_12 = _T_4414_12; // @[NV_NVDLA_CSC_wl.scala 836:30:@19575.4]
  assign io_sc2mac_wt_b_bits_data_13 = _T_4414_13; // @[NV_NVDLA_CSC_wl.scala 836:30:@19576.4]
  assign io_sc2mac_wt_b_bits_data_14 = _T_4414_14; // @[NV_NVDLA_CSC_wl.scala 836:30:@19577.4]
  assign io_sc2mac_wt_b_bits_data_15 = _T_4414_15; // @[NV_NVDLA_CSC_wl.scala 836:30:@19578.4]
  assign io_sc2mac_wt_b_bits_data_16 = _T_4414_16; // @[NV_NVDLA_CSC_wl.scala 836:30:@19579.4]
  assign io_sc2mac_wt_b_bits_data_17 = _T_4414_17; // @[NV_NVDLA_CSC_wl.scala 836:30:@19580.4]
  assign io_sc2mac_wt_b_bits_data_18 = _T_4414_18; // @[NV_NVDLA_CSC_wl.scala 836:30:@19581.4]
  assign io_sc2mac_wt_b_bits_data_19 = _T_4414_19; // @[NV_NVDLA_CSC_wl.scala 836:30:@19582.4]
  assign io_sc2mac_wt_b_bits_data_20 = _T_4414_20; // @[NV_NVDLA_CSC_wl.scala 836:30:@19583.4]
  assign io_sc2mac_wt_b_bits_data_21 = _T_4414_21; // @[NV_NVDLA_CSC_wl.scala 836:30:@19584.4]
  assign io_sc2mac_wt_b_bits_data_22 = _T_4414_22; // @[NV_NVDLA_CSC_wl.scala 836:30:@19585.4]
  assign io_sc2mac_wt_b_bits_data_23 = _T_4414_23; // @[NV_NVDLA_CSC_wl.scala 836:30:@19586.4]
  assign io_sc2mac_wt_b_bits_data_24 = _T_4414_24; // @[NV_NVDLA_CSC_wl.scala 836:30:@19587.4]
  assign io_sc2mac_wt_b_bits_data_25 = _T_4414_25; // @[NV_NVDLA_CSC_wl.scala 836:30:@19588.4]
  assign io_sc2mac_wt_b_bits_data_26 = _T_4414_26; // @[NV_NVDLA_CSC_wl.scala 836:30:@19589.4]
  assign io_sc2mac_wt_b_bits_data_27 = _T_4414_27; // @[NV_NVDLA_CSC_wl.scala 836:30:@19590.4]
  assign io_sc2mac_wt_b_bits_data_28 = _T_4414_28; // @[NV_NVDLA_CSC_wl.scala 836:30:@19591.4]
  assign io_sc2mac_wt_b_bits_data_29 = _T_4414_29; // @[NV_NVDLA_CSC_wl.scala 836:30:@19592.4]
  assign io_sc2mac_wt_b_bits_data_30 = _T_4414_30; // @[NV_NVDLA_CSC_wl.scala 836:30:@19593.4]
  assign io_sc2mac_wt_b_bits_data_31 = _T_4414_31; // @[NV_NVDLA_CSC_wl.scala 836:30:@19594.4]
  assign io_sc2mac_wt_b_bits_data_32 = _T_4414_32; // @[NV_NVDLA_CSC_wl.scala 836:30:@19595.4]
  assign io_sc2mac_wt_b_bits_data_33 = _T_4414_33; // @[NV_NVDLA_CSC_wl.scala 836:30:@19596.4]
  assign io_sc2mac_wt_b_bits_data_34 = _T_4414_34; // @[NV_NVDLA_CSC_wl.scala 836:30:@19597.4]
  assign io_sc2mac_wt_b_bits_data_35 = _T_4414_35; // @[NV_NVDLA_CSC_wl.scala 836:30:@19598.4]
  assign io_sc2mac_wt_b_bits_data_36 = _T_4414_36; // @[NV_NVDLA_CSC_wl.scala 836:30:@19599.4]
  assign io_sc2mac_wt_b_bits_data_37 = _T_4414_37; // @[NV_NVDLA_CSC_wl.scala 836:30:@19600.4]
  assign io_sc2mac_wt_b_bits_data_38 = _T_4414_38; // @[NV_NVDLA_CSC_wl.scala 836:30:@19601.4]
  assign io_sc2mac_wt_b_bits_data_39 = _T_4414_39; // @[NV_NVDLA_CSC_wl.scala 836:30:@19602.4]
  assign io_sc2mac_wt_b_bits_data_40 = _T_4414_40; // @[NV_NVDLA_CSC_wl.scala 836:30:@19603.4]
  assign io_sc2mac_wt_b_bits_data_41 = _T_4414_41; // @[NV_NVDLA_CSC_wl.scala 836:30:@19604.4]
  assign io_sc2mac_wt_b_bits_data_42 = _T_4414_42; // @[NV_NVDLA_CSC_wl.scala 836:30:@19605.4]
  assign io_sc2mac_wt_b_bits_data_43 = _T_4414_43; // @[NV_NVDLA_CSC_wl.scala 836:30:@19606.4]
  assign io_sc2mac_wt_b_bits_data_44 = _T_4414_44; // @[NV_NVDLA_CSC_wl.scala 836:30:@19607.4]
  assign io_sc2mac_wt_b_bits_data_45 = _T_4414_45; // @[NV_NVDLA_CSC_wl.scala 836:30:@19608.4]
  assign io_sc2mac_wt_b_bits_data_46 = _T_4414_46; // @[NV_NVDLA_CSC_wl.scala 836:30:@19609.4]
  assign io_sc2mac_wt_b_bits_data_47 = _T_4414_47; // @[NV_NVDLA_CSC_wl.scala 836:30:@19610.4]
  assign io_sc2mac_wt_b_bits_data_48 = _T_4414_48; // @[NV_NVDLA_CSC_wl.scala 836:30:@19611.4]
  assign io_sc2mac_wt_b_bits_data_49 = _T_4414_49; // @[NV_NVDLA_CSC_wl.scala 836:30:@19612.4]
  assign io_sc2mac_wt_b_bits_data_50 = _T_4414_50; // @[NV_NVDLA_CSC_wl.scala 836:30:@19613.4]
  assign io_sc2mac_wt_b_bits_data_51 = _T_4414_51; // @[NV_NVDLA_CSC_wl.scala 836:30:@19614.4]
  assign io_sc2mac_wt_b_bits_data_52 = _T_4414_52; // @[NV_NVDLA_CSC_wl.scala 836:30:@19615.4]
  assign io_sc2mac_wt_b_bits_data_53 = _T_4414_53; // @[NV_NVDLA_CSC_wl.scala 836:30:@19616.4]
  assign io_sc2mac_wt_b_bits_data_54 = _T_4414_54; // @[NV_NVDLA_CSC_wl.scala 836:30:@19617.4]
  assign io_sc2mac_wt_b_bits_data_55 = _T_4414_55; // @[NV_NVDLA_CSC_wl.scala 836:30:@19618.4]
  assign io_sc2mac_wt_b_bits_data_56 = _T_4414_56; // @[NV_NVDLA_CSC_wl.scala 836:30:@19619.4]
  assign io_sc2mac_wt_b_bits_data_57 = _T_4414_57; // @[NV_NVDLA_CSC_wl.scala 836:30:@19620.4]
  assign io_sc2mac_wt_b_bits_data_58 = _T_4414_58; // @[NV_NVDLA_CSC_wl.scala 836:30:@19621.4]
  assign io_sc2mac_wt_b_bits_data_59 = _T_4414_59; // @[NV_NVDLA_CSC_wl.scala 836:30:@19622.4]
  assign io_sc2mac_wt_b_bits_data_60 = _T_4414_60; // @[NV_NVDLA_CSC_wl.scala 836:30:@19623.4]
  assign io_sc2mac_wt_b_bits_data_61 = _T_4414_61; // @[NV_NVDLA_CSC_wl.scala 836:30:@19624.4]
  assign io_sc2mac_wt_b_bits_data_62 = _T_4414_62; // @[NV_NVDLA_CSC_wl.scala 836:30:@19625.4]
  assign io_sc2mac_wt_b_bits_data_63 = _T_4414_63; // @[NV_NVDLA_CSC_wl.scala 836:30:@19626.4]
  assign NV_NVDLA_CSC_WL_dec_reset = reset; // @[:@17925.4]
  assign NV_NVDLA_CSC_WL_dec_io_nvdla_core_clk = io_nvdla_core_clk; // @[NV_NVDLA_CSC_wl.scala 779:29:@17926.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_valid = _T_2472; // @[NV_NVDLA_CSC_wl.scala 783:26:@18056.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_0 = _T_2739_0; // @[NV_NVDLA_CSC_wl.scala 781:30:@17991.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_1 = _T_2739_1; // @[NV_NVDLA_CSC_wl.scala 781:30:@17992.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_2 = _T_2739_2; // @[NV_NVDLA_CSC_wl.scala 781:30:@17993.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_3 = _T_2739_3; // @[NV_NVDLA_CSC_wl.scala 781:30:@17994.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_4 = _T_2739_4; // @[NV_NVDLA_CSC_wl.scala 781:30:@17995.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_5 = _T_2739_5; // @[NV_NVDLA_CSC_wl.scala 781:30:@17996.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_6 = _T_2739_6; // @[NV_NVDLA_CSC_wl.scala 781:30:@17997.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_7 = _T_2739_7; // @[NV_NVDLA_CSC_wl.scala 781:30:@17998.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_8 = _T_2739_8; // @[NV_NVDLA_CSC_wl.scala 781:30:@17999.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_9 = _T_2739_9; // @[NV_NVDLA_CSC_wl.scala 781:30:@18000.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_10 = _T_2739_10; // @[NV_NVDLA_CSC_wl.scala 781:30:@18001.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_11 = _T_2739_11; // @[NV_NVDLA_CSC_wl.scala 781:30:@18002.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_12 = _T_2739_12; // @[NV_NVDLA_CSC_wl.scala 781:30:@18003.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_13 = _T_2739_13; // @[NV_NVDLA_CSC_wl.scala 781:30:@18004.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_14 = _T_2739_14; // @[NV_NVDLA_CSC_wl.scala 781:30:@18005.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_15 = _T_2739_15; // @[NV_NVDLA_CSC_wl.scala 781:30:@18006.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_16 = _T_2739_16; // @[NV_NVDLA_CSC_wl.scala 781:30:@18007.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_17 = _T_2739_17; // @[NV_NVDLA_CSC_wl.scala 781:30:@18008.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_18 = _T_2739_18; // @[NV_NVDLA_CSC_wl.scala 781:30:@18009.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_19 = _T_2739_19; // @[NV_NVDLA_CSC_wl.scala 781:30:@18010.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_20 = _T_2739_20; // @[NV_NVDLA_CSC_wl.scala 781:30:@18011.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_21 = _T_2739_21; // @[NV_NVDLA_CSC_wl.scala 781:30:@18012.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_22 = _T_2739_22; // @[NV_NVDLA_CSC_wl.scala 781:30:@18013.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_23 = _T_2739_23; // @[NV_NVDLA_CSC_wl.scala 781:30:@18014.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_24 = _T_2739_24; // @[NV_NVDLA_CSC_wl.scala 781:30:@18015.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_25 = _T_2739_25; // @[NV_NVDLA_CSC_wl.scala 781:30:@18016.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_26 = _T_2739_26; // @[NV_NVDLA_CSC_wl.scala 781:30:@18017.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_27 = _T_2739_27; // @[NV_NVDLA_CSC_wl.scala 781:30:@18018.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_28 = _T_2739_28; // @[NV_NVDLA_CSC_wl.scala 781:30:@18019.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_29 = _T_2739_29; // @[NV_NVDLA_CSC_wl.scala 781:30:@18020.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_30 = _T_2739_30; // @[NV_NVDLA_CSC_wl.scala 781:30:@18021.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_31 = _T_2739_31; // @[NV_NVDLA_CSC_wl.scala 781:30:@18022.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_32 = _T_2739_32; // @[NV_NVDLA_CSC_wl.scala 781:30:@18023.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_33 = _T_2739_33; // @[NV_NVDLA_CSC_wl.scala 781:30:@18024.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_34 = _T_2739_34; // @[NV_NVDLA_CSC_wl.scala 781:30:@18025.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_35 = _T_2739_35; // @[NV_NVDLA_CSC_wl.scala 781:30:@18026.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_36 = _T_2739_36; // @[NV_NVDLA_CSC_wl.scala 781:30:@18027.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_37 = _T_2739_37; // @[NV_NVDLA_CSC_wl.scala 781:30:@18028.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_38 = _T_2739_38; // @[NV_NVDLA_CSC_wl.scala 781:30:@18029.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_39 = _T_2739_39; // @[NV_NVDLA_CSC_wl.scala 781:30:@18030.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_40 = _T_2739_40; // @[NV_NVDLA_CSC_wl.scala 781:30:@18031.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_41 = _T_2739_41; // @[NV_NVDLA_CSC_wl.scala 781:30:@18032.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_42 = _T_2739_42; // @[NV_NVDLA_CSC_wl.scala 781:30:@18033.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_43 = _T_2739_43; // @[NV_NVDLA_CSC_wl.scala 781:30:@18034.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_44 = _T_2739_44; // @[NV_NVDLA_CSC_wl.scala 781:30:@18035.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_45 = _T_2739_45; // @[NV_NVDLA_CSC_wl.scala 781:30:@18036.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_46 = _T_2739_46; // @[NV_NVDLA_CSC_wl.scala 781:30:@18037.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_47 = _T_2739_47; // @[NV_NVDLA_CSC_wl.scala 781:30:@18038.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_48 = _T_2739_48; // @[NV_NVDLA_CSC_wl.scala 781:30:@18039.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_49 = _T_2739_49; // @[NV_NVDLA_CSC_wl.scala 781:30:@18040.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_50 = _T_2739_50; // @[NV_NVDLA_CSC_wl.scala 781:30:@18041.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_51 = _T_2739_51; // @[NV_NVDLA_CSC_wl.scala 781:30:@18042.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_52 = _T_2739_52; // @[NV_NVDLA_CSC_wl.scala 781:30:@18043.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_53 = _T_2739_53; // @[NV_NVDLA_CSC_wl.scala 781:30:@18044.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_54 = _T_2739_54; // @[NV_NVDLA_CSC_wl.scala 781:30:@18045.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_55 = _T_2739_55; // @[NV_NVDLA_CSC_wl.scala 781:30:@18046.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_56 = _T_2739_56; // @[NV_NVDLA_CSC_wl.scala 781:30:@18047.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_57 = _T_2739_57; // @[NV_NVDLA_CSC_wl.scala 781:30:@18048.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_58 = _T_2739_58; // @[NV_NVDLA_CSC_wl.scala 781:30:@18049.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_59 = _T_2739_59; // @[NV_NVDLA_CSC_wl.scala 781:30:@18050.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_60 = _T_2739_60; // @[NV_NVDLA_CSC_wl.scala 781:30:@18051.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_61 = _T_2739_61; // @[NV_NVDLA_CSC_wl.scala 781:30:@18052.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_62 = _T_2739_62; // @[NV_NVDLA_CSC_wl.scala 781:30:@18053.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_63 = _T_2739_63; // @[NV_NVDLA_CSC_wl.scala 781:30:@18054.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_0 = _T_2095_0; // @[NV_NVDLA_CSC_wl.scala 780:30:@17927.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_1 = _T_2095_1; // @[NV_NVDLA_CSC_wl.scala 780:30:@17928.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_2 = _T_2095_2; // @[NV_NVDLA_CSC_wl.scala 780:30:@17929.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_3 = _T_2095_3; // @[NV_NVDLA_CSC_wl.scala 780:30:@17930.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_4 = _T_2095_4; // @[NV_NVDLA_CSC_wl.scala 780:30:@17931.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_5 = _T_2095_5; // @[NV_NVDLA_CSC_wl.scala 780:30:@17932.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_6 = _T_2095_6; // @[NV_NVDLA_CSC_wl.scala 780:30:@17933.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_7 = _T_2095_7; // @[NV_NVDLA_CSC_wl.scala 780:30:@17934.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_8 = _T_2095_8; // @[NV_NVDLA_CSC_wl.scala 780:30:@17935.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_9 = _T_2095_9; // @[NV_NVDLA_CSC_wl.scala 780:30:@17936.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_10 = _T_2095_10; // @[NV_NVDLA_CSC_wl.scala 780:30:@17937.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_11 = _T_2095_11; // @[NV_NVDLA_CSC_wl.scala 780:30:@17938.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_12 = _T_2095_12; // @[NV_NVDLA_CSC_wl.scala 780:30:@17939.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_13 = _T_2095_13; // @[NV_NVDLA_CSC_wl.scala 780:30:@17940.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_14 = _T_2095_14; // @[NV_NVDLA_CSC_wl.scala 780:30:@17941.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_15 = _T_2095_15; // @[NV_NVDLA_CSC_wl.scala 780:30:@17942.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_16 = _T_2095_16; // @[NV_NVDLA_CSC_wl.scala 780:30:@17943.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_17 = _T_2095_17; // @[NV_NVDLA_CSC_wl.scala 780:30:@17944.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_18 = _T_2095_18; // @[NV_NVDLA_CSC_wl.scala 780:30:@17945.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_19 = _T_2095_19; // @[NV_NVDLA_CSC_wl.scala 780:30:@17946.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_20 = _T_2095_20; // @[NV_NVDLA_CSC_wl.scala 780:30:@17947.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_21 = _T_2095_21; // @[NV_NVDLA_CSC_wl.scala 780:30:@17948.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_22 = _T_2095_22; // @[NV_NVDLA_CSC_wl.scala 780:30:@17949.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_23 = _T_2095_23; // @[NV_NVDLA_CSC_wl.scala 780:30:@17950.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_24 = _T_2095_24; // @[NV_NVDLA_CSC_wl.scala 780:30:@17951.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_25 = _T_2095_25; // @[NV_NVDLA_CSC_wl.scala 780:30:@17952.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_26 = _T_2095_26; // @[NV_NVDLA_CSC_wl.scala 780:30:@17953.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_27 = _T_2095_27; // @[NV_NVDLA_CSC_wl.scala 780:30:@17954.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_28 = _T_2095_28; // @[NV_NVDLA_CSC_wl.scala 780:30:@17955.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_29 = _T_2095_29; // @[NV_NVDLA_CSC_wl.scala 780:30:@17956.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_30 = _T_2095_30; // @[NV_NVDLA_CSC_wl.scala 780:30:@17957.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_31 = _T_2095_31; // @[NV_NVDLA_CSC_wl.scala 780:30:@17958.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_32 = _T_2095_32; // @[NV_NVDLA_CSC_wl.scala 780:30:@17959.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_33 = _T_2095_33; // @[NV_NVDLA_CSC_wl.scala 780:30:@17960.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_34 = _T_2095_34; // @[NV_NVDLA_CSC_wl.scala 780:30:@17961.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_35 = _T_2095_35; // @[NV_NVDLA_CSC_wl.scala 780:30:@17962.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_36 = _T_2095_36; // @[NV_NVDLA_CSC_wl.scala 780:30:@17963.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_37 = _T_2095_37; // @[NV_NVDLA_CSC_wl.scala 780:30:@17964.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_38 = _T_2095_38; // @[NV_NVDLA_CSC_wl.scala 780:30:@17965.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_39 = _T_2095_39; // @[NV_NVDLA_CSC_wl.scala 780:30:@17966.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_40 = _T_2095_40; // @[NV_NVDLA_CSC_wl.scala 780:30:@17967.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_41 = _T_2095_41; // @[NV_NVDLA_CSC_wl.scala 780:30:@17968.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_42 = _T_2095_42; // @[NV_NVDLA_CSC_wl.scala 780:30:@17969.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_43 = _T_2095_43; // @[NV_NVDLA_CSC_wl.scala 780:30:@17970.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_44 = _T_2095_44; // @[NV_NVDLA_CSC_wl.scala 780:30:@17971.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_45 = _T_2095_45; // @[NV_NVDLA_CSC_wl.scala 780:30:@17972.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_46 = _T_2095_46; // @[NV_NVDLA_CSC_wl.scala 780:30:@17973.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_47 = _T_2095_47; // @[NV_NVDLA_CSC_wl.scala 780:30:@17974.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_48 = _T_2095_48; // @[NV_NVDLA_CSC_wl.scala 780:30:@17975.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_49 = _T_2095_49; // @[NV_NVDLA_CSC_wl.scala 780:30:@17976.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_50 = _T_2095_50; // @[NV_NVDLA_CSC_wl.scala 780:30:@17977.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_51 = _T_2095_51; // @[NV_NVDLA_CSC_wl.scala 780:30:@17978.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_52 = _T_2095_52; // @[NV_NVDLA_CSC_wl.scala 780:30:@17979.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_53 = _T_2095_53; // @[NV_NVDLA_CSC_wl.scala 780:30:@17980.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_54 = _T_2095_54; // @[NV_NVDLA_CSC_wl.scala 780:30:@17981.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_55 = _T_2095_55; // @[NV_NVDLA_CSC_wl.scala 780:30:@17982.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_56 = _T_2095_56; // @[NV_NVDLA_CSC_wl.scala 780:30:@17983.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_57 = _T_2095_57; // @[NV_NVDLA_CSC_wl.scala 780:30:@17984.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_58 = _T_2095_58; // @[NV_NVDLA_CSC_wl.scala 780:30:@17985.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_59 = _T_2095_59; // @[NV_NVDLA_CSC_wl.scala 780:30:@17986.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_60 = _T_2095_60; // @[NV_NVDLA_CSC_wl.scala 780:30:@17987.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_61 = _T_2095_61; // @[NV_NVDLA_CSC_wl.scala 780:30:@17988.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_62 = _T_2095_62; // @[NV_NVDLA_CSC_wl.scala 780:30:@17989.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_63 = _T_2095_63; // @[NV_NVDLA_CSC_wl.scala 780:30:@17990.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_0 = _T_2362[0]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18057.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_1 = _T_2362[1]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18058.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_2 = _T_2362[2]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18059.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_3 = _T_2362[3]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18060.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_4 = _T_2362[4]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18061.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_5 = _T_2362[5]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18062.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_6 = _T_2362[6]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18063.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_7 = _T_2362[7]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18064.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_8 = _T_2362[8]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18065.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_9 = _T_2362[9]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18066.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_10 = _T_2362[10]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18067.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_11 = _T_2362[11]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18068.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_12 = _T_2362[12]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18069.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_13 = _T_2362[13]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18070.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_14 = _T_2362[14]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18071.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_15 = _T_2362[15]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18072.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_16 = _T_2362[16]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18073.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_17 = _T_2362[17]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18074.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_18 = _T_2362[18]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18075.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_19 = _T_2362[19]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18076.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_20 = _T_2362[20]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18077.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_21 = _T_2362[21]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18078.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_22 = _T_2362[22]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18079.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_23 = _T_2362[23]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18080.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_24 = _T_2362[24]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18081.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_25 = _T_2362[25]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18082.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_26 = _T_2362[26]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18083.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_27 = _T_2362[27]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18084.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_28 = _T_2362[28]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18085.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_29 = _T_2362[29]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18086.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_30 = _T_2362[30]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18087.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_31 = _T_2362[31]; // @[NV_NVDLA_CSC_wl.scala 784:29:@18088.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_mask_en = _T_2938; // @[NV_NVDLA_CSC_wl.scala 782:28:@18055.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_698 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_715 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_722 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_729 = _RAND_3[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_736 = _RAND_4[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_739 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_742 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1692 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{`RANDOM}};
  _T_1712 = _RAND_8[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_798 = _RAND_9[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_863 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_867 = _RAND_11[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_871 = _RAND_12[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_877 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_882 = _RAND_14[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_893 = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_896 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_920 = _RAND_17[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_923 = _RAND_18[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_1003 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_1006 = _RAND_20[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_1041 = _RAND_21[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_1044 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_1047 = _RAND_23[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_1050 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_1053 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_1056 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_1059 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_1062 = _RAND_28[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_1081 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_1084 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_1087 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_1090 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_1093 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_1096 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_1101 = _RAND_35[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_1104 = _RAND_36[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_1107 = _RAND_37[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_1110 = _RAND_38[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_1113 = _RAND_39[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_1116 = _RAND_40[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {10{`RANDOM}};
  _T_1156 = _RAND_41[318:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {16{`RANDOM}};
  _T_1163 = _RAND_42[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {16{`RANDOM}};
  _T_1193 = _RAND_43[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_1223 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_1226 = _RAND_45[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_1229 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_1232 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_1235 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_1238 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_1241 = _RAND_50[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_1244 = _RAND_51[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_1247 = _RAND_52[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {2{`RANDOM}};
  _T_1447 = _RAND_53[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_1537 = _RAND_54[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_1540 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_1563 = _RAND_56[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_1566 = _RAND_57[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_1605 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_1608 = _RAND_59[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_1631 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_1634 = _RAND_61[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_1637 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_1640 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_1643 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_1646 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_1649 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_1652 = _RAND_67[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_1655 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_1658 = _RAND_69[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_1661 = _RAND_70[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_1677 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_1680 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_1683 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_1686 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_1689 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {2{`RANDOM}};
  _T_1697 = _RAND_76[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {2{`RANDOM}};
  _T_1700 = _RAND_77[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {2{`RANDOM}};
  _T_1703 = _RAND_78[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {2{`RANDOM}};
  _T_1706 = _RAND_79[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {2{`RANDOM}};
  _T_1709 = _RAND_80[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_1717 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_1720 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_1723 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_1726 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_1729 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_1732 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {2{`RANDOM}};
  _T_1737 = _RAND_87[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {2{`RANDOM}};
  _T_1740 = _RAND_88[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {2{`RANDOM}};
  _T_1743 = _RAND_89[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {2{`RANDOM}};
  _T_1746 = _RAND_90[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {2{`RANDOM}};
  _T_1749 = _RAND_91[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {2{`RANDOM}};
  _T_1752 = _RAND_92[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_1762 = _RAND_93[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_1765 = _RAND_94[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {16{`RANDOM}};
  _T_1786 = _RAND_95[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {16{`RANDOM}};
  _T_1788 = _RAND_96[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_2095_0 = _RAND_97[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_2095_1 = _RAND_98[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_2095_2 = _RAND_99[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_2095_3 = _RAND_100[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_2095_4 = _RAND_101[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_2095_5 = _RAND_102[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_2095_6 = _RAND_103[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_2095_7 = _RAND_104[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_2095_8 = _RAND_105[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_2095_9 = _RAND_106[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_2095_10 = _RAND_107[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_2095_11 = _RAND_108[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_2095_12 = _RAND_109[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_2095_13 = _RAND_110[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_2095_14 = _RAND_111[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_2095_15 = _RAND_112[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_2095_16 = _RAND_113[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_2095_17 = _RAND_114[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_2095_18 = _RAND_115[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_2095_19 = _RAND_116[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_2095_20 = _RAND_117[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_2095_21 = _RAND_118[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_2095_22 = _RAND_119[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_2095_23 = _RAND_120[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_2095_24 = _RAND_121[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_2095_25 = _RAND_122[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_2095_26 = _RAND_123[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_2095_27 = _RAND_124[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_2095_28 = _RAND_125[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_2095_29 = _RAND_126[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_2095_30 = _RAND_127[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_2095_31 = _RAND_128[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_2095_32 = _RAND_129[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_2095_33 = _RAND_130[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_2095_34 = _RAND_131[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_2095_35 = _RAND_132[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_2095_36 = _RAND_133[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_2095_37 = _RAND_134[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_2095_38 = _RAND_135[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_2095_39 = _RAND_136[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_2095_40 = _RAND_137[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_2095_41 = _RAND_138[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_2095_42 = _RAND_139[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_2095_43 = _RAND_140[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_2095_44 = _RAND_141[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_2095_45 = _RAND_142[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_2095_46 = _RAND_143[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_2095_47 = _RAND_144[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_2095_48 = _RAND_145[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_2095_49 = _RAND_146[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_2095_50 = _RAND_147[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_2095_51 = _RAND_148[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_2095_52 = _RAND_149[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_2095_53 = _RAND_150[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_2095_54 = _RAND_151[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_2095_55 = _RAND_152[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_2095_56 = _RAND_153[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_2095_57 = _RAND_154[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_2095_58 = _RAND_155[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_2095_59 = _RAND_156[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_2095_60 = _RAND_157[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_2095_61 = _RAND_158[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_2095_62 = _RAND_159[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_2095_63 = _RAND_160[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_2359 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_2362 = _RAND_162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_2472 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_2739_0 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_2739_1 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_2739_2 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_2739_3 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_2739_4 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_2739_5 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_2739_6 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_2739_7 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_2739_8 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_2739_9 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_2739_10 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_2739_11 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_2739_12 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_2739_13 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_2739_14 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_2739_15 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_2739_16 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_2739_17 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_2739_18 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_2739_19 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_2739_20 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_2739_21 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_2739_22 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_2739_23 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_2739_24 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_2739_25 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_2739_26 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_2739_27 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_2739_28 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_2739_29 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_2739_30 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_2739_31 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_2739_32 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_2739_33 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_2739_34 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_2739_35 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_2739_36 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_2739_37 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_2739_38 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_2739_39 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_2739_40 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_2739_41 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_2739_42 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_2739_43 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_2739_44 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_2739_45 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_2739_46 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_2739_47 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_2739_48 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_2739_49 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_2739_50 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_2739_51 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_2739_52 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_2739_53 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_2739_54 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_2739_55 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_2739_56 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_2739_57 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_2739_58 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_2739_59 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_2739_60 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_2739_61 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_2739_62 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_2739_63 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_2938 = _RAND_228[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_3157 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_3160 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_3427_0 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_3427_1 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_3427_2 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_3427_3 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_3427_4 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_3427_5 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_3427_6 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_3427_7 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_3427_8 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_3427_9 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_3427_10 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_3427_11 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_3427_12 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_3427_13 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_3427_14 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_3427_15 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_3427_16 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_3427_17 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_3427_18 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_3427_19 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_3427_20 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_3427_21 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_3427_22 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_3427_23 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_3427_24 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_3427_25 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_3427_26 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_3427_27 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_3427_28 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_3427_29 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_3427_30 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_3427_31 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_3427_32 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_3427_33 = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_3427_34 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_3427_35 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_3427_36 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_3427_37 = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_3427_38 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_3427_39 = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_3427_40 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_3427_41 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_3427_42 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_3427_43 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_3427_44 = _RAND_275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_3427_45 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_3427_46 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_3427_47 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_3427_48 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_3427_49 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_3427_50 = _RAND_281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_3427_51 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_3427_52 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_3427_53 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_3427_54 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_3427_55 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_3427_56 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_3427_57 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_3427_58 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_3427_59 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_3427_60 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_3427_61 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_3427_62 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_3427_63 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_3890_0 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_3890_1 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_3890_2 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_3890_3 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_3890_4 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_3890_5 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_3890_6 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_3890_7 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_3890_8 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_3890_9 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_3890_10 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_3890_11 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_3890_12 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_3890_13 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_3890_14 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_3890_15 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_3890_16 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_3890_17 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_3890_18 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_3890_19 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_3890_20 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_3890_21 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_3890_22 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_3890_23 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_3890_24 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_3890_25 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_3890_26 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_3890_27 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_3890_28 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_3890_29 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_3890_30 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_3890_31 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_3890_32 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_3890_33 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_3890_34 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_3890_35 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_3890_36 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_3890_37 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_3890_38 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_3890_39 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_3890_40 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_3890_41 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_3890_42 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_3890_43 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_3890_44 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_3890_45 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_3890_46 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_3890_47 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_3890_48 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_3890_49 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_3890_50 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_3890_51 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_3890_52 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_3890_53 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_3890_54 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_3890_55 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_3890_56 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_3890_57 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_3890_58 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_3890_59 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_3890_60 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_3890_61 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_3890_62 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_3890_63 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_4161_0 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_4161_1 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_4161_2 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_4161_3 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_4161_4 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_4161_5 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_4161_6 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_4161_7 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_4161_8 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_4161_9 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_4161_10 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_4161_11 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_4161_12 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_4161_13 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_4161_14 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_4161_15 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_4288_0 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_4288_1 = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_4288_2 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_4288_3 = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_4288_4 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_4288_5 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_4288_6 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_4288_7 = _RAND_382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_4288_8 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_4288_9 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_4288_10 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_4288_11 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_4288_12 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_4288_13 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_4288_14 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_4288_15 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_4344_0 = _RAND_391[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_4344_1 = _RAND_392[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_4344_2 = _RAND_393[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_4344_3 = _RAND_394[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_4344_4 = _RAND_395[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_4344_5 = _RAND_396[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_4344_6 = _RAND_397[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_4344_7 = _RAND_398[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_4344_8 = _RAND_399[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_4344_9 = _RAND_400[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_4344_10 = _RAND_401[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_4344_11 = _RAND_402[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_4344_12 = _RAND_403[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_4344_13 = _RAND_404[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_4344_14 = _RAND_405[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_4344_15 = _RAND_406[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_4344_16 = _RAND_407[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_4344_17 = _RAND_408[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_4344_18 = _RAND_409[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_4344_19 = _RAND_410[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_4344_20 = _RAND_411[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_4344_21 = _RAND_412[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_4344_22 = _RAND_413[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_4344_23 = _RAND_414[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_4344_24 = _RAND_415[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_4344_25 = _RAND_416[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_4344_26 = _RAND_417[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_4344_27 = _RAND_418[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_4344_28 = _RAND_419[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_4344_29 = _RAND_420[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_4344_30 = _RAND_421[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_4344_31 = _RAND_422[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_4344_32 = _RAND_423[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_4344_33 = _RAND_424[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_4344_34 = _RAND_425[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_4344_35 = _RAND_426[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_4344_36 = _RAND_427[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_4344_37 = _RAND_428[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_4344_38 = _RAND_429[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_4344_39 = _RAND_430[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_4344_40 = _RAND_431[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_4344_41 = _RAND_432[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_4344_42 = _RAND_433[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_4344_43 = _RAND_434[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_4344_44 = _RAND_435[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_4344_45 = _RAND_436[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_4344_46 = _RAND_437[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_4344_47 = _RAND_438[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_4344_48 = _RAND_439[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_4344_49 = _RAND_440[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_4344_50 = _RAND_441[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_4344_51 = _RAND_442[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_4344_52 = _RAND_443[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_4344_53 = _RAND_444[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_4344_54 = _RAND_445[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_4344_55 = _RAND_446[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_4344_56 = _RAND_447[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_4344_57 = _RAND_448[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_4344_58 = _RAND_449[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_4344_59 = _RAND_450[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_4344_60 = _RAND_451[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_4344_61 = _RAND_452[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_4344_62 = _RAND_453[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_4344_63 = _RAND_454[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_4414_0 = _RAND_455[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_4414_1 = _RAND_456[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_4414_2 = _RAND_457[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_4414_3 = _RAND_458[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_4414_4 = _RAND_459[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_4414_5 = _RAND_460[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_4414_6 = _RAND_461[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_4414_7 = _RAND_462[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_4414_8 = _RAND_463[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_4414_9 = _RAND_464[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_4414_10 = _RAND_465[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_4414_11 = _RAND_466[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_4414_12 = _RAND_467[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_4414_13 = _RAND_468[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_4414_14 = _RAND_469[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_4414_15 = _RAND_470[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_4414_16 = _RAND_471[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_4414_17 = _RAND_472[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_4414_18 = _RAND_473[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_4414_19 = _RAND_474[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_4414_20 = _RAND_475[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_4414_21 = _RAND_476[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_4414_22 = _RAND_477[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_4414_23 = _RAND_478[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_4414_24 = _RAND_479[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_4414_25 = _RAND_480[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_4414_26 = _RAND_481[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_4414_27 = _RAND_482[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_4414_28 = _RAND_483[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_4414_29 = _RAND_484[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_4414_30 = _RAND_485[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_4414_31 = _RAND_486[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_4414_32 = _RAND_487[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_4414_33 = _RAND_488[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_4414_34 = _RAND_489[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_4414_35 = _RAND_490[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_4414_36 = _RAND_491[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_4414_37 = _RAND_492[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_4414_38 = _RAND_493[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_4414_39 = _RAND_494[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_4414_40 = _RAND_495[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_4414_41 = _RAND_496[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_4414_42 = _RAND_497[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_4414_43 = _RAND_498[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_4414_44 = _RAND_499[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_4414_45 = _RAND_500[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_4414_46 = _RAND_501[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_4414_47 = _RAND_502[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_4414_48 = _RAND_503[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_4414_49 = _RAND_504[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_4414_50 = _RAND_505[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_4414_51 = _RAND_506[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_4414_52 = _RAND_507[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_4414_53 = _RAND_508[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_4414_54 = _RAND_509[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_4414_55 = _RAND_510[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_4414_56 = _RAND_511[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_4414_57 = _RAND_512[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_4414_58 = _RAND_513[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_4414_59 = _RAND_514[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_4414_60 = _RAND_515[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_4414_61 = _RAND_516[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_4414_62 = _RAND_517[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_4414_63 = _RAND_518[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_698 <= 1'h0;
    end else begin
      _T_698 <= _T_704;
    end
    if (reset) begin
      _T_715 <= 5'h0;
    end else begin
      if (_T_743) begin
        _T_715 <= _T_750;
      end
    end
    if (reset) begin
      _T_722 <= 5'h0;
    end else begin
      if (_T_743) begin
        _T_722 <= _T_753;
      end
    end
    if (reset) begin
      _T_729 <= 15'h0;
    end else begin
      if (_T_757) begin
        _T_729 <= _T_758;
      end
    end
    if (reset) begin
      _T_736 <= 9'h0;
    end else begin
      if (_T_757) begin
        if (_T_742) begin
          _T_736 <= _T_759;
        end else begin
          _T_736 <= 9'h0;
        end
      end
    end
    if (reset) begin
      _T_739 <= 3'h1;
    end else begin
      if (_T_743) begin
        _T_739 <= _T_756;
      end
    end
    if (reset) begin
      _T_742 <= 1'h0;
    end else begin
      if (_T_743) begin
        _T_742 <= io_reg2dp_weight_format;
      end
    end
    if (reset) begin
      _T_1692 <= 1'h0;
    end else begin
      _T_1692 <= _T_1689;
    end
    if (reset) begin
      _T_1712 <= 36'h0;
    end else begin
      if (_T_1689) begin
        _T_1712 <= _T_1709;
      end
    end
    if (reset) begin
      _T_863 <= 1'h0;
    end else begin
      _T_863 <= _T_858;
    end
    if (reset) begin
      _T_867 <= 15'h0;
    end else begin
      if (_T_858) begin
        if (io_sg2wl_reuse_rls) begin
          _T_867 <= _T_729;
        end else begin
          _T_867 <= _T_1755;
        end
      end
    end
    if (reset) begin
      _T_871 <= 9'h0;
    end else begin
      if (_T_858) begin
        if (io_sg2wl_reuse_rls) begin
          _T_871 <= _T_736;
        end else begin
          _T_871 <= _T_1754;
        end
      end
    end
    if (reset) begin
      _T_877 <= 1'h0;
    end else begin
      _T_877 <= io_sg2wl_pd_valid;
    end
    if (reset) begin
      _T_882 <= 18'h0;
    end else begin
      if (io_sg2wl_pd_valid) begin
        _T_882 <= {{17'd0}, _T_879};
      end
    end
    if (reset) begin
      _T_893 <= 5'h0;
    end else begin
      if (_T_913) begin
        if (_T_743) begin
          _T_893 <= 5'h0;
        end else begin
          if (_T_905) begin
            _T_893 <= 5'h0;
          end else begin
            _T_893 <= _T_899;
          end
        end
      end
    end
    if (reset) begin
      _T_896 <= 1'h0;
    end else begin
      if (_T_877) begin
        _T_896 <= 1'h1;
      end else begin
        if (_T_909) begin
          _T_896 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_920 <= 11'h0;
    end else begin
      if (_T_972) begin
        if (_T_743) begin
          _T_920 <= 11'h0;
        end else begin
          if (_T_938) begin
            _T_920 <= _T_923;
          end else begin
            _T_920 <= _T_934;
          end
        end
      end
    end
    if (reset) begin
      _T_923 <= 11'h0;
    end else begin
      if (_T_976) begin
        if (_T_743) begin
          _T_923 <= 11'h0;
        end else begin
          if (!(_T_938)) begin
            _T_923 <= _T_934;
          end
        end
      end
    end
    if (reset) begin
      _T_1003 <= 1'h0;
    end else begin
      if (_T_1008) begin
        _T_1003 <= 1'h0;
      end else begin
        if (_T_1010) begin
          _T_1003 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_1006 <= 9'h0;
    end else begin
      if (_T_1029) begin
        if (_T_743) begin
          _T_1006 <= 9'h0;
        end else begin
          if (_T_1018) begin
            _T_1006 <= 9'h0;
          end else begin
            _T_1006 <= _T_1016;
          end
        end
      end
    end
    if (reset) begin
      _T_1041 <= 7'h0;
    end else begin
      if (_T_912) begin
        _T_1041 <= _T_883;
      end
    end
    if (reset) begin
      _T_1044 <= 8'h0;
    end else begin
      if (_T_912) begin
        _T_1044 <= _T_917;
      end
    end
    if (reset) begin
      _T_1047 <= 9'h0;
    end else begin
      if (_T_1064) begin
        if (_T_1031) begin
          _T_1047 <= _T_1006;
        end else begin
          _T_1047 <= _T_1016;
        end
      end
    end
    if (reset) begin
      _T_1050 <= 1'h0;
    end else begin
      if (_T_912) begin
        _T_1050 <= _T_905;
      end
    end
    if (reset) begin
      _T_1053 <= 1'h0;
    end else begin
      if (_T_912) begin
        _T_1053 <= _T_1010;
      end
    end
    if (reset) begin
      _T_1056 <= 1'h0;
    end else begin
      if (_T_912) begin
        _T_1056 <= _T_1007;
      end
    end
    if (reset) begin
      _T_1059 <= 1'h0;
    end else begin
      if (_T_912) begin
        _T_1059 <= _T_1067;
      end
    end
    if (reset) begin
      _T_1062 <= 2'h0;
    end else begin
      if (_T_912) begin
        _T_1062 <= _T_885;
      end
    end
    if (reset) begin
      _T_1081 <= 1'h0;
    end else begin
      _T_1081 <= _T_896;
    end
    if (reset) begin
      _T_1084 <= 1'h0;
    end else begin
      _T_1084 <= _T_1081;
    end
    if (reset) begin
      _T_1087 <= 1'h0;
    end else begin
      _T_1087 <= _T_1084;
    end
    if (reset) begin
      _T_1090 <= 1'h0;
    end else begin
      _T_1090 <= _T_1087;
    end
    if (reset) begin
      _T_1093 <= 1'h0;
    end else begin
      _T_1093 <= _T_1090;
    end
    if (reset) begin
      _T_1096 <= 1'h0;
    end else begin
      _T_1096 <= _T_1093;
    end
    if (reset) begin
      _T_1101 <= 31'h0;
    end else begin
      if (_T_896) begin
        _T_1101 <= _T_1076;
      end
    end
    if (reset) begin
      _T_1104 <= 31'h0;
    end else begin
      if (_T_1081) begin
        _T_1104 <= _T_1101;
      end
    end
    if (reset) begin
      _T_1107 <= 31'h0;
    end else begin
      if (_T_1084) begin
        _T_1107 <= _T_1104;
      end
    end
    if (reset) begin
      _T_1110 <= 31'h0;
    end else begin
      if (_T_1087) begin
        _T_1110 <= _T_1107;
      end
    end
    if (reset) begin
      _T_1113 <= 31'h0;
    end else begin
      if (_T_1090) begin
        _T_1113 <= _T_1110;
      end
    end
    if (reset) begin
      _T_1116 <= 31'h0;
    end else begin
      if (_T_1093) begin
        _T_1116 <= _T_1113;
      end
    end
    if (reset) begin
      _T_1156 <= 319'h0;
    end else begin
      if (_T_1096) begin
        _T_1156 <= _T_1186;
      end
    end
    if (reset) begin
      _T_1163 <= 512'h0;
    end else begin
      if (_T_1149) begin
        if (_T_743) begin
          _T_1163 <= 512'h0;
        end else begin
          if (_T_1138) begin
            _T_1163 <= _T_1193;
          end else begin
            _T_1163 <= _T_1199;
          end
        end
      end
    end
    if (reset) begin
      _T_1193 <= 512'h0;
    end else begin
      if (_T_1147) begin
        if (_T_743) begin
          _T_1193 <= 512'h0;
        end else begin
          if (!(_T_1138)) begin
            _T_1193 <= _T_1199;
          end
        end
      end
    end
    if (reset) begin
      _T_1223 <= 1'h0;
    end else begin
      _T_1223 <= _T_1096;
    end
    if (reset) begin
      _T_1226 <= 7'h0;
    end else begin
      if (_T_1096) begin
        _T_1226 <= _T_1117;
      end
    end
    if (reset) begin
      _T_1229 <= 1'h0;
    end else begin
      if (_T_1096) begin
        _T_1229 <= _T_1120;
      end
    end
    if (reset) begin
      _T_1232 <= 1'h0;
    end else begin
      if (_T_1096) begin
        _T_1232 <= _T_1121;
      end
    end
    if (reset) begin
      _T_1235 <= 1'h0;
    end else begin
      if (_T_1096) begin
        _T_1235 <= _T_1122;
      end
    end
    if (reset) begin
      _T_1238 <= 1'h0;
    end else begin
      if (_T_1096) begin
        _T_1238 <= _T_1123;
      end
    end
    if (reset) begin
      _T_1241 <= 9'h0;
    end else begin
      if (_T_1096) begin
        _T_1241 <= _T_1119;
      end
    end
    if (reset) begin
      _T_1244 <= 2'h0;
    end else begin
      if (_T_1096) begin
        _T_1244 <= _T_1124;
      end
    end
    if (reset) begin
      _T_1247 <= 7'h0;
    end else begin
      if (_T_1096) begin
        _T_1247 <= {{1'd0}, _T_1220};
      end
    end
    if (reset) begin
      _T_1447 <= 64'h0;
    end else begin
      _T_1447 <= _GEN_60[63:0];
    end
    if (reset) begin
      _T_1537 <= 8'h0;
    end else begin
      _T_1537 <= _GEN_49[7:0];
    end
    if (reset) begin
      _T_1540 <= 8'h0;
    end else begin
      _T_1540 <= _GEN_50[7:0];
    end
    if (reset) begin
      _T_1563 <= 13'h0;
    end else begin
      if (_T_1591) begin
        if (_T_708) begin
          _T_1563 <= _T_1583;
        end else begin
          if (_T_1554) begin
            _T_1563 <= _T_1566;
          end else begin
            if (_T_1542) begin
              if (_T_1576) begin
                _T_1563 <= 13'h0;
              end else begin
                _T_1563 <= _T_1569;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1566 <= 13'h0;
    end else begin
      if (_T_1594) begin
        if (_T_708) begin
          _T_1566 <= _T_1583;
        end else begin
          if (!(_T_1554)) begin
            if (_T_1542) begin
              if (_T_1576) begin
                _T_1566 <= 13'h0;
              end else begin
                _T_1566 <= _T_1569;
              end
            end else begin
              _T_1566 <= _T_1563;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1605 <= 1'h0;
    end else begin
      if (_T_1609) begin
        _T_1605 <= 1'h0;
      end else begin
        if (_T_1232) begin
          _T_1605 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_1608 <= 15'h0;
    end else begin
      if (_T_1625) begin
        if (_T_743) begin
          _T_1608 <= 15'h0;
        end else begin
          if (_T_1235) begin
            _T_1608 <= 15'h0;
          end else begin
            _T_1608 <= _T_1616;
          end
        end
      end
    end
    if (reset) begin
      _T_1631 <= 1'h0;
    end else begin
      _T_1631 <= _T_1542;
    end
    if (reset) begin
      _T_1634 <= 13'h0;
    end else begin
      _T_1634 <= _GEN_54[12:0];
    end
    if (reset) begin
      _T_1637 <= 1'h0;
    end else begin
      _T_1637 <= _T_1223;
    end
    if (reset) begin
      _T_1640 <= 1'h0;
    end else begin
      if (_T_1223) begin
        _T_1640 <= _T_1229;
      end
    end
    if (reset) begin
      _T_1643 <= 1'h0;
    end else begin
      if (_T_1223) begin
        _T_1643 <= _T_1232;
      end
    end
    if (reset) begin
      _T_1646 <= 1'h0;
    end else begin
      if (_T_1223) begin
        _T_1646 <= _T_1235;
      end
    end
    if (reset) begin
      _T_1649 <= 1'h0;
    end else begin
      if (_T_1223) begin
        _T_1649 <= _T_1238;
      end
    end
    if (reset) begin
      _T_1652 <= 8'h0;
    end else begin
      _T_1652 <= _GEN_59[7:0];
    end
    if (reset) begin
      _T_1655 <= 1'h0;
    end else begin
      _T_1655 <= _T_1534;
    end
    if (reset) begin
      _T_1658 <= 9'h0;
    end else begin
      if (_T_1223) begin
        _T_1658 <= _T_1241;
      end
    end
    if (reset) begin
      _T_1661 <= 15'h0;
    end else begin
      if (_T_1663) begin
        if (_T_1627) begin
          _T_1661 <= _T_1608;
        end else begin
          _T_1661 <= _T_1616;
        end
      end
    end
    if (reset) begin
      _T_1677 <= 1'h0;
    end else begin
      _T_1677 <= _T_1637;
    end
    if (reset) begin
      _T_1680 <= 1'h0;
    end else begin
      _T_1680 <= _T_1677;
    end
    if (reset) begin
      _T_1683 <= 1'h0;
    end else begin
      _T_1683 <= _T_1680;
    end
    if (reset) begin
      _T_1686 <= 1'h0;
    end else begin
      _T_1686 <= _T_1683;
    end
    if (reset) begin
      _T_1689 <= 1'h0;
    end else begin
      _T_1689 <= _T_1686;
    end
    if (reset) begin
      _T_1697 <= 36'h0;
    end else begin
      if (_T_1637) begin
        _T_1697 <= _T_1672;
      end
    end
    if (reset) begin
      _T_1700 <= 36'h0;
    end else begin
      if (_T_1677) begin
        _T_1700 <= _T_1697;
      end
    end
    if (reset) begin
      _T_1703 <= 36'h0;
    end else begin
      if (_T_1680) begin
        _T_1703 <= _T_1700;
      end
    end
    if (reset) begin
      _T_1706 <= 36'h0;
    end else begin
      if (_T_1683) begin
        _T_1706 <= _T_1703;
      end
    end
    if (reset) begin
      _T_1709 <= 36'h0;
    end else begin
      if (_T_1686) begin
        _T_1709 <= _T_1706;
      end
    end
    if (reset) begin
      _T_1717 <= 1'h0;
    end else begin
      _T_1717 <= _T_1655;
    end
    if (reset) begin
      _T_1720 <= 1'h0;
    end else begin
      _T_1720 <= _T_1717;
    end
    if (reset) begin
      _T_1723 <= 1'h0;
    end else begin
      _T_1723 <= _T_1720;
    end
    if (reset) begin
      _T_1726 <= 1'h0;
    end else begin
      _T_1726 <= _T_1723;
    end
    if (reset) begin
      _T_1729 <= 1'h0;
    end else begin
      _T_1729 <= _T_1726;
    end
    if (reset) begin
      _T_1732 <= 1'h0;
    end else begin
      _T_1732 <= _T_1729;
    end
    if (reset) begin
      _T_1737 <= 64'h0;
    end else begin
      if (_T_1655) begin
        _T_1737 <= _T_1447;
      end
    end
    if (reset) begin
      _T_1740 <= 64'h0;
    end else begin
      if (_T_1717) begin
        _T_1740 <= _T_1737;
      end
    end
    if (reset) begin
      _T_1743 <= 64'h0;
    end else begin
      if (_T_1720) begin
        _T_1743 <= _T_1740;
      end
    end
    if (reset) begin
      _T_1746 <= 64'h0;
    end else begin
      if (_T_1723) begin
        _T_1746 <= _T_1743;
      end
    end
    if (reset) begin
      _T_1749 <= 64'h0;
    end else begin
      if (_T_1726) begin
        _T_1749 <= _T_1746;
      end
    end
    if (reset) begin
      _T_1752 <= 64'h0;
    end else begin
      if (_T_1729) begin
        _T_1752 <= _T_1749;
      end
    end
    if (reset) begin
      _T_1762 <= 7'h0;
    end else begin
      if (_T_1782) begin
        _T_1762 <= _T_1781;
      end
    end
    if (reset) begin
      _T_1765 <= 7'h0;
    end else begin
      if (_T_1784) begin
        _T_1765 <= _T_1781;
      end
    end
    if (_T_1817) begin
      if (_T_743) begin
        _T_1786 <= 512'h0;
      end else begin
        if (_T_1810) begin
          _T_1786 <= _T_1788;
        end else begin
          if (io_sc2buf_wt_rd_data_valid) begin
            _T_1786 <= _T_1796;
          end else begin
            _T_1786 <= _T_1804;
          end
        end
      end
    end
    if (_T_1822) begin
      if (_T_743) begin
        _T_1788 <= 512'h0;
      end else begin
        if (!(_T_1810)) begin
          if (io_sc2buf_wt_rd_data_valid) begin
            _T_1788 <= _T_1796;
          end else begin
            _T_1788 <= _T_1804;
          end
        end
      end
    end
    if (reset) begin
      _T_2095_0 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_0 <= _T_2293;
      end
    end
    if (reset) begin
      _T_2095_1 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_1 <= _T_2294;
      end
    end
    if (reset) begin
      _T_2095_2 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_2 <= _T_2295;
      end
    end
    if (reset) begin
      _T_2095_3 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_3 <= _T_2296;
      end
    end
    if (reset) begin
      _T_2095_4 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_4 <= _T_2297;
      end
    end
    if (reset) begin
      _T_2095_5 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_5 <= _T_2298;
      end
    end
    if (reset) begin
      _T_2095_6 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_6 <= _T_2299;
      end
    end
    if (reset) begin
      _T_2095_7 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_7 <= _T_2300;
      end
    end
    if (reset) begin
      _T_2095_8 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_8 <= _T_2301;
      end
    end
    if (reset) begin
      _T_2095_9 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_9 <= _T_2302;
      end
    end
    if (reset) begin
      _T_2095_10 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_10 <= _T_2303;
      end
    end
    if (reset) begin
      _T_2095_11 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_11 <= _T_2304;
      end
    end
    if (reset) begin
      _T_2095_12 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_12 <= _T_2305;
      end
    end
    if (reset) begin
      _T_2095_13 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_13 <= _T_2306;
      end
    end
    if (reset) begin
      _T_2095_14 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_14 <= _T_2307;
      end
    end
    if (reset) begin
      _T_2095_15 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_15 <= _T_2308;
      end
    end
    if (reset) begin
      _T_2095_16 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_16 <= _T_2309;
      end
    end
    if (reset) begin
      _T_2095_17 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_17 <= _T_2310;
      end
    end
    if (reset) begin
      _T_2095_18 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_18 <= _T_2311;
      end
    end
    if (reset) begin
      _T_2095_19 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_19 <= _T_2312;
      end
    end
    if (reset) begin
      _T_2095_20 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_20 <= _T_2313;
      end
    end
    if (reset) begin
      _T_2095_21 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_21 <= _T_2314;
      end
    end
    if (reset) begin
      _T_2095_22 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_22 <= _T_2315;
      end
    end
    if (reset) begin
      _T_2095_23 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_23 <= _T_2316;
      end
    end
    if (reset) begin
      _T_2095_24 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_24 <= _T_2317;
      end
    end
    if (reset) begin
      _T_2095_25 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_25 <= _T_2318;
      end
    end
    if (reset) begin
      _T_2095_26 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_26 <= _T_2319;
      end
    end
    if (reset) begin
      _T_2095_27 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_27 <= _T_2320;
      end
    end
    if (reset) begin
      _T_2095_28 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_28 <= _T_2321;
      end
    end
    if (reset) begin
      _T_2095_29 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_29 <= _T_2322;
      end
    end
    if (reset) begin
      _T_2095_30 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_30 <= _T_2323;
      end
    end
    if (reset) begin
      _T_2095_31 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_31 <= _T_2324;
      end
    end
    if (reset) begin
      _T_2095_32 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_32 <= _T_2325;
      end
    end
    if (reset) begin
      _T_2095_33 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_33 <= _T_2326;
      end
    end
    if (reset) begin
      _T_2095_34 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_34 <= _T_2327;
      end
    end
    if (reset) begin
      _T_2095_35 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_35 <= _T_2328;
      end
    end
    if (reset) begin
      _T_2095_36 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_36 <= _T_2329;
      end
    end
    if (reset) begin
      _T_2095_37 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_37 <= _T_2330;
      end
    end
    if (reset) begin
      _T_2095_38 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_38 <= _T_2331;
      end
    end
    if (reset) begin
      _T_2095_39 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_39 <= _T_2332;
      end
    end
    if (reset) begin
      _T_2095_40 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_40 <= _T_2333;
      end
    end
    if (reset) begin
      _T_2095_41 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_41 <= _T_2334;
      end
    end
    if (reset) begin
      _T_2095_42 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_42 <= _T_2335;
      end
    end
    if (reset) begin
      _T_2095_43 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_43 <= _T_2336;
      end
    end
    if (reset) begin
      _T_2095_44 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_44 <= _T_2337;
      end
    end
    if (reset) begin
      _T_2095_45 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_45 <= _T_2338;
      end
    end
    if (reset) begin
      _T_2095_46 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_46 <= _T_2339;
      end
    end
    if (reset) begin
      _T_2095_47 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_47 <= _T_2340;
      end
    end
    if (reset) begin
      _T_2095_48 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_48 <= _T_2341;
      end
    end
    if (reset) begin
      _T_2095_49 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_49 <= _T_2342;
      end
    end
    if (reset) begin
      _T_2095_50 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_50 <= _T_2343;
      end
    end
    if (reset) begin
      _T_2095_51 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_51 <= _T_2344;
      end
    end
    if (reset) begin
      _T_2095_52 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_52 <= _T_2345;
      end
    end
    if (reset) begin
      _T_2095_53 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_53 <= _T_2346;
      end
    end
    if (reset) begin
      _T_2095_54 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_54 <= _T_2347;
      end
    end
    if (reset) begin
      _T_2095_55 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_55 <= _T_2348;
      end
    end
    if (reset) begin
      _T_2095_56 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_56 <= _T_2349;
      end
    end
    if (reset) begin
      _T_2095_57 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_57 <= _T_2350;
      end
    end
    if (reset) begin
      _T_2095_58 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_58 <= _T_2351;
      end
    end
    if (reset) begin
      _T_2095_59 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_59 <= _T_2352;
      end
    end
    if (reset) begin
      _T_2095_60 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_60 <= _T_2353;
      end
    end
    if (reset) begin
      _T_2095_61 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_61 <= _T_2354;
      end
    end
    if (reset) begin
      _T_2095_62 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_62 <= _T_2355;
      end
    end
    if (reset) begin
      _T_2095_63 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_63 <= _T_2356;
      end
    end
    if (reset) begin
      _T_2359 <= 1'h0;
    end else begin
      if (_T_1692) begin
        _T_2359 <= _T_1756;
      end
    end
    if (reset) begin
      _T_2362 <= 32'h1;
    end else begin
      if (_T_1692) begin
        if (_T_2359) begin
          _T_2362 <= 32'h1;
        end else begin
          _T_2362 <= _T_2366;
        end
      end
    end
    if (reset) begin
      _T_2472 <= 1'h0;
    end else begin
      _T_2472 <= _T_1692;
    end
    if (reset) begin
      _T_2739_0 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_0 <= _T_2939;
      end
    end
    if (reset) begin
      _T_2739_1 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_1 <= _T_2940;
      end
    end
    if (reset) begin
      _T_2739_2 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_2 <= _T_2941;
      end
    end
    if (reset) begin
      _T_2739_3 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_3 <= _T_2942;
      end
    end
    if (reset) begin
      _T_2739_4 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_4 <= _T_2943;
      end
    end
    if (reset) begin
      _T_2739_5 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_5 <= _T_2944;
      end
    end
    if (reset) begin
      _T_2739_6 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_6 <= _T_2945;
      end
    end
    if (reset) begin
      _T_2739_7 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_7 <= _T_2946;
      end
    end
    if (reset) begin
      _T_2739_8 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_8 <= _T_2947;
      end
    end
    if (reset) begin
      _T_2739_9 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_9 <= _T_2948;
      end
    end
    if (reset) begin
      _T_2739_10 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_10 <= _T_2949;
      end
    end
    if (reset) begin
      _T_2739_11 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_11 <= _T_2950;
      end
    end
    if (reset) begin
      _T_2739_12 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_12 <= _T_2951;
      end
    end
    if (reset) begin
      _T_2739_13 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_13 <= _T_2952;
      end
    end
    if (reset) begin
      _T_2739_14 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_14 <= _T_2953;
      end
    end
    if (reset) begin
      _T_2739_15 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_15 <= _T_2954;
      end
    end
    if (reset) begin
      _T_2739_16 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_16 <= _T_2955;
      end
    end
    if (reset) begin
      _T_2739_17 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_17 <= _T_2956;
      end
    end
    if (reset) begin
      _T_2739_18 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_18 <= _T_2957;
      end
    end
    if (reset) begin
      _T_2739_19 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_19 <= _T_2958;
      end
    end
    if (reset) begin
      _T_2739_20 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_20 <= _T_2959;
      end
    end
    if (reset) begin
      _T_2739_21 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_21 <= _T_2960;
      end
    end
    if (reset) begin
      _T_2739_22 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_22 <= _T_2961;
      end
    end
    if (reset) begin
      _T_2739_23 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_23 <= _T_2962;
      end
    end
    if (reset) begin
      _T_2739_24 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_24 <= _T_2963;
      end
    end
    if (reset) begin
      _T_2739_25 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_25 <= _T_2964;
      end
    end
    if (reset) begin
      _T_2739_26 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_26 <= _T_2965;
      end
    end
    if (reset) begin
      _T_2739_27 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_27 <= _T_2966;
      end
    end
    if (reset) begin
      _T_2739_28 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_28 <= _T_2967;
      end
    end
    if (reset) begin
      _T_2739_29 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_29 <= _T_2968;
      end
    end
    if (reset) begin
      _T_2739_30 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_30 <= _T_2969;
      end
    end
    if (reset) begin
      _T_2739_31 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_31 <= _T_2970;
      end
    end
    if (reset) begin
      _T_2739_32 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_32 <= _T_2971;
      end
    end
    if (reset) begin
      _T_2739_33 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_33 <= _T_2972;
      end
    end
    if (reset) begin
      _T_2739_34 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_34 <= _T_2973;
      end
    end
    if (reset) begin
      _T_2739_35 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_35 <= _T_2974;
      end
    end
    if (reset) begin
      _T_2739_36 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_36 <= _T_2975;
      end
    end
    if (reset) begin
      _T_2739_37 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_37 <= _T_2976;
      end
    end
    if (reset) begin
      _T_2739_38 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_38 <= _T_2977;
      end
    end
    if (reset) begin
      _T_2739_39 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_39 <= _T_2978;
      end
    end
    if (reset) begin
      _T_2739_40 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_40 <= _T_2979;
      end
    end
    if (reset) begin
      _T_2739_41 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_41 <= _T_2980;
      end
    end
    if (reset) begin
      _T_2739_42 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_42 <= _T_2981;
      end
    end
    if (reset) begin
      _T_2739_43 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_43 <= _T_2982;
      end
    end
    if (reset) begin
      _T_2739_44 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_44 <= _T_2983;
      end
    end
    if (reset) begin
      _T_2739_45 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_45 <= _T_2984;
      end
    end
    if (reset) begin
      _T_2739_46 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_46 <= _T_2985;
      end
    end
    if (reset) begin
      _T_2739_47 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_47 <= _T_2986;
      end
    end
    if (reset) begin
      _T_2739_48 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_48 <= _T_2987;
      end
    end
    if (reset) begin
      _T_2739_49 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_49 <= _T_2988;
      end
    end
    if (reset) begin
      _T_2739_50 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_50 <= _T_2989;
      end
    end
    if (reset) begin
      _T_2739_51 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_51 <= _T_2990;
      end
    end
    if (reset) begin
      _T_2739_52 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_52 <= _T_2991;
      end
    end
    if (reset) begin
      _T_2739_53 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_53 <= _T_2992;
      end
    end
    if (reset) begin
      _T_2739_54 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_54 <= _T_2993;
      end
    end
    if (reset) begin
      _T_2739_55 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_55 <= _T_2994;
      end
    end
    if (reset) begin
      _T_2739_56 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_56 <= _T_2995;
      end
    end
    if (reset) begin
      _T_2739_57 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_57 <= _T_2996;
      end
    end
    if (reset) begin
      _T_2739_58 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_58 <= _T_2997;
      end
    end
    if (reset) begin
      _T_2739_59 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_59 <= _T_2998;
      end
    end
    if (reset) begin
      _T_2739_60 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_60 <= _T_2999;
      end
    end
    if (reset) begin
      _T_2739_61 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_61 <= _T_3000;
      end
    end
    if (reset) begin
      _T_2739_62 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_62 <= _T_3001;
      end
    end
    if (reset) begin
      _T_2739_63 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_63 <= _T_3002;
      end
    end
    if (reset) begin
      _T_2938 <= 10'h0;
    end else begin
      if (_T_1732) begin
        _T_2938 <= 10'h3ff;
      end else begin
        _T_2938 <= 10'h0;
      end
    end
    if (reset) begin
      _T_3157 <= 1'h0;
    end else begin
      _T_3157 <= _T_3152;
    end
    if (reset) begin
      _T_3160 <= 1'h0;
    end else begin
      _T_3160 <= _T_3154;
    end
    if (reset) begin
      _T_3427_0 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_0 <= _T_4482;
      end
    end
    if (reset) begin
      _T_3427_1 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_1 <= _T_4484;
      end
    end
    if (reset) begin
      _T_3427_2 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_2 <= _T_4486;
      end
    end
    if (reset) begin
      _T_3427_3 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_3 <= _T_4488;
      end
    end
    if (reset) begin
      _T_3427_4 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_4 <= _T_4490;
      end
    end
    if (reset) begin
      _T_3427_5 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_5 <= _T_4492;
      end
    end
    if (reset) begin
      _T_3427_6 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_6 <= _T_4494;
      end
    end
    if (reset) begin
      _T_3427_7 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_7 <= _T_4496;
      end
    end
    if (reset) begin
      _T_3427_8 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_8 <= _T_4498;
      end
    end
    if (reset) begin
      _T_3427_9 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_9 <= _T_4500;
      end
    end
    if (reset) begin
      _T_3427_10 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_10 <= _T_4502;
      end
    end
    if (reset) begin
      _T_3427_11 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_11 <= _T_4504;
      end
    end
    if (reset) begin
      _T_3427_12 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_12 <= _T_4506;
      end
    end
    if (reset) begin
      _T_3427_13 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_13 <= _T_4508;
      end
    end
    if (reset) begin
      _T_3427_14 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_14 <= _T_4510;
      end
    end
    if (reset) begin
      _T_3427_15 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_15 <= _T_4512;
      end
    end
    if (reset) begin
      _T_3427_16 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_16 <= _T_4514;
      end
    end
    if (reset) begin
      _T_3427_17 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_17 <= _T_4516;
      end
    end
    if (reset) begin
      _T_3427_18 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_18 <= _T_4518;
      end
    end
    if (reset) begin
      _T_3427_19 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_19 <= _T_4520;
      end
    end
    if (reset) begin
      _T_3427_20 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_20 <= _T_4522;
      end
    end
    if (reset) begin
      _T_3427_21 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_21 <= _T_4524;
      end
    end
    if (reset) begin
      _T_3427_22 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_22 <= _T_4526;
      end
    end
    if (reset) begin
      _T_3427_23 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_23 <= _T_4528;
      end
    end
    if (reset) begin
      _T_3427_24 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_24 <= _T_4530;
      end
    end
    if (reset) begin
      _T_3427_25 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_25 <= _T_4532;
      end
    end
    if (reset) begin
      _T_3427_26 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_26 <= _T_4534;
      end
    end
    if (reset) begin
      _T_3427_27 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_27 <= _T_4536;
      end
    end
    if (reset) begin
      _T_3427_28 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_28 <= _T_4538;
      end
    end
    if (reset) begin
      _T_3427_29 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_29 <= _T_4540;
      end
    end
    if (reset) begin
      _T_3427_30 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_30 <= _T_4542;
      end
    end
    if (reset) begin
      _T_3427_31 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_31 <= _T_4544;
      end
    end
    if (reset) begin
      _T_3427_32 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_32 <= _T_4546;
      end
    end
    if (reset) begin
      _T_3427_33 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_33 <= _T_4548;
      end
    end
    if (reset) begin
      _T_3427_34 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_34 <= _T_4550;
      end
    end
    if (reset) begin
      _T_3427_35 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_35 <= _T_4552;
      end
    end
    if (reset) begin
      _T_3427_36 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_36 <= _T_4554;
      end
    end
    if (reset) begin
      _T_3427_37 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_37 <= _T_4556;
      end
    end
    if (reset) begin
      _T_3427_38 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_38 <= _T_4558;
      end
    end
    if (reset) begin
      _T_3427_39 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_39 <= _T_4560;
      end
    end
    if (reset) begin
      _T_3427_40 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_40 <= _T_4562;
      end
    end
    if (reset) begin
      _T_3427_41 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_41 <= _T_4564;
      end
    end
    if (reset) begin
      _T_3427_42 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_42 <= _T_4566;
      end
    end
    if (reset) begin
      _T_3427_43 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_43 <= _T_4568;
      end
    end
    if (reset) begin
      _T_3427_44 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_44 <= _T_4570;
      end
    end
    if (reset) begin
      _T_3427_45 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_45 <= _T_4572;
      end
    end
    if (reset) begin
      _T_3427_46 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_46 <= _T_4574;
      end
    end
    if (reset) begin
      _T_3427_47 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_47 <= _T_4576;
      end
    end
    if (reset) begin
      _T_3427_48 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_48 <= _T_4578;
      end
    end
    if (reset) begin
      _T_3427_49 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_49 <= _T_4580;
      end
    end
    if (reset) begin
      _T_3427_50 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_50 <= _T_4582;
      end
    end
    if (reset) begin
      _T_3427_51 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_51 <= _T_4584;
      end
    end
    if (reset) begin
      _T_3427_52 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_52 <= _T_4586;
      end
    end
    if (reset) begin
      _T_3427_53 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_53 <= _T_4588;
      end
    end
    if (reset) begin
      _T_3427_54 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_54 <= _T_4590;
      end
    end
    if (reset) begin
      _T_3427_55 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_55 <= _T_4592;
      end
    end
    if (reset) begin
      _T_3427_56 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_56 <= _T_4594;
      end
    end
    if (reset) begin
      _T_3427_57 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_57 <= _T_4596;
      end
    end
    if (reset) begin
      _T_3427_58 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_58 <= _T_4598;
      end
    end
    if (reset) begin
      _T_3427_59 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_59 <= _T_4600;
      end
    end
    if (reset) begin
      _T_3427_60 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_60 <= _T_4602;
      end
    end
    if (reset) begin
      _T_3427_61 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_61 <= _T_4604;
      end
    end
    if (reset) begin
      _T_3427_62 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_62 <= _T_4606;
      end
    end
    if (reset) begin
      _T_3427_63 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_63 <= _T_4608;
      end
    end
    if (reset) begin
      _T_3890_0 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_0 <= _T_4680;
      end
    end
    if (reset) begin
      _T_3890_1 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_1 <= _T_4682;
      end
    end
    if (reset) begin
      _T_3890_2 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_2 <= _T_4684;
      end
    end
    if (reset) begin
      _T_3890_3 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_3 <= _T_4686;
      end
    end
    if (reset) begin
      _T_3890_4 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_4 <= _T_4688;
      end
    end
    if (reset) begin
      _T_3890_5 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_5 <= _T_4690;
      end
    end
    if (reset) begin
      _T_3890_6 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_6 <= _T_4692;
      end
    end
    if (reset) begin
      _T_3890_7 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_7 <= _T_4694;
      end
    end
    if (reset) begin
      _T_3890_8 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_8 <= _T_4696;
      end
    end
    if (reset) begin
      _T_3890_9 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_9 <= _T_4698;
      end
    end
    if (reset) begin
      _T_3890_10 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_10 <= _T_4700;
      end
    end
    if (reset) begin
      _T_3890_11 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_11 <= _T_4702;
      end
    end
    if (reset) begin
      _T_3890_12 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_12 <= _T_4704;
      end
    end
    if (reset) begin
      _T_3890_13 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_13 <= _T_4706;
      end
    end
    if (reset) begin
      _T_3890_14 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_14 <= _T_4708;
      end
    end
    if (reset) begin
      _T_3890_15 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_15 <= _T_4710;
      end
    end
    if (reset) begin
      _T_3890_16 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_16 <= _T_4712;
      end
    end
    if (reset) begin
      _T_3890_17 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_17 <= _T_4714;
      end
    end
    if (reset) begin
      _T_3890_18 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_18 <= _T_4716;
      end
    end
    if (reset) begin
      _T_3890_19 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_19 <= _T_4718;
      end
    end
    if (reset) begin
      _T_3890_20 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_20 <= _T_4720;
      end
    end
    if (reset) begin
      _T_3890_21 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_21 <= _T_4722;
      end
    end
    if (reset) begin
      _T_3890_22 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_22 <= _T_4724;
      end
    end
    if (reset) begin
      _T_3890_23 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_23 <= _T_4726;
      end
    end
    if (reset) begin
      _T_3890_24 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_24 <= _T_4728;
      end
    end
    if (reset) begin
      _T_3890_25 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_25 <= _T_4730;
      end
    end
    if (reset) begin
      _T_3890_26 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_26 <= _T_4732;
      end
    end
    if (reset) begin
      _T_3890_27 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_27 <= _T_4734;
      end
    end
    if (reset) begin
      _T_3890_28 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_28 <= _T_4736;
      end
    end
    if (reset) begin
      _T_3890_29 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_29 <= _T_4738;
      end
    end
    if (reset) begin
      _T_3890_30 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_30 <= _T_4740;
      end
    end
    if (reset) begin
      _T_3890_31 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_31 <= _T_4742;
      end
    end
    if (reset) begin
      _T_3890_32 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_32 <= _T_4744;
      end
    end
    if (reset) begin
      _T_3890_33 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_33 <= _T_4746;
      end
    end
    if (reset) begin
      _T_3890_34 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_34 <= _T_4748;
      end
    end
    if (reset) begin
      _T_3890_35 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_35 <= _T_4750;
      end
    end
    if (reset) begin
      _T_3890_36 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_36 <= _T_4752;
      end
    end
    if (reset) begin
      _T_3890_37 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_37 <= _T_4754;
      end
    end
    if (reset) begin
      _T_3890_38 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_38 <= _T_4756;
      end
    end
    if (reset) begin
      _T_3890_39 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_39 <= _T_4758;
      end
    end
    if (reset) begin
      _T_3890_40 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_40 <= _T_4760;
      end
    end
    if (reset) begin
      _T_3890_41 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_41 <= _T_4762;
      end
    end
    if (reset) begin
      _T_3890_42 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_42 <= _T_4764;
      end
    end
    if (reset) begin
      _T_3890_43 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_43 <= _T_4766;
      end
    end
    if (reset) begin
      _T_3890_44 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_44 <= _T_4768;
      end
    end
    if (reset) begin
      _T_3890_45 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_45 <= _T_4770;
      end
    end
    if (reset) begin
      _T_3890_46 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_46 <= _T_4772;
      end
    end
    if (reset) begin
      _T_3890_47 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_47 <= _T_4774;
      end
    end
    if (reset) begin
      _T_3890_48 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_48 <= _T_4776;
      end
    end
    if (reset) begin
      _T_3890_49 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_49 <= _T_4778;
      end
    end
    if (reset) begin
      _T_3890_50 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_50 <= _T_4780;
      end
    end
    if (reset) begin
      _T_3890_51 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_51 <= _T_4782;
      end
    end
    if (reset) begin
      _T_3890_52 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_52 <= _T_4784;
      end
    end
    if (reset) begin
      _T_3890_53 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_53 <= _T_4786;
      end
    end
    if (reset) begin
      _T_3890_54 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_54 <= _T_4788;
      end
    end
    if (reset) begin
      _T_3890_55 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_55 <= _T_4790;
      end
    end
    if (reset) begin
      _T_3890_56 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_56 <= _T_4792;
      end
    end
    if (reset) begin
      _T_3890_57 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_57 <= _T_4794;
      end
    end
    if (reset) begin
      _T_3890_58 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_58 <= _T_4796;
      end
    end
    if (reset) begin
      _T_3890_59 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_59 <= _T_4798;
      end
    end
    if (reset) begin
      _T_3890_60 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_60 <= _T_4800;
      end
    end
    if (reset) begin
      _T_3890_61 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_61 <= _T_4802;
      end
    end
    if (reset) begin
      _T_3890_62 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_62 <= _T_4804;
      end
    end
    if (reset) begin
      _T_3890_63 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_63 <= _T_4806;
      end
    end
    if (reset) begin
      _T_4161_0 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_0 <= _T_4878;
      end
    end
    if (reset) begin
      _T_4161_1 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_1 <= _T_4879;
      end
    end
    if (reset) begin
      _T_4161_2 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_2 <= _T_4880;
      end
    end
    if (reset) begin
      _T_4161_3 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_3 <= _T_4881;
      end
    end
    if (reset) begin
      _T_4161_4 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_4 <= _T_4882;
      end
    end
    if (reset) begin
      _T_4161_5 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_5 <= _T_4883;
      end
    end
    if (reset) begin
      _T_4161_6 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_6 <= _T_4884;
      end
    end
    if (reset) begin
      _T_4161_7 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_7 <= _T_4885;
      end
    end
    if (reset) begin
      _T_4161_8 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_8 <= _T_4886;
      end
    end
    if (reset) begin
      _T_4161_9 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_9 <= _T_4887;
      end
    end
    if (reset) begin
      _T_4161_10 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_10 <= _T_4888;
      end
    end
    if (reset) begin
      _T_4161_11 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_11 <= _T_4889;
      end
    end
    if (reset) begin
      _T_4161_12 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_12 <= _T_4890;
      end
    end
    if (reset) begin
      _T_4161_13 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_13 <= _T_4891;
      end
    end
    if (reset) begin
      _T_4161_14 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_14 <= _T_4892;
      end
    end
    if (reset) begin
      _T_4161_15 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_15 <= _T_4893;
      end
    end
    if (reset) begin
      _T_4288_0 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_0 <= _T_4917;
      end
    end
    if (reset) begin
      _T_4288_1 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_1 <= _T_4918;
      end
    end
    if (reset) begin
      _T_4288_2 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_2 <= _T_4919;
      end
    end
    if (reset) begin
      _T_4288_3 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_3 <= _T_4920;
      end
    end
    if (reset) begin
      _T_4288_4 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_4 <= _T_4921;
      end
    end
    if (reset) begin
      _T_4288_5 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_5 <= _T_4922;
      end
    end
    if (reset) begin
      _T_4288_6 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_6 <= _T_4923;
      end
    end
    if (reset) begin
      _T_4288_7 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_7 <= _T_4924;
      end
    end
    if (reset) begin
      _T_4288_8 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_8 <= _T_4925;
      end
    end
    if (reset) begin
      _T_4288_9 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_9 <= _T_4926;
      end
    end
    if (reset) begin
      _T_4288_10 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_10 <= _T_4927;
      end
    end
    if (reset) begin
      _T_4288_11 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_11 <= _T_4928;
      end
    end
    if (reset) begin
      _T_4288_12 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_12 <= _T_4929;
      end
    end
    if (reset) begin
      _T_4288_13 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_13 <= _T_4930;
      end
    end
    if (reset) begin
      _T_4288_14 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_14 <= _T_4931;
      end
    end
    if (reset) begin
      _T_4288_15 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_15 <= _T_4932;
      end
    end
    if (_T_4482) begin
      _T_4344_0 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_0;
    end
    if (_T_4484) begin
      _T_4344_1 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_1;
    end
    if (_T_4486) begin
      _T_4344_2 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_2;
    end
    if (_T_4488) begin
      _T_4344_3 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_3;
    end
    if (_T_4490) begin
      _T_4344_4 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_4;
    end
    if (_T_4492) begin
      _T_4344_5 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_5;
    end
    if (_T_4494) begin
      _T_4344_6 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_6;
    end
    if (_T_4496) begin
      _T_4344_7 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_7;
    end
    if (_T_4498) begin
      _T_4344_8 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_8;
    end
    if (_T_4500) begin
      _T_4344_9 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_9;
    end
    if (_T_4502) begin
      _T_4344_10 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_10;
    end
    if (_T_4504) begin
      _T_4344_11 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_11;
    end
    if (_T_4506) begin
      _T_4344_12 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_12;
    end
    if (_T_4508) begin
      _T_4344_13 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_13;
    end
    if (_T_4510) begin
      _T_4344_14 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_14;
    end
    if (_T_4512) begin
      _T_4344_15 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_15;
    end
    if (_T_4514) begin
      _T_4344_16 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_16;
    end
    if (_T_4516) begin
      _T_4344_17 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_17;
    end
    if (_T_4518) begin
      _T_4344_18 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_18;
    end
    if (_T_4520) begin
      _T_4344_19 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_19;
    end
    if (_T_4522) begin
      _T_4344_20 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_20;
    end
    if (_T_4524) begin
      _T_4344_21 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_21;
    end
    if (_T_4526) begin
      _T_4344_22 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_22;
    end
    if (_T_4528) begin
      _T_4344_23 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_23;
    end
    if (_T_4530) begin
      _T_4344_24 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_24;
    end
    if (_T_4532) begin
      _T_4344_25 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_25;
    end
    if (_T_4534) begin
      _T_4344_26 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_26;
    end
    if (_T_4536) begin
      _T_4344_27 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_27;
    end
    if (_T_4538) begin
      _T_4344_28 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_28;
    end
    if (_T_4540) begin
      _T_4344_29 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_29;
    end
    if (_T_4542) begin
      _T_4344_30 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_30;
    end
    if (_T_4544) begin
      _T_4344_31 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_31;
    end
    if (_T_4546) begin
      _T_4344_32 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_32;
    end
    if (_T_4548) begin
      _T_4344_33 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_33;
    end
    if (_T_4550) begin
      _T_4344_34 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_34;
    end
    if (_T_4552) begin
      _T_4344_35 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_35;
    end
    if (_T_4554) begin
      _T_4344_36 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_36;
    end
    if (_T_4556) begin
      _T_4344_37 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_37;
    end
    if (_T_4558) begin
      _T_4344_38 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_38;
    end
    if (_T_4560) begin
      _T_4344_39 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_39;
    end
    if (_T_4562) begin
      _T_4344_40 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_40;
    end
    if (_T_4564) begin
      _T_4344_41 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_41;
    end
    if (_T_4566) begin
      _T_4344_42 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_42;
    end
    if (_T_4568) begin
      _T_4344_43 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_43;
    end
    if (_T_4570) begin
      _T_4344_44 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_44;
    end
    if (_T_4572) begin
      _T_4344_45 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_45;
    end
    if (_T_4574) begin
      _T_4344_46 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_46;
    end
    if (_T_4576) begin
      _T_4344_47 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_47;
    end
    if (_T_4578) begin
      _T_4344_48 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_48;
    end
    if (_T_4580) begin
      _T_4344_49 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_49;
    end
    if (_T_4582) begin
      _T_4344_50 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_50;
    end
    if (_T_4584) begin
      _T_4344_51 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_51;
    end
    if (_T_4586) begin
      _T_4344_52 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_52;
    end
    if (_T_4588) begin
      _T_4344_53 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_53;
    end
    if (_T_4590) begin
      _T_4344_54 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_54;
    end
    if (_T_4592) begin
      _T_4344_55 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_55;
    end
    if (_T_4594) begin
      _T_4344_56 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_56;
    end
    if (_T_4596) begin
      _T_4344_57 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_57;
    end
    if (_T_4598) begin
      _T_4344_58 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_58;
    end
    if (_T_4600) begin
      _T_4344_59 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_59;
    end
    if (_T_4602) begin
      _T_4344_60 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_60;
    end
    if (_T_4604) begin
      _T_4344_61 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_61;
    end
    if (_T_4606) begin
      _T_4344_62 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_62;
    end
    if (_T_4608) begin
      _T_4344_63 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_63;
    end
    if (_T_4680) begin
      _T_4414_0 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_0;
    end
    if (_T_4682) begin
      _T_4414_1 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_1;
    end
    if (_T_4684) begin
      _T_4414_2 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_2;
    end
    if (_T_4686) begin
      _T_4414_3 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_3;
    end
    if (_T_4688) begin
      _T_4414_4 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_4;
    end
    if (_T_4690) begin
      _T_4414_5 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_5;
    end
    if (_T_4692) begin
      _T_4414_6 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_6;
    end
    if (_T_4694) begin
      _T_4414_7 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_7;
    end
    if (_T_4696) begin
      _T_4414_8 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_8;
    end
    if (_T_4698) begin
      _T_4414_9 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_9;
    end
    if (_T_4700) begin
      _T_4414_10 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_10;
    end
    if (_T_4702) begin
      _T_4414_11 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_11;
    end
    if (_T_4704) begin
      _T_4414_12 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_12;
    end
    if (_T_4706) begin
      _T_4414_13 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_13;
    end
    if (_T_4708) begin
      _T_4414_14 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_14;
    end
    if (_T_4710) begin
      _T_4414_15 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_15;
    end
    if (_T_4712) begin
      _T_4414_16 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_16;
    end
    if (_T_4714) begin
      _T_4414_17 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_17;
    end
    if (_T_4716) begin
      _T_4414_18 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_18;
    end
    if (_T_4718) begin
      _T_4414_19 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_19;
    end
    if (_T_4720) begin
      _T_4414_20 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_20;
    end
    if (_T_4722) begin
      _T_4414_21 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_21;
    end
    if (_T_4724) begin
      _T_4414_22 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_22;
    end
    if (_T_4726) begin
      _T_4414_23 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_23;
    end
    if (_T_4728) begin
      _T_4414_24 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_24;
    end
    if (_T_4730) begin
      _T_4414_25 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_25;
    end
    if (_T_4732) begin
      _T_4414_26 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_26;
    end
    if (_T_4734) begin
      _T_4414_27 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_27;
    end
    if (_T_4736) begin
      _T_4414_28 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_28;
    end
    if (_T_4738) begin
      _T_4414_29 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_29;
    end
    if (_T_4740) begin
      _T_4414_30 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_30;
    end
    if (_T_4742) begin
      _T_4414_31 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_31;
    end
    if (_T_4744) begin
      _T_4414_32 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_32;
    end
    if (_T_4746) begin
      _T_4414_33 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_33;
    end
    if (_T_4748) begin
      _T_4414_34 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_34;
    end
    if (_T_4750) begin
      _T_4414_35 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_35;
    end
    if (_T_4752) begin
      _T_4414_36 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_36;
    end
    if (_T_4754) begin
      _T_4414_37 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_37;
    end
    if (_T_4756) begin
      _T_4414_38 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_38;
    end
    if (_T_4758) begin
      _T_4414_39 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_39;
    end
    if (_T_4760) begin
      _T_4414_40 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_40;
    end
    if (_T_4762) begin
      _T_4414_41 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_41;
    end
    if (_T_4764) begin
      _T_4414_42 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_42;
    end
    if (_T_4766) begin
      _T_4414_43 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_43;
    end
    if (_T_4768) begin
      _T_4414_44 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_44;
    end
    if (_T_4770) begin
      _T_4414_45 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_45;
    end
    if (_T_4772) begin
      _T_4414_46 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_46;
    end
    if (_T_4774) begin
      _T_4414_47 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_47;
    end
    if (_T_4776) begin
      _T_4414_48 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_48;
    end
    if (_T_4778) begin
      _T_4414_49 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_49;
    end
    if (_T_4780) begin
      _T_4414_50 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_50;
    end
    if (_T_4782) begin
      _T_4414_51 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_51;
    end
    if (_T_4784) begin
      _T_4414_52 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_52;
    end
    if (_T_4786) begin
      _T_4414_53 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_53;
    end
    if (_T_4788) begin
      _T_4414_54 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_54;
    end
    if (_T_4790) begin
      _T_4414_55 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_55;
    end
    if (_T_4792) begin
      _T_4414_56 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_56;
    end
    if (_T_4794) begin
      _T_4414_57 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_57;
    end
    if (_T_4796) begin
      _T_4414_58 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_58;
    end
    if (_T_4798) begin
      _T_4414_59 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_59;
    end
    if (_T_4800) begin
      _T_4414_60 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_60;
    end
    if (_T_4802) begin
      _T_4414_61 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_61;
    end
    if (_T_4804) begin
      _T_4414_62 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_62;
    end
    if (_T_4806) begin
      _T_4414_63 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_63;
    end
  end
  always @(posedge io_nvdla_core_ng_clk) begin
    if (reset) begin
      _T_798 <= 15'h0;
    end else begin
      if (_T_847) begin
        if (io_sc2cdma_wt_pending_req) begin
          _T_798 <= 15'h0;
        end else begin
          if (!(_T_810)) begin
            if (_T_808) begin
              _T_798 <= _T_805;
            end else begin
              _T_798 <= _T_800;
            end
          end
        end
      end
    end
  end
endmodule
module NV_NVDLA_CSC_dl( // @[:@19628.2]
  input          reset, // @[:@19630.4]
  input          io_nvdla_core_clk, // @[:@19631.4]
  input          io_nvdla_core_ng_clk, // @[:@19631.4]
  input  [1:0]   io_sc_state, // @[:@19631.4]
  input          io_sg2dl_pd_valid, // @[:@19631.4]
  input          io_sg2dl_reuse_rls, // @[:@19631.4]
  input          io_sc2cdma_dat_pending_req, // @[:@19631.4]
  output         io_sc2cdma_dat_updt_valid, // @[:@19631.4]
  output [14:0]  io_sc2cdma_dat_updt_bits_entries, // @[:@19631.4]
  output [13:0]  io_sc2cdma_dat_updt_bits_slices, // @[:@19631.4]
  output         io_sc2buf_dat_rd_addr_valid, // @[:@19631.4]
  output [12:0]  io_sc2buf_dat_rd_addr_bits, // @[:@19631.4]
  input          io_sc2buf_dat_rd_data_valid, // @[:@19631.4]
  input  [511:0] io_sc2buf_dat_rd_data_bits, // @[:@19631.4]
  output         io_sc2mac_dat_a_valid, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_0, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_1, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_2, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_3, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_4, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_5, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_6, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_7, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_8, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_9, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_10, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_11, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_12, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_13, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_14, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_15, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_16, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_17, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_18, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_19, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_20, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_21, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_22, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_23, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_24, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_25, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_26, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_27, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_28, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_29, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_30, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_31, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_32, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_33, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_34, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_35, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_36, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_37, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_38, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_39, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_40, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_41, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_42, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_43, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_44, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_45, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_46, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_47, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_48, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_49, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_50, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_51, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_52, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_53, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_54, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_55, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_56, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_57, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_58, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_59, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_60, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_61, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_62, // @[:@19631.4]
  output         io_sc2mac_dat_a_bits_mask_63, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_0, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_1, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_2, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_3, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_4, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_5, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_6, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_7, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_8, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_9, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_10, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_11, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_12, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_13, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_14, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_15, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_16, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_17, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_18, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_19, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_20, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_21, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_22, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_23, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_24, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_25, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_26, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_27, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_28, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_29, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_30, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_31, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_32, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_33, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_34, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_35, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_36, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_37, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_38, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_39, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_40, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_41, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_42, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_43, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_44, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_45, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_46, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_47, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_48, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_49, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_50, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_51, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_52, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_53, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_54, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_55, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_56, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_57, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_58, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_59, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_60, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_61, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_62, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_63, // @[:@19631.4]
  output [8:0]   io_sc2mac_dat_a_bits_pd, // @[:@19631.4]
  output         io_sc2mac_dat_b_valid, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_0, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_1, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_2, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_3, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_4, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_5, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_6, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_7, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_8, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_9, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_10, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_11, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_12, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_13, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_14, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_15, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_16, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_17, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_18, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_19, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_20, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_21, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_22, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_23, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_24, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_25, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_26, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_27, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_28, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_29, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_30, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_31, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_32, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_33, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_34, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_35, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_36, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_37, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_38, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_39, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_40, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_41, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_42, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_43, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_44, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_45, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_46, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_47, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_48, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_49, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_50, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_51, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_52, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_53, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_54, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_55, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_56, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_57, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_58, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_59, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_60, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_61, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_62, // @[:@19631.4]
  output         io_sc2mac_dat_b_bits_mask_63, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_0, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_1, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_2, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_3, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_4, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_5, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_6, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_7, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_8, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_9, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_10, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_11, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_12, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_13, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_14, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_15, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_16, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_17, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_18, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_19, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_20, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_21, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_22, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_23, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_24, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_25, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_26, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_27, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_28, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_29, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_30, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_31, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_32, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_33, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_34, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_35, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_36, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_37, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_38, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_39, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_40, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_41, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_42, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_43, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_44, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_45, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_46, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_47, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_48, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_49, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_50, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_51, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_52, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_53, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_54, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_55, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_56, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_57, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_58, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_59, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_60, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_61, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_62, // @[:@19631.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_63, // @[:@19631.4]
  output [8:0]   io_sc2mac_dat_b_bits_pd, // @[:@19631.4]
  input          io_reg2dp_op_en, // @[:@19631.4]
  input          io_reg2dp_conv_mode, // @[:@19631.4]
  input          io_reg2dp_datain_format, // @[:@19631.4]
  input          io_reg2dp_skip_data_rls, // @[:@19631.4]
  input  [12:0]  io_reg2dp_datain_channel_ext, // @[:@19631.4]
  input  [12:0]  io_reg2dp_datain_height_ext, // @[:@19631.4]
  input  [12:0]  io_reg2dp_datain_width_ext, // @[:@19631.4]
  input  [1:0]   io_reg2dp_y_extension, // @[:@19631.4]
  input  [12:0]  io_reg2dp_weight_channel_ext, // @[:@19631.4]
  input  [13:0]  io_reg2dp_entries, // @[:@19631.4]
  input  [12:0]  io_reg2dp_dataout_width, // @[:@19631.4]
  input  [11:0]  io_reg2dp_rls_slices, // @[:@19631.4]
  input  [2:0]   io_reg2dp_conv_x_stride_ext, // @[:@19631.4]
  input  [2:0]   io_reg2dp_conv_y_stride_ext, // @[:@19631.4]
  input  [4:0]   io_reg2dp_x_dilation_ext, // @[:@19631.4]
  input  [4:0]   io_reg2dp_y_dilation_ext, // @[:@19631.4]
  input  [4:0]   io_reg2dp_pad_left, // @[:@19631.4]
  input  [4:0]   io_reg2dp_pad_top, // @[:@19631.4]
  input  [15:0]  io_reg2dp_pad_value, // @[:@19631.4]
  input  [4:0]   io_reg2dp_data_bank // @[:@19631.4]
);
  wire  _T_622; // @[NV_NVDLA_CSC_dl.scala 75:31:@19633.4]
  wire  _T_626; // @[NV_NVDLA_CSC_dl.scala 77:31:@19635.4]
  wire  _T_630; // @[NV_NVDLA_CSC_dl.scala 84:32:@19638.4]
  wire  _T_634; // @[NV_NVDLA_CSC_dl.scala 86:35:@19640.4]
  wire  _T_635; // @[NV_NVDLA_CSC_dl.scala 87:22:@19641.4]
  wire [6:0] _T_640; // @[NV_NVDLA_CSC_dl.scala 94:53:@19642.4]
  wire [6:0] _T_642; // @[NV_NVDLA_CSC_dl.scala 94:24:@19643.4]
  wire [2:0] _T_643; // @[NV_NVDLA_CSC_dl.scala 94:100:@19644.4]
  wire [2:0] _T_645; // @[NV_NVDLA_CSC_dl.scala 95:22:@19645.4]
  wire [3:0] _T_647; // @[NV_NVDLA_CSC_dl.scala 96:34:@19646.4]
  wire [3:0] _T_648; // @[NV_NVDLA_CSC_dl.scala 96:34:@19647.4]
  wire [3:0] _T_650; // @[NV_NVDLA_CSC_dl.scala 97:51:@19648.4]
  wire [1:0] _T_651; // @[NV_NVDLA_CSC_dl.scala 98:62:@19649.4]
  wire [5:0] _T_654; // @[Cat.scala 30:58:@19650.4]
  wire [4:0] _T_657; // @[Cat.scala 30:58:@19651.4]
  wire [4:0] _GEN_671; // @[NV_NVDLA_CSC_dl.scala 100:74:@19652.4]
  wire [5:0] _T_658; // @[NV_NVDLA_CSC_dl.scala 100:74:@19652.4]
  wire  _T_659; // @[Mux.scala 46:19:@19653.4]
  wire [5:0] _T_660; // @[Mux.scala 46:16:@19654.4]
  wire  _T_661; // @[Mux.scala 46:19:@19655.4]
  wire [5:0] _T_662; // @[Mux.scala 46:16:@19656.4]
  wire  _T_664; // @[NV_NVDLA_CSC_dl.scala 102:88:@19657.4]
  wire [5:0] _T_670; // @[NV_NVDLA_CSC_dl.scala 102:172:@19659.4]
  wire [5:0] _T_671; // @[NV_NVDLA_CSC_dl.scala 102:58:@19660.4]
  wire [6:0] _T_674; // @[Cat.scala 30:58:@19661.4]
  wire [6:0] _GEN_672; // @[NV_NVDLA_CSC_dl.scala 103:81:@19662.4]
  wire [7:0] _T_675; // @[NV_NVDLA_CSC_dl.scala 103:81:@19662.4]
  wire [6:0] _T_676; // @[NV_NVDLA_CSC_dl.scala 103:81:@19663.4]
  wire [6:0] _GEN_673; // @[NV_NVDLA_CSC_dl.scala 103:100:@19665.4]
  wire [7:0] _T_678; // @[NV_NVDLA_CSC_dl.scala 103:100:@19665.4]
  wire [6:0] _T_679; // @[NV_NVDLA_CSC_dl.scala 103:100:@19666.4]
  wire [6:0] _T_682; // @[NV_NVDLA_CSC_dl.scala 104:58:@19668.4]
  wire [5:0] _T_683; // @[NV_NVDLA_CSC_dl.scala 104:58:@19669.4]
  wire  _T_684; // @[Mux.scala 46:19:@19670.4]
  wire [5:0] _T_685; // @[Mux.scala 46:16:@19671.4]
  wire  _T_686; // @[Mux.scala 46:19:@19672.4]
  wire [6:0] _T_687; // @[Mux.scala 46:16:@19673.4]
  wire [6:0] _T_690; // @[NV_NVDLA_CSC_dl.scala 105:80:@19675.4]
  wire [7:0] _T_693; // @[Cat.scala 30:58:@19676.4]
  wire [6:0] _T_698; // @[Mux.scala 46:16:@19679.4]
  wire [7:0] _T_700; // @[Mux.scala 46:16:@19681.4]
  wire [11:0] _T_702; // @[Cat.scala 30:58:@19682.4]
  wire [3:0] _T_704; // @[NV_NVDLA_CSC_dl.scala 115:52:@19683.4]
  wire [5:0] _T_707; // @[NV_NVDLA_CSC_dl.scala 116:60:@19684.4]
  wire [5:0] _T_708; // @[NV_NVDLA_CSC_dl.scala 116:21:@19685.4]
  wire [5:0] _T_711; // @[NV_NVDLA_CSC_dl.scala 117:60:@19686.4]
  wire [5:0] _T_712; // @[NV_NVDLA_CSC_dl.scala 117:21:@19687.4]
  reg  _T_715; // @[NV_NVDLA_CSC_dl.scala 119:26:@19688.4]
  reg [31:0] _RAND_0;
  reg [5:0] _T_722; // @[NV_NVDLA_CSC_dl.scala 120:25:@19690.4]
  reg [31:0] _RAND_1;
  reg [13:0] _T_729; // @[NV_NVDLA_CSC_dl.scala 121:25:@19692.4]
  reg [31:0] _RAND_2;
  reg [13:0] _T_736; // @[NV_NVDLA_CSC_dl.scala 122:29:@19694.4]
  reg [31:0] _RAND_3;
  reg [14:0] _T_743; // @[NV_NVDLA_CSC_dl.scala 123:22:@19696.4]
  reg [31:0] _RAND_4;
  reg [14:0] _T_750; // @[NV_NVDLA_CSC_dl.scala 124:28:@19698.4]
  reg [31:0] _RAND_5;
  reg [12:0] _T_757; // @[NV_NVDLA_CSC_dl.scala 125:32:@19700.4]
  reg [31:0] _RAND_6;
  reg [14:0] _T_771; // @[NV_NVDLA_CSC_dl.scala 127:26:@19704.4]
  reg [31:0] _RAND_7;
  reg [11:0] _T_778; // @[NV_NVDLA_CSC_dl.scala 128:30:@19706.4]
  reg [31:0] _RAND_8;
  reg [11:0] _T_785; // @[NV_NVDLA_CSC_dl.scala 129:30:@19708.4]
  reg [31:0] _RAND_9;
  reg [13:0] _T_792; // @[NV_NVDLA_CSC_dl.scala 130:25:@19710.4]
  reg [31:0] _RAND_10;
  wire [14:0] _T_794; // @[NV_NVDLA_CSC_dl.scala 133:43:@19711.4]
  wire [20:0] _T_796; // @[NV_NVDLA_CSC_dl.scala 134:41:@19713.4]
  wire [14:0] _T_797; // @[NV_NVDLA_CSC_dl.scala 134:56:@19714.4]
  wire [11:0] _T_798; // @[NV_NVDLA_CSC_dl.scala 136:37:@19715.4]
  wire [14:0] _GEN_674; // @[NV_NVDLA_CSC_dl.scala 137:34:@19716.4]
  wire [20:0] _T_799; // @[NV_NVDLA_CSC_dl.scala 137:34:@19716.4]
  wire [11:0] _T_800; // @[NV_NVDLA_CSC_dl.scala 137:47:@19717.4]
  wire [14:0] _GEN_675; // @[NV_NVDLA_CSC_dl.scala 138:34:@19718.4]
  wire [28:0] _T_801; // @[NV_NVDLA_CSC_dl.scala 138:34:@19718.4]
  wire [11:0] _T_802; // @[NV_NVDLA_CSC_dl.scala 138:51:@19719.4]
  wire [12:0] _T_804; // @[NV_NVDLA_CSC_dl.scala 139:41:@19720.4]
  wire [11:0] _T_805; // @[NV_NVDLA_CSC_dl.scala 139:41:@19721.4]
  wire [13:0] _T_807; // @[NV_NVDLA_CSC_dl.scala 140:77:@19722.4]
  wire [12:0] _GEN_676; // @[NV_NVDLA_CSC_dl.scala 140:113:@19723.4]
  wire [13:0] _T_808; // @[NV_NVDLA_CSC_dl.scala 140:113:@19723.4]
  wire [13:0] _T_809; // @[NV_NVDLA_CSC_dl.scala 140:113:@19724.4]
  wire [13:0] _T_810; // @[NV_NVDLA_CSC_dl.scala 140:23:@19725.4]
  wire [13:0] _T_811; // @[NV_NVDLA_CSC_dl.scala 141:24:@19726.4]
  wire [14:0] _GEN_677; // @[NV_NVDLA_CSC_dl.scala 142:38:@19727.4]
  wire [28:0] _T_812; // @[NV_NVDLA_CSC_dl.scala 142:38:@19727.4]
  wire [14:0] _T_813; // @[NV_NVDLA_CSC_dl.scala 142:54:@19728.4]
  reg [33:0] _T_831; // @[NV_NVDLA_CSC_dl.scala 147:24:@19734.4]
  reg [63:0] _RAND_11;
  reg [4:0] _T_838; // @[NV_NVDLA_CSC_dl.scala 148:24:@19736.4]
  reg [31:0] _RAND_12;
  reg [13:0] _T_845; // @[NV_NVDLA_CSC_dl.scala 149:27:@19738.4]
  reg [31:0] _RAND_13;
  reg [12:0] _T_852; // @[NV_NVDLA_CSC_dl.scala 150:31:@19740.4]
  reg [31:0] _RAND_14;
  reg [12:0] _T_859; // @[NV_NVDLA_CSC_dl.scala 151:32:@19742.4]
  reg [31:0] _RAND_15;
  reg [10:0] _T_866; // @[NV_NVDLA_CSC_dl.scala 152:33:@19744.4]
  reg [31:0] _RAND_16;
  reg [2:0] _T_869; // @[NV_NVDLA_CSC_dl.scala 153:29:@19745.4]
  reg [31:0] _RAND_17;
  reg [2:0] _T_872; // @[NV_NVDLA_CSC_dl.scala 154:29:@19746.4]
  reg [31:0] _RAND_18;
  reg [2:0] _T_878; // @[NV_NVDLA_CSC_dl.scala 156:29:@19748.4]
  reg [31:0] _RAND_19;
  reg [2:0] _T_881; // @[NV_NVDLA_CSC_dl.scala 157:29:@19749.4]
  reg [31:0] _RAND_20;
  reg [2:0] _T_884; // @[NV_NVDLA_CSC_dl.scala 158:29:@19750.4]
  reg [31:0] _RAND_21;
  reg [2:0] _T_887; // @[NV_NVDLA_CSC_dl.scala 159:29:@19751.4]
  reg [31:0] _RAND_22;
  reg [2:0] _T_893; // @[NV_NVDLA_CSC_dl.scala 161:29:@19753.4]
  reg [31:0] _RAND_23;
  reg [2:0] _T_896; // @[NV_NVDLA_CSC_dl.scala 162:29:@19754.4]
  reg [31:0] _RAND_24;
  reg [2:0] _T_902; // @[NV_NVDLA_CSC_dl.scala 164:30:@19756.4]
  reg [31:0] _RAND_25;
  reg [2:0] _T_905; // @[NV_NVDLA_CSC_dl.scala 165:27:@19757.4]
  reg [31:0] _RAND_26;
  reg [2:0] _T_908; // @[NV_NVDLA_CSC_dl.scala 166:27:@19758.4]
  reg [31:0] _RAND_27;
  reg [3:0] _T_915; // @[NV_NVDLA_CSC_dl.scala 167:28:@19760.4]
  reg [31:0] _RAND_28;
  reg [3:0] _T_922; // @[NV_NVDLA_CSC_dl.scala 168:28:@19762.4]
  reg [31:0] _RAND_29;
  reg [4:0] _T_932; // @[NV_NVDLA_CSC_dl.scala 170:24:@19765.4]
  reg [31:0] _RAND_30;
  reg [6:0] _T_939; // @[NV_NVDLA_CSC_dl.scala 171:27:@19767.4]
  reg [31:0] _RAND_31;
  reg [6:0] _T_946; // @[NV_NVDLA_CSC_dl.scala 172:34:@19769.4]
  reg [31:0] _RAND_32;
  reg [7:0] _T_953; // @[NV_NVDLA_CSC_dl.scala 173:26:@19771.4]
  reg [31:0] _RAND_33;
  reg [6:0] _T_960; // @[NV_NVDLA_CSC_dl.scala 174:34:@19773.4]
  reg [31:0] _RAND_34;
  reg [11:0] _T_967; // @[NV_NVDLA_CSC_dl.scala 175:30:@19775.4]
  reg [31:0] _RAND_35;
  reg [5:0] _T_974; // @[NV_NVDLA_CSC_dl.scala 176:23:@19777.4]
  reg [31:0] _RAND_36;
  reg [5:0] _T_981; // @[NV_NVDLA_CSC_dl.scala 177:23:@19779.4]
  reg [31:0] _RAND_37;
  reg [15:0] _T_988; // @[NV_NVDLA_CSC_dl.scala 178:24:@19781.4]
  reg [31:0] _RAND_38;
  reg [14:0] _T_995; // @[NV_NVDLA_CSC_dl.scala 179:26:@19783.4]
  reg [31:0] _RAND_39;
  reg [14:0] _T_1002; // @[NV_NVDLA_CSC_dl.scala 180:30:@19785.4]
  reg [31:0] _RAND_40;
  reg [14:0] _T_1009; // @[NV_NVDLA_CSC_dl.scala 181:30:@19787.4]
  reg [31:0] _RAND_41;
  reg [13:0] _T_1016; // @[NV_NVDLA_CSC_dl.scala 183:26:@19789.4]
  reg [31:0] _RAND_42;
  reg [14:0] _T_1023; // @[NV_NVDLA_CSC_dl.scala 184:27:@19791.4]
  reg [31:0] _RAND_43;
  wire [33:0] _T_1038; // @[Bitwise.scala 72:12:@19799.6]
  wire [5:0] _T_1040; // @[NV_NVDLA_CSC_dl.scala 191:38:@19801.6]
  wire [4:0] _T_1041; // @[NV_NVDLA_CSC_dl.scala 191:38:@19802.6]
  wire [13:0] _T_1043; // @[NV_NVDLA_CSC_dl.scala 192:48:@19804.6]
  wire [6:0] _T_1049; // @[NV_NVDLA_CSC_dl.scala 195:93:@19809.6]
  wire [10:0] _T_1050; // @[Cat.scala 30:58:@19810.6]
  wire [14:0] _T_1054; // @[Cat.scala 30:58:@19843.6]
  wire [33:0] _GEN_1; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [4:0] _GEN_2; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [13:0] _GEN_3; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [12:0] _GEN_4; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [12:0] _GEN_5; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [10:0] _GEN_6; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [2:0] _GEN_7; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [2:0] _GEN_8; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [2:0] _GEN_10; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [2:0] _GEN_11; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [2:0] _GEN_12; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [2:0] _GEN_13; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [2:0] _GEN_15; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [2:0] _GEN_16; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [2:0] _GEN_18; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [2:0] _GEN_19; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [2:0] _GEN_20; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [3:0] _GEN_21; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [3:0] _GEN_22; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [5:0] _GEN_24; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [4:0] _GEN_25; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [6:0] _GEN_26; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [6:0] _GEN_27; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [7:0] _GEN_28; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [6:0] _GEN_29; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [11:0] _GEN_30; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [5:0] _GEN_31; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [5:0] _GEN_32; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [15:0] _GEN_33; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [14:0] _GEN_34; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [14:0] _GEN_35; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [14:0] _GEN_36; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [13:0] _GEN_37; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [13:0] _GEN_38; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [13:0] _GEN_39; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [12:0] _GEN_40; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  wire [11:0] _GEN_43; // @[NV_NVDLA_CSC_dl.scala 233:18:@19856.4]
  wire [11:0] _GEN_44; // @[NV_NVDLA_CSC_dl.scala 233:18:@19856.4]
  wire [14:0] _GEN_45; // @[NV_NVDLA_CSC_dl.scala 233:18:@19856.4]
  wire [14:0] _GEN_46; // @[NV_NVDLA_CSC_dl.scala 233:18:@19856.4]
  wire [14:0] _GEN_47; // @[NV_NVDLA_CSC_dl.scala 233:18:@19856.4]
  wire [13:0] _GEN_48; // @[NV_NVDLA_CSC_dl.scala 240:17:@19863.4]
  wire [14:0] _GEN_49; // @[NV_NVDLA_CSC_dl.scala 240:17:@19863.4]
  reg [14:0] _T_1076; // @[NV_NVDLA_CSC_dl.scala 263:59:@19875.4]
  reg [31:0] _RAND_44;
  wire  _T_1156; // @[NV_NVDLA_CSC_dl.scala 304:37:@19938.4]
  wire  _T_1157; // @[NV_NVDLA_CSC_dl.scala 304:23:@19939.4]
  wire  _T_2241; // @[NV_NVDLA_CSC_dl.scala 894:32:@20853.4]
  reg  _T_2217; // @[NV_NVDLA_CSC_dl.scala 879:41:@20821.4]
  reg [31:0] _RAND_45;
  wire  _T_2242; // @[NV_NVDLA_CSC_dl.scala 894:36:@20854.4]
  wire  _T_2243; // @[NV_NVDLA_CSC_dl.scala 895:35:@20855.4]
  reg  _T_2211; // @[NV_NVDLA_CSC_dl.scala 879:41:@20819.4]
  reg [31:0] _RAND_46;
  wire  _T_2244; // @[NV_NVDLA_CSC_dl.scala 895:39:@20856.4]
  wire  _T_2245; // @[NV_NVDLA_CSC_dl.scala 894:57:@20857.4]
  wire  _T_2246; // @[NV_NVDLA_CSC_dl.scala 896:35:@20858.4]
  reg  _T_2208; // @[NV_NVDLA_CSC_dl.scala 879:41:@20818.4]
  reg [31:0] _RAND_47;
  wire  _T_2247; // @[NV_NVDLA_CSC_dl.scala 896:39:@20859.4]
  wire  _T_2248; // @[NV_NVDLA_CSC_dl.scala 895:60:@20860.4]
  wire  _T_2249; // @[NV_NVDLA_CSC_dl.scala 903:42:@20862.4]
  wire [26:0] _T_2253; // @[Bitwise.scala 72:12:@20864.4]
  reg [26:0] _T_2231; // @[NV_NVDLA_CSC_dl.scala 881:41:@20826.4]
  reg [31:0] _RAND_48;
  wire [26:0] _T_2254; // @[NV_NVDLA_CSC_dl.scala 903:47:@20865.4]
  wire  _T_2255; // @[NV_NVDLA_CSC_dl.scala 904:42:@20866.4]
  wire [26:0] _T_2259; // @[Bitwise.scala 72:12:@20868.4]
  reg [26:0] _T_2225; // @[NV_NVDLA_CSC_dl.scala 881:41:@20824.4]
  reg [31:0] _RAND_49;
  wire [26:0] _T_2260; // @[NV_NVDLA_CSC_dl.scala 904:47:@20869.4]
  wire [26:0] _T_2261; // @[NV_NVDLA_CSC_dl.scala 903:66:@20870.4]
  wire  _T_2262; // @[NV_NVDLA_CSC_dl.scala 905:42:@20871.4]
  wire [26:0] _T_2266; // @[Bitwise.scala 72:12:@20873.4]
  reg [26:0] _T_2222; // @[NV_NVDLA_CSC_dl.scala 881:41:@20823.4]
  reg [31:0] _RAND_50;
  wire [26:0] _T_2267; // @[NV_NVDLA_CSC_dl.scala 905:47:@20874.4]
  wire [26:0] _T_2268; // @[NV_NVDLA_CSC_dl.scala 904:66:@20875.4]
  wire  _T_2287; // @[NV_NVDLA_CSC_dl.scala 929:26:@20894.4]
  wire  _T_1154; // @[NV_NVDLA_CSC_dl.scala 301:29:@19937.4]
  wire  _T_1159; // @[NV_NVDLA_CSC_dl.scala 304:66:@19940.4]
  wire  _T_1160; // @[NV_NVDLA_CSC_dl.scala 304:53:@19941.4]
  wire  _T_1161; // @[NV_NVDLA_CSC_dl.scala 304:42:@19942.4]
  wire [13:0] _T_1162; // @[NV_NVDLA_CSC_dl.scala 305:28:@19944.4]
  wire [14:0] _T_1163; // @[NV_NVDLA_CSC_dl.scala 306:29:@19946.4]
  wire [14:0] _T_1094; // @[NV_NVDLA_CSC_dl.scala 273:28:@19886.4]
  wire [15:0] _T_1102; // @[NV_NVDLA_CSC_dl.scala 278:37:@19893.4]
  wire [14:0] _T_1103; // @[NV_NVDLA_CSC_dl.scala 278:37:@19894.4]
  wire [13:0] _T_1109; // @[Cat.scala 30:58:@19896.4]
  wire [14:0] _GEN_678; // @[NV_NVDLA_CSC_dl.scala 279:46:@19897.4]
  wire [15:0] _T_1110; // @[NV_NVDLA_CSC_dl.scala 279:46:@19897.4]
  wire [15:0] _T_1111; // @[NV_NVDLA_CSC_dl.scala 279:46:@19898.4]
  wire [14:0] _T_1112; // @[NV_NVDLA_CSC_dl.scala 279:46:@19899.4]
  wire  _T_1119; // @[NV_NVDLA_CSC_dl.scala 280:45:@19902.4]
  wire [14:0] _T_1121; // @[NV_NVDLA_CSC_dl.scala 281:83:@19903.4]
  wire [14:0] _T_1122; // @[NV_NVDLA_CSC_dl.scala 281:25:@19904.4]
  wire  _T_1148; // @[NV_NVDLA_CSC_dl.scala 292:13:@19927.4]
  wire [14:0] _GEN_52; // @[NV_NVDLA_CSC_dl.scala 292:25:@19928.4]
  reg  _T_1166; // @[NV_NVDLA_CSC_dl.scala 308:37:@19948.4]
  reg [31:0] _RAND_51;
  reg [13:0] _T_1169; // @[Reg.scala 19:20:@19951.4]
  reg [31:0] _RAND_52;
  wire [13:0] _GEN_54; // @[Reg.scala 20:19:@19952.4]
  reg [14:0] _T_1172; // @[Reg.scala 19:20:@19956.4]
  reg [31:0] _RAND_53;
  wire [14:0] _GEN_55; // @[Reg.scala 20:19:@19957.4]
  reg  _T_1177; // @[NV_NVDLA_CSC_dl.scala 321:50:@19962.4]
  reg [31:0] _RAND_54;
  reg  _T_1180; // @[NV_NVDLA_CSC_dl.scala 321:50:@19963.4]
  reg [31:0] _RAND_55;
  reg  _T_1183; // @[NV_NVDLA_CSC_dl.scala 321:50:@19964.4]
  reg [31:0] _RAND_56;
  reg  _T_1186; // @[NV_NVDLA_CSC_dl.scala 321:50:@19965.4]
  reg [31:0] _RAND_57;
  reg  _T_1189; // @[NV_NVDLA_CSC_dl.scala 321:50:@19966.4]
  reg [31:0] _RAND_58;
  reg  _T_1211; // @[NV_NVDLA_CSC_dl.scala 340:36:@19996.4]
  reg [31:0] _RAND_59;
  reg  _T_1214; // @[NV_NVDLA_CSC_dl.scala 340:36:@19997.4]
  reg [31:0] _RAND_60;
  reg  _T_1217; // @[NV_NVDLA_CSC_dl.scala 340:36:@19998.4]
  reg [31:0] _RAND_61;
  reg  _T_1220; // @[NV_NVDLA_CSC_dl.scala 340:36:@19999.4]
  reg [31:0] _RAND_62;
  reg [30:0] _T_1225; // @[NV_NVDLA_CSC_dl.scala 342:34:@20001.4]
  reg [31:0] _RAND_63;
  reg [30:0] _T_1228; // @[NV_NVDLA_CSC_dl.scala 342:34:@20002.4]
  reg [31:0] _RAND_64;
  reg [30:0] _T_1231; // @[NV_NVDLA_CSC_dl.scala 342:34:@20003.4]
  reg [31:0] _RAND_65;
  reg [30:0] _T_1234; // @[NV_NVDLA_CSC_dl.scala 342:34:@20004.4]
  reg [31:0] _RAND_66;
  wire [30:0] _T_1222; // @[NV_NVDLA_CSC_dl.scala 341:19:@20000.4 NV_NVDLA_CSC_dl.scala 345:12:@20006.4]
  wire [30:0] _GEN_61; // @[NV_NVDLA_CSC_dl.scala 349:23:@20008.4]
  wire [30:0] _GEN_62; // @[NV_NVDLA_CSC_dl.scala 349:23:@20012.4]
  wire [30:0] _GEN_63; // @[NV_NVDLA_CSC_dl.scala 349:23:@20016.4]
  wire [30:0] _GEN_64; // @[NV_NVDLA_CSC_dl.scala 349:23:@20020.4]
  wire  _T_1235; // @[NV_NVDLA_CSC_dl.scala 354:30:@20023.4]
  wire  _T_1236; // @[NV_NVDLA_CSC_dl.scala 354:34:@20024.4]
  wire  _T_1237; // @[NV_NVDLA_CSC_dl.scala 355:30:@20025.4]
  wire  _T_1238; // @[NV_NVDLA_CSC_dl.scala 355:34:@20026.4]
  wire  _T_1239; // @[NV_NVDLA_CSC_dl.scala 354:50:@20027.4]
  wire  _T_1240; // @[NV_NVDLA_CSC_dl.scala 356:30:@20028.4]
  wire  _T_1241; // @[NV_NVDLA_CSC_dl.scala 356:34:@20029.4]
  wire  _T_1242; // @[NV_NVDLA_CSC_dl.scala 355:50:@20030.4]
  wire  _T_1243; // @[NV_NVDLA_CSC_dl.scala 358:37:@20031.4]
  wire [30:0] _T_1247; // @[Bitwise.scala 72:12:@20033.4]
  wire [30:0] _T_1248; // @[NV_NVDLA_CSC_dl.scala 358:42:@20034.4]
  wire  _T_1249; // @[NV_NVDLA_CSC_dl.scala 359:37:@20035.4]
  wire [30:0] _T_1253; // @[Bitwise.scala 72:12:@20037.4]
  wire [30:0] _T_1254; // @[NV_NVDLA_CSC_dl.scala 359:42:@20038.4]
  wire [30:0] _T_1255; // @[NV_NVDLA_CSC_dl.scala 358:56:@20039.4]
  wire  _T_1256; // @[NV_NVDLA_CSC_dl.scala 360:37:@20040.4]
  wire [30:0] _T_1260; // @[Bitwise.scala 72:12:@20042.4]
  wire [30:0] _T_1261; // @[NV_NVDLA_CSC_dl.scala 360:42:@20043.4]
  wire [30:0] _T_1262; // @[NV_NVDLA_CSC_dl.scala 359:56:@20044.4]
  wire [4:0] _T_1263; // @[NV_NVDLA_CSC_dl.scala 363:24:@20045.4]
  wire [4:0] _T_1264; // @[NV_NVDLA_CSC_dl.scala 364:24:@20046.4]
  wire [6:0] _T_1265; // @[NV_NVDLA_CSC_dl.scala 365:28:@20047.4]
  wire [6:0] _T_1266; // @[NV_NVDLA_CSC_dl.scala 366:29:@20048.4]
  wire [1:0] _T_1267; // @[NV_NVDLA_CSC_dl.scala 367:25:@20049.4]
  wire  _T_1268; // @[NV_NVDLA_CSC_dl.scala 368:25:@20050.4]
  wire  _T_1269; // @[NV_NVDLA_CSC_dl.scala 369:27:@20051.4]
  wire  _T_1270; // @[NV_NVDLA_CSC_dl.scala 370:25:@20052.4]
  wire  _T_1271; // @[NV_NVDLA_CSC_dl.scala 371:25:@20053.4]
  wire  _T_1272; // @[NV_NVDLA_CSC_dl.scala 372:27:@20054.4]
  reg [4:0] _T_1279; // @[NV_NVDLA_CSC_dl.scala 377:24:@20057.4]
  reg [31:0] _RAND_67;
  wire [5:0] _T_1283; // @[NV_NVDLA_CSC_dl.scala 381:24:@20058.4]
  wire [4:0] _T_1284; // @[NV_NVDLA_CSC_dl.scala 381:24:@20059.4]
  wire  _T_1287; // @[NV_NVDLA_CSC_dl.scala 383:27:@20063.4]
  wire [4:0] _T_1285; // @[NV_NVDLA_CSC_dl.scala 380:17:@20060.4]
  wire [4:0] _T_1286; // @[NV_NVDLA_CSC_dl.scala 379:17:@20061.4]
  reg [1:0] _T_1290; // @[NV_NVDLA_CSC_dl.scala 386:24:@20065.4]
  reg [31:0] _RAND_68;
  wire [2:0] _T_1294; // @[NV_NVDLA_CSC_dl.scala 389:31:@20067.4]
  wire [1:0] _T_1295; // @[NV_NVDLA_CSC_dl.scala 389:31:@20068.4]
  wire [2:0] _GEN_682; // @[NV_NVDLA_CSC_dl.scala 390:32:@20069.4]
  wire  _T_1296; // @[NV_NVDLA_CSC_dl.scala 390:32:@20069.4]
  wire  _T_1298; // @[NV_NVDLA_CSC_dl.scala 391:61:@20071.4]
  reg [6:0] _T_1306; // @[NV_NVDLA_CSC_dl.scala 397:25:@20079.4]
  reg [31:0] _RAND_69;
  wire  _T_1346; // @[NV_NVDLA_CSC_dl.scala 424:37:@20108.4]
  wire  _T_1347; // @[NV_NVDLA_CSC_dl.scala 424:24:@20109.4]
  wire  _T_1349; // @[NV_NVDLA_CSC_dl.scala 424:56:@20110.4]
  wire  _T_1350; // @[NV_NVDLA_CSC_dl.scala 424:44:@20111.4]
  wire  _T_1351; // @[NV_NVDLA_CSC_dl.scala 424:42:@20112.4]
  wire  _T_1353; // @[NV_NVDLA_CSC_dl.scala 424:75:@20113.4]
  wire  _T_1354; // @[NV_NVDLA_CSC_dl.scala 424:63:@20114.4]
  wire  _T_1355; // @[NV_NVDLA_CSC_dl.scala 424:61:@20115.4]
  reg  _T_1335; // @[NV_NVDLA_CSC_dl.scala 416:32:@20101.4]
  reg [31:0] _RAND_70;
  wire  _T_1357; // @[NV_NVDLA_CSC_dl.scala 424:22:@20116.4]
  wire  _T_1358; // @[NV_NVDLA_CSC_dl.scala 423:22:@20117.4]
  wire  _T_1299; // @[NV_NVDLA_CSC_dl.scala 391:66:@20072.4]
  wire  _T_1300; // @[NV_NVDLA_CSC_dl.scala 391:33:@20073.4]
  wire  _T_1301; // @[NV_NVDLA_CSC_dl.scala 393:31:@20075.6]
  wire [1:0] _T_1303; // @[NV_NVDLA_CSC_dl.scala 393:21:@20076.6]
  wire [1:0] _GEN_65; // @[NV_NVDLA_CSC_dl.scala 392:23:@20074.4]
  wire [7:0] _T_1312; // @[NV_NVDLA_CSC_dl.scala 401:33:@20082.4]
  wire [6:0] _T_1313; // @[NV_NVDLA_CSC_dl.scala 401:33:@20083.4]
  wire  _T_1314; // @[NV_NVDLA_CSC_dl.scala 402:51:@20084.4]
  wire  _T_1315; // @[NV_NVDLA_CSC_dl.scala 402:33:@20085.4]
  wire  _T_1316; // @[NV_NVDLA_CSC_dl.scala 403:34:@20087.4]
  wire  _T_1317; // @[NV_NVDLA_CSC_dl.scala 404:52:@20089.4]
  wire  _T_1318; // @[NV_NVDLA_CSC_dl.scala 404:34:@20090.4]
  wire  _T_1320; // @[NV_NVDLA_CSC_dl.scala 408:41:@20092.6]
  wire  _T_1321; // @[NV_NVDLA_CSC_dl.scala 408:39:@20093.6]
  wire [6:0] _T_1324; // @[NV_NVDLA_CSC_dl.scala 409:22:@20094.6]
  wire [6:0] _T_1325; // @[NV_NVDLA_CSC_dl.scala 408:22:@20095.6]
  wire [6:0] _T_1326; // @[NV_NVDLA_CSC_dl.scala 407:22:@20096.6]
  wire [6:0] _GEN_66; // @[NV_NVDLA_CSC_dl.scala 406:24:@20091.4]
  reg  _T_1329; // @[NV_NVDLA_CSC_dl.scala 414:35:@20099.4]
  reg [31:0] _RAND_71;
  reg  _T_1332; // @[NV_NVDLA_CSC_dl.scala 415:32:@20100.4]
  reg [31:0] _RAND_72;
  wire  _T_1343; // @[NV_NVDLA_CSC_dl.scala 422:27:@20106.4]
  wire  _T_1338; // @[NV_NVDLA_CSC_dl.scala 419:49:@20103.4]
  wire  _T_1341; // @[NV_NVDLA_CSC_dl.scala 420:32:@20104.4]
  wire  _T_1342; // @[NV_NVDLA_CSC_dl.scala 419:33:@20105.4]
  reg [7:0] _T_1361; // @[NV_NVDLA_CSC_dl.scala 432:31:@20122.4]
  reg [31:0] _RAND_73;
  wire [7:0] _T_1363; // @[Cat.scala 30:58:@20123.4]
  wire [7:0] _GEN_67; // @[NV_NVDLA_CSC_dl.scala 434:21:@20124.4]
  reg [12:0] _T_1366; // @[NV_NVDLA_CSC_dl.scala 440:28:@20127.4]
  reg [31:0] _RAND_74;
  reg [12:0] _T_1369; // @[NV_NVDLA_CSC_dl.scala 441:28:@20128.4]
  reg [31:0] _RAND_75;
  wire [12:0] _GEN_683; // @[NV_NVDLA_CSC_dl.scala 444:39:@20129.4]
  wire [13:0] _T_1370; // @[NV_NVDLA_CSC_dl.scala 444:39:@20129.4]
  wire [12:0] _T_1371; // @[NV_NVDLA_CSC_dl.scala 444:39:@20130.4]
  wire  _T_1372; // @[NV_NVDLA_CSC_dl.scala 445:29:@20131.4]
  wire  _T_1373; // @[NV_NVDLA_CSC_dl.scala 445:61:@20132.4]
  wire  _T_1374; // @[NV_NVDLA_CSC_dl.scala 445:44:@20133.4]
  wire  _T_1377; // @[NV_NVDLA_CSC_dl.scala 448:43:@20136.4]
  wire  _T_1378; // @[NV_NVDLA_CSC_dl.scala 448:41:@20137.4]
  wire [12:0] _T_1379; // @[NV_NVDLA_CSC_dl.scala 449:26:@20138.4]
  wire [12:0] _T_1380; // @[NV_NVDLA_CSC_dl.scala 448:26:@20139.4]
  wire [12:0] _T_1381; // @[NV_NVDLA_CSC_dl.scala 447:26:@20140.4]
  wire  _T_1383; // @[NV_NVDLA_CSC_dl.scala 450:70:@20142.4]
  wire  _T_1384; // @[NV_NVDLA_CSC_dl.scala 450:37:@20143.4]
  wire  _T_1385; // @[NV_NVDLA_CSC_dl.scala 451:55:@20144.4]
  wire  _T_1386; // @[NV_NVDLA_CSC_dl.scala 451:71:@20145.4]
  wire  _T_1387; // @[NV_NVDLA_CSC_dl.scala 451:37:@20146.4]
  wire [12:0] _GEN_68; // @[NV_NVDLA_CSC_dl.scala 453:27:@20147.4]
  wire [12:0] _GEN_69; // @[NV_NVDLA_CSC_dl.scala 456:27:@20150.4]
  reg [10:0] _T_1390; // @[NV_NVDLA_CSC_dl.scala 461:27:@20153.4]
  reg [31:0] _RAND_76;
  wire  _T_1391; // @[NV_NVDLA_CSC_dl.scala 463:37:@20154.4]
  wire  _T_1393; // @[NV_NVDLA_CSC_dl.scala 464:70:@20156.4]
  wire  _T_1394; // @[NV_NVDLA_CSC_dl.scala 464:36:@20157.4]
  wire [11:0] _T_1398; // @[NV_NVDLA_CSC_dl.scala 469:34:@20159.6]
  wire [10:0] _T_1399; // @[NV_NVDLA_CSC_dl.scala 469:34:@20160.6]
  wire [10:0] _T_1400; // @[NV_NVDLA_CSC_dl.scala 468:24:@20161.6]
  wire [10:0] _T_1401; // @[NV_NVDLA_CSC_dl.scala 467:24:@20162.6]
  wire [10:0] _GEN_70; // @[NV_NVDLA_CSC_dl.scala 466:26:@20158.4]
  reg [13:0] _T_1404; // @[NV_NVDLA_CSC_dl.scala 473:27:@20165.4]
  reg [31:0] _RAND_77;
  reg [13:0] _T_1407; // @[NV_NVDLA_CSC_dl.scala 474:27:@20166.4]
  reg [31:0] _RAND_78;
  reg [15:0] _T_1410; // @[NV_NVDLA_CSC_dl.scala 475:26:@20167.4]
  reg [31:0] _RAND_79;
  reg [15:0] _T_1413; // @[NV_NVDLA_CSC_dl.scala 476:26:@20168.4]
  reg [31:0] _RAND_80;
  reg [15:0] _T_1416; // @[NV_NVDLA_CSC_dl.scala 477:29:@20169.4]
  reg [31:0] _RAND_81;
  reg [12:0] _T_1419; // @[NV_NVDLA_CSC_dl.scala 478:29:@20170.4]
  reg [31:0] _RAND_82;
  reg  _T_1424; // @[NV_NVDLA_CSC_dl.scala 480:33:@20172.4]
  reg [31:0] _RAND_83;
  reg  _T_1427; // @[NV_NVDLA_CSC_dl.scala 481:35:@20173.4]
  reg [31:0] _RAND_84;
  wire [12:0] _GEN_684; // @[NV_NVDLA_CSC_dl.scala 484:41:@20174.4]
  wire [13:0] _T_1430; // @[NV_NVDLA_CSC_dl.scala 484:41:@20174.4]
  wire [13:0] _T_1431; // @[NV_NVDLA_CSC_dl.scala 484:41:@20175.4]
  wire [13:0] _T_1432; // @[NV_NVDLA_CSC_dl.scala 483:26:@20176.4]
  wire [13:0] _GEN_685; // @[NV_NVDLA_CSC_dl.scala 485:37:@20177.4]
  wire [14:0] _T_1433; // @[NV_NVDLA_CSC_dl.scala 485:37:@20177.4]
  wire [13:0] _T_1434; // @[NV_NVDLA_CSC_dl.scala 485:37:@20178.4]
  wire [13:0] _T_1437; // @[NV_NVDLA_CSC_dl.scala 490:25:@20181.4]
  wire [13:0] _T_1438; // @[NV_NVDLA_CSC_dl.scala 489:25:@20182.4]
  wire [13:0] _T_1439; // @[NV_NVDLA_CSC_dl.scala 488:25:@20183.4]
  wire [5:0] _GEN_686; // @[NV_NVDLA_CSC_dl.scala 492:35:@20184.4]
  wire [10:0] _T_1440; // @[NV_NVDLA_CSC_dl.scala 492:35:@20184.4]
  wire [13:0] _GEN_687; // @[NV_NVDLA_CSC_dl.scala 493:33:@20185.4]
  wire [14:0] _T_1441; // @[NV_NVDLA_CSC_dl.scala 493:33:@20185.4]
  wire [13:0] _T_1442; // @[NV_NVDLA_CSC_dl.scala 493:33:@20186.4]
  wire  _T_1445; // @[NV_NVDLA_CSC_dl.scala 494:96:@20189.4]
  wire  _T_1446; // @[NV_NVDLA_CSC_dl.scala 494:86:@20190.4]
  wire  _T_1447; // @[NV_NVDLA_CSC_dl.scala 494:84:@20191.4]
  wire  _T_1448; // @[NV_NVDLA_CSC_dl.scala 494:36:@20192.4]
  wire  _T_1451; // @[NV_NVDLA_CSC_dl.scala 495:99:@20195.4]
  wire  _T_1452; // @[NV_NVDLA_CSC_dl.scala 495:89:@20196.4]
  wire  _T_1453; // @[NV_NVDLA_CSC_dl.scala 495:87:@20197.4]
  wire  _T_1454; // @[NV_NVDLA_CSC_dl.scala 495:36:@20198.4]
  wire [7:0] _T_1456; // @[NV_NVDLA_CSC_dl.scala 498:26:@20199.4]
  wire  _T_1459; // @[NV_NVDLA_CSC_dl.scala 500:79:@20201.4]
  wire [7:0] _T_1463; // @[NV_NVDLA_CSC_dl.scala 501:74:@20204.4]
  wire [6:0] _T_1464; // @[NV_NVDLA_CSC_dl.scala 501:74:@20205.4]
  wire [6:0] _T_1465; // @[NV_NVDLA_CSC_dl.scala 500:27:@20206.4]
  wire  _T_1466; // @[NV_NVDLA_CSC_dl.scala 502:37:@20207.4]
  wire  _T_1468; // @[NV_NVDLA_CSC_dl.scala 503:35:@20208.4]
  wire [13:0] _T_1470; // @[NV_NVDLA_CSC_dl.scala 503:66:@20209.4]
  wire [12:0] _T_1471; // @[NV_NVDLA_CSC_dl.scala 503:66:@20210.4]
  wire [12:0] _T_1472; // @[NV_NVDLA_CSC_dl.scala 503:22:@20211.4]
  wire [12:0] _T_1473; // @[NV_NVDLA_CSC_dl.scala 502:22:@20212.4]
  wire [12:0] _GEN_688; // @[NV_NVDLA_CSC_dl.scala 505:44:@20214.4]
  wire  _T_1474; // @[NV_NVDLA_CSC_dl.scala 505:44:@20214.4]
  wire  _T_1475; // @[NV_NVDLA_CSC_dl.scala 509:39:@20215.4]
  wire  _T_1476; // @[NV_NVDLA_CSC_dl.scala 509:54:@20216.4]
  wire  _T_1477; // @[NV_NVDLA_CSC_dl.scala 509:71:@20217.4]
  wire  _T_1480; // @[NV_NVDLA_CSC_dl.scala 510:73:@20220.4]
  wire  _T_1481; // @[NV_NVDLA_CSC_dl.scala 510:71:@20221.4]
  wire [15:0] _GEN_689; // @[NV_NVDLA_CSC_dl.scala 510:99:@20222.4]
  wire [16:0] _T_1482; // @[NV_NVDLA_CSC_dl.scala 510:99:@20222.4]
  wire [15:0] _T_1483; // @[NV_NVDLA_CSC_dl.scala 510:99:@20223.4]
  wire  _T_1485; // @[NV_NVDLA_CSC_dl.scala 511:54:@20225.4]
  wire [15:0] _GEN_690; // @[NV_NVDLA_CSC_dl.scala 511:90:@20226.4]
  wire [16:0] _T_1486; // @[NV_NVDLA_CSC_dl.scala 511:90:@20226.4]
  wire [15:0] _T_1487; // @[NV_NVDLA_CSC_dl.scala 511:90:@20227.4]
  wire  _T_1489; // @[NV_NVDLA_CSC_dl.scala 512:56:@20229.4]
  wire  _T_1490; // @[NV_NVDLA_CSC_dl.scala 512:54:@20230.4]
  wire [16:0] _T_1492; // @[NV_NVDLA_CSC_dl.scala 512:91:@20231.4]
  wire [15:0] _T_1493; // @[NV_NVDLA_CSC_dl.scala 512:91:@20232.4]
  wire  _T_1494; // @[NV_NVDLA_CSC_dl.scala 513:41:@20233.4]
  wire  _T_1495; // @[NV_NVDLA_CSC_dl.scala 513:39:@20234.4]
  wire [15:0] _GEN_691; // @[NV_NVDLA_CSC_dl.scala 513:81:@20235.4]
  wire [16:0] _T_1496; // @[NV_NVDLA_CSC_dl.scala 513:81:@20235.4]
  wire [15:0] _T_1497; // @[NV_NVDLA_CSC_dl.scala 513:81:@20236.4]
  wire [15:0] _T_1498; // @[NV_NVDLA_CSC_dl.scala 513:24:@20237.4]
  wire [15:0] _T_1499; // @[NV_NVDLA_CSC_dl.scala 512:24:@20238.4]
  wire [15:0] _T_1500; // @[NV_NVDLA_CSC_dl.scala 511:24:@20239.4]
  wire [15:0] _T_1501; // @[NV_NVDLA_CSC_dl.scala 510:24:@20240.4]
  wire [15:0] _T_1502; // @[NV_NVDLA_CSC_dl.scala 509:24:@20241.4]
  wire [15:0] _T_1503; // @[NV_NVDLA_CSC_dl.scala 508:24:@20242.4]
  wire [9:0] _T_1509; // @[NV_NVDLA_CSC_dl.scala 515:68:@20244.4]
  wire [14:0] _T_1510; // @[Cat.scala 30:58:@20245.4]
  wire  _T_1521; // @[NV_NVDLA_CSC_dl.scala 518:68:@20256.4]
  wire  _T_1522; // @[NV_NVDLA_CSC_dl.scala 518:57:@20257.4]
  wire  _T_1523; // @[NV_NVDLA_CSC_dl.scala 518:72:@20258.4]
  wire  _T_1524; // @[NV_NVDLA_CSC_dl.scala 518:88:@20259.4]
  wire  _T_1525; // @[NV_NVDLA_CSC_dl.scala 518:103:@20260.4]
  wire  _T_1526; // @[NV_NVDLA_CSC_dl.scala 518:39:@20261.4]
  wire  _T_1528; // @[NV_NVDLA_CSC_dl.scala 520:42:@20263.4]
  wire  _T_1531; // @[NV_NVDLA_CSC_dl.scala 520:74:@20264.4]
  wire  _T_1532; // @[NV_NVDLA_CSC_dl.scala 520:28:@20265.4]
  wire  _T_1534; // @[NV_NVDLA_CSC_dl.scala 521:36:@20267.4]
  wire  _T_1535; // @[NV_NVDLA_CSC_dl.scala 521:72:@20268.4]
  wire  _T_1536; // @[NV_NVDLA_CSC_dl.scala 521:51:@20269.4]
  wire [13:0] _GEN_71; // @[NV_NVDLA_CSC_dl.scala 523:26:@20270.4]
  wire [15:0] _GEN_72; // @[NV_NVDLA_CSC_dl.scala 523:26:@20270.4]
  wire [13:0] _GEN_73; // @[NV_NVDLA_CSC_dl.scala 527:26:@20274.4]
  wire [15:0] _GEN_74; // @[NV_NVDLA_CSC_dl.scala 527:26:@20274.4]
  wire [15:0] _GEN_75; // @[NV_NVDLA_CSC_dl.scala 531:26:@20278.4]
  reg [13:0] _T_1539; // @[NV_NVDLA_CSC_dl.scala 537:27:@20281.4]
  reg [31:0] _RAND_85;
  reg [13:0] _T_1542; // @[NV_NVDLA_CSC_dl.scala 538:27:@20282.4]
  reg [31:0] _RAND_86;
  wire [13:0] _GEN_692; // @[NV_NVDLA_CSC_dl.scala 540:41:@20283.4]
  wire [14:0] _T_1544; // @[NV_NVDLA_CSC_dl.scala 540:41:@20283.4]
  wire [14:0] _T_1545; // @[NV_NVDLA_CSC_dl.scala 540:41:@20284.4]
  wire [13:0] _T_1546; // @[NV_NVDLA_CSC_dl.scala 540:41:@20285.4]
  wire [13:0] _GEN_693; // @[NV_NVDLA_CSC_dl.scala 541:37:@20286.4]
  wire [14:0] _T_1547; // @[NV_NVDLA_CSC_dl.scala 541:37:@20286.4]
  wire [13:0] _T_1548; // @[NV_NVDLA_CSC_dl.scala 541:37:@20287.4]
  wire  _T_1549; // @[NV_NVDLA_CSC_dl.scala 542:52:@20288.4]
  wire  _T_1550; // @[NV_NVDLA_CSC_dl.scala 542:35:@20289.4]
  wire [13:0] _T_1553; // @[NV_NVDLA_CSC_dl.scala 544:25:@20292.4]
  wire [13:0] _T_1554; // @[NV_NVDLA_CSC_dl.scala 543:25:@20293.4]
  wire [13:0] _T_1555; // @[NV_NVDLA_CSC_dl.scala 542:25:@20294.4]
  wire  _T_1558; // @[NV_NVDLA_CSC_dl.scala 545:91:@20297.4]
  wire  _T_1559; // @[NV_NVDLA_CSC_dl.scala 545:54:@20298.4]
  wire  _T_1560; // @[NV_NVDLA_CSC_dl.scala 545:36:@20299.4]
  wire [5:0] _GEN_694; // @[NV_NVDLA_CSC_dl.scala 547:35:@20303.4]
  wire [10:0] _T_1564; // @[NV_NVDLA_CSC_dl.scala 547:35:@20303.4]
  wire [13:0] _GEN_695; // @[NV_NVDLA_CSC_dl.scala 548:33:@20304.4]
  wire [14:0] _T_1565; // @[NV_NVDLA_CSC_dl.scala 548:33:@20304.4]
  wire [13:0] _T_1566; // @[NV_NVDLA_CSC_dl.scala 548:33:@20305.4]
  wire [13:0] _GEN_696; // @[NV_NVDLA_CSC_dl.scala 548:51:@20306.4]
  wire [14:0] _T_1567; // @[NV_NVDLA_CSC_dl.scala 548:51:@20306.4]
  wire [13:0] _T_1568; // @[NV_NVDLA_CSC_dl.scala 548:51:@20307.4]
  wire [13:0] _GEN_76; // @[NV_NVDLA_CSC_dl.scala 550:26:@20308.4]
  wire [13:0] _GEN_77; // @[NV_NVDLA_CSC_dl.scala 551:26:@20311.4]
  wire  _T_1569; // @[NV_NVDLA_CSC_dl.scala 554:39:@20314.4]
  wire [13:0] _GEN_697; // @[NV_NVDLA_CSC_dl.scala 554:59:@20315.4]
  wire  _T_1570; // @[NV_NVDLA_CSC_dl.scala 554:59:@20315.4]
  wire  _T_1571; // @[NV_NVDLA_CSC_dl.scala 554:44:@20316.4]
  wire  _T_1572; // @[NV_NVDLA_CSC_dl.scala 554:92:@20317.4]
  wire  _T_1573; // @[NV_NVDLA_CSC_dl.scala 554:78:@20318.4]
  wire [13:0] _GEN_698; // @[NV_NVDLA_CSC_dl.scala 554:112:@20319.4]
  wire  _T_1574; // @[NV_NVDLA_CSC_dl.scala 554:112:@20319.4]
  wire  _T_1575; // @[NV_NVDLA_CSC_dl.scala 554:97:@20320.4]
  wire  _T_1588; // @[NV_NVDLA_CSC_dl.scala 557:42:@20330.4]
  wire  _T_1698; // @[NV_NVDLA_CSC_dl.scala 642:33:@20416.4]
  wire  _T_1699; // @[NV_NVDLA_CSC_dl.scala 643:24:@20417.4]
  wire [12:0] _T_1701; // @[NV_NVDLA_CSC_dl.scala 643:77:@20418.4]
  wire [14:0] _T_1702; // @[Cat.scala 30:58:@20419.4]
  wire  _T_1704; // @[NV_NVDLA_CSC_dl.scala 644:38:@20420.4]
  wire [11:0] _T_1709; // @[NV_NVDLA_CSC_dl.scala 645:54:@20423.4]
  wire [14:0] _T_1710; // @[Cat.scala 30:58:@20424.4]
  wire [14:0] _T_1711; // @[NV_NVDLA_CSC_dl.scala 644:23:@20425.4]
  wire [14:0] _T_1712; // @[NV_NVDLA_CSC_dl.scala 643:23:@20426.4]
  wire [14:0] _T_1713; // @[NV_NVDLA_CSC_dl.scala 642:23:@20427.4]
  wire [13:0] _T_1714; // @[NV_NVDLA_CSC_dl.scala 654:24:@20429.4]
  wire [11:0] _T_1591; // @[NV_NVDLA_CSC_dl.scala 561:32:@20332.4]
  wire [14:0] _GEN_700; // @[NV_NVDLA_CSC_dl.scala 561:40:@20333.4]
  wire  _T_1592; // @[NV_NVDLA_CSC_dl.scala 561:40:@20333.4]
  wire  _T_1593; // @[NV_NVDLA_CSC_dl.scala 562:34:@20334.4]
  wire  _T_1594; // @[NV_NVDLA_CSC_dl.scala 562:24:@20335.4]
  wire  _T_1595; // @[NV_NVDLA_CSC_dl.scala 563:29:@20336.4]
  wire  _T_1596; // @[NV_NVDLA_CSC_dl.scala 563:33:@20337.4]
  wire  _T_1597; // @[NV_NVDLA_CSC_dl.scala 564:39:@20338.4]
  wire  _T_1598; // @[NV_NVDLA_CSC_dl.scala 564:37:@20339.4]
  wire  _T_1599; // @[NV_NVDLA_CSC_dl.scala 564:56:@20340.4]
  wire  _T_1600; // @[NV_NVDLA_CSC_dl.scala 564:54:@20341.4]
  wire  _T_1601; // @[NV_NVDLA_CSC_dl.scala 567:37:@20342.4]
  wire  _T_1602; // @[NV_NVDLA_CSC_dl.scala 567:27:@20343.4]
  wire  _T_1603; // @[NV_NVDLA_CSC_dl.scala 567:54:@20344.4]
  wire  _T_1604; // @[NV_NVDLA_CSC_dl.scala 567:26:@20345.4]
  wire [1:0] _T_1605; // @[NV_NVDLA_CSC_dl.scala 568:35:@20346.4]
  wire  _T_1607; // @[NV_NVDLA_CSC_dl.scala 569:55:@20347.4]
  wire  _T_1608; // @[NV_NVDLA_CSC_dl.scala 569:42:@20348.4]
  wire  _T_1609; // @[NV_NVDLA_CSC_dl.scala 572:42:@20350.4]
  wire [8:0] _T_1613; // @[Cat.scala 30:58:@20354.4]
  reg  _T_1616; // @[NV_NVDLA_CSC_dl.scala 579:31:@20355.4]
  reg [31:0] _RAND_87;
  reg [1:0] _T_1619; // @[NV_NVDLA_CSC_dl.scala 580:31:@20356.4]
  reg [31:0] _RAND_88;
  reg [1:0] _T_1622; // @[NV_NVDLA_CSC_dl.scala 581:31:@20357.4]
  reg [31:0] _RAND_89;
  reg  _T_1625; // @[NV_NVDLA_CSC_dl.scala 582:31:@20358.4]
  reg [31:0] _RAND_90;
  reg  _T_1628; // @[NV_NVDLA_CSC_dl.scala 583:32:@20359.4]
  reg [31:0] _RAND_91;
  reg  _T_1631; // @[NV_NVDLA_CSC_dl.scala 584:31:@20360.4]
  reg [31:0] _RAND_92;
  reg [1:0] _T_1634; // @[NV_NVDLA_CSC_dl.scala 585:35:@20361.4]
  reg [31:0] _RAND_93;
  reg  _T_1637; // @[NV_NVDLA_CSC_dl.scala 586:34:@20362.4]
  reg [31:0] _RAND_94;
  reg [8:0] _T_1640; // @[NV_NVDLA_CSC_dl.scala 587:30:@20363.4]
  reg [31:0] _RAND_95;
  reg  _T_1643; // @[NV_NVDLA_CSC_dl.scala 588:29:@20364.4]
  reg [31:0] _RAND_96;
  wire  _T_1644; // @[NV_NVDLA_CSC_dl.scala 599:38:@20374.6]
  wire  _T_1645; // @[NV_NVDLA_CSC_dl.scala 599:56:@20375.6]
  wire [1:0] _GEN_78; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  wire [1:0] _GEN_79; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  wire  _GEN_80; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  wire  _GEN_81; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  wire  _GEN_82; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  wire [1:0] _GEN_83; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  wire [8:0] _GEN_84; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  wire  _GEN_85; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  wire  _GEN_86; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  wire  _GEN_87; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  wire  _GEN_88; // @[NV_NVDLA_CSC_dl.scala 603:26:@20380.4]
  reg [12:0] _T_1648; // @[NV_NVDLA_CSC_dl.scala 611:21:@20383.4]
  reg [31:0] _RAND_97;
  reg [12:0] _T_1651; // @[NV_NVDLA_CSC_dl.scala 612:24:@20384.4]
  reg [31:0] _RAND_98;
  reg [12:0] _T_1654; // @[NV_NVDLA_CSC_dl.scala 613:26:@20385.4]
  reg [31:0] _RAND_99;
  reg [12:0] _T_1657; // @[NV_NVDLA_CSC_dl.scala 614:26:@20386.4]
  reg [31:0] _RAND_100;
  reg [12:0] _T_1660; // @[NV_NVDLA_CSC_dl.scala 615:26:@20387.4]
  reg [31:0] _RAND_101;
  reg [12:0] _T_1663; // @[NV_NVDLA_CSC_dl.scala 616:26:@20388.4]
  reg [31:0] _RAND_102;
  reg [12:0] _T_1666; // @[NV_NVDLA_CSC_dl.scala 617:24:@20389.4]
  reg [31:0] _RAND_103;
  wire  _T_1667; // @[NV_NVDLA_CSC_dl.scala 620:32:@20390.4]
  wire  _T_1668; // @[NV_NVDLA_CSC_dl.scala 620:22:@20391.4]
  wire [11:0] _T_1669; // @[NV_NVDLA_CSC_dl.scala 620:49:@20392.4]
  wire [11:0] _T_1671; // @[NV_NVDLA_CSC_dl.scala 620:21:@20393.4]
  wire  _T_1673; // @[NV_NVDLA_CSC_dl.scala 622:34:@20394.4]
  wire [12:0] _GEN_701; // @[NV_NVDLA_CSC_dl.scala 622:64:@20395.4]
  wire [13:0] _T_1675; // @[NV_NVDLA_CSC_dl.scala 622:64:@20395.4]
  wire [12:0] _T_1676; // @[NV_NVDLA_CSC_dl.scala 622:64:@20396.4]
  wire [12:0] _T_1677; // @[NV_NVDLA_CSC_dl.scala 622:19:@20397.4]
  wire [12:0] _T_1678; // @[NV_NVDLA_CSC_dl.scala 621:19:@20398.4]
  wire  _T_1682; // @[NV_NVDLA_CSC_dl.scala 624:31:@20402.4]
  wire [13:0] _GEN_702; // @[NV_NVDLA_CSC_dl.scala 627:32:@20403.4]
  wire [25:0] _T_1683; // @[NV_NVDLA_CSC_dl.scala 627:32:@20403.4]
  wire [12:0] _T_1684; // @[NV_NVDLA_CSC_dl.scala 627:50:@20404.4]
  wire [11:0] _GEN_703; // @[NV_NVDLA_CSC_dl.scala 628:31:@20405.4]
  wire [16:0] _T_1685; // @[NV_NVDLA_CSC_dl.scala 628:31:@20405.4]
  wire [12:0] _T_1686; // @[NV_NVDLA_CSC_dl.scala 628:49:@20406.4]
  wire [14:0] _GEN_704; // @[NV_NVDLA_CSC_dl.scala 629:29:@20407.4]
  wire [19:0] _T_1687; // @[NV_NVDLA_CSC_dl.scala 629:29:@20407.4]
  wire [12:0] _T_1688; // @[NV_NVDLA_CSC_dl.scala 629:47:@20408.4]
  wire [14:0] _GEN_705; // @[NV_NVDLA_CSC_dl.scala 630:47:@20409.4]
  wire [16:0] _T_1690; // @[NV_NVDLA_CSC_dl.scala 630:47:@20409.4]
  wire [16:0] _T_1691; // @[NV_NVDLA_CSC_dl.scala 630:21:@20410.4]
  wire [12:0] _T_1692; // @[NV_NVDLA_CSC_dl.scala 630:65:@20411.4]
  wire  _T_1693; // @[NV_NVDLA_CSC_dl.scala 631:45:@20412.4]
  wire  _T_1694; // @[NV_NVDLA_CSC_dl.scala 631:34:@20413.4]
  wire [1:0] _T_1695; // @[Cat.scala 30:58:@20414.4]
  wire [12:0] _GEN_89; // @[NV_NVDLA_CSC_dl.scala 658:20:@20431.4]
  wire [12:0] _GEN_90; // @[NV_NVDLA_CSC_dl.scala 661:23:@20434.4]
  wire  _T_1715; // @[NV_NVDLA_CSC_dl.scala 664:19:@20437.4]
  wire [12:0] _GEN_91; // @[NV_NVDLA_CSC_dl.scala 664:23:@20438.4]
  wire [12:0] _GEN_92; // @[NV_NVDLA_CSC_dl.scala 664:23:@20438.4]
  wire [12:0] _GEN_93; // @[NV_NVDLA_CSC_dl.scala 664:23:@20438.4]
  wire  _T_1716; // @[NV_NVDLA_CSC_dl.scala 669:19:@20443.4]
  wire [12:0] _GEN_94; // @[NV_NVDLA_CSC_dl.scala 669:23:@20444.4]
  wire [13:0] _GEN_95; // @[NV_NVDLA_CSC_dl.scala 672:20:@20447.4]
  reg [12:0] _T_1759_0; // @[NV_NVDLA_CSC_dl.scala 680:33:@20459.4]
  reg [31:0] _RAND_104;
  reg [12:0] _T_1759_1; // @[NV_NVDLA_CSC_dl.scala 680:33:@20459.4]
  reg [31:0] _RAND_105;
  reg [12:0] _T_1759_2; // @[NV_NVDLA_CSC_dl.scala 680:33:@20459.4]
  reg [31:0] _RAND_106;
  reg [12:0] _T_1759_3; // @[NV_NVDLA_CSC_dl.scala 680:33:@20459.4]
  reg [31:0] _RAND_107;
  reg  _T_1778; // @[NV_NVDLA_CSC_dl.scala 681:35:@20460.4]
  reg [31:0] _RAND_108;
  reg [14:0] _T_1785; // @[NV_NVDLA_CSC_dl.scala 682:37:@20462.4]
  reg [31:0] _RAND_109;
  reg  _T_1788; // @[NV_NVDLA_CSC_dl.scala 683:32:@20463.4]
  reg [31:0] _RAND_110;
  reg [1:0] _T_1794; // @[NV_NVDLA_CSC_dl.scala 685:33:@20465.4]
  reg [31:0] _RAND_111;
  reg [1:0] _T_1797; // @[NV_NVDLA_CSC_dl.scala 686:33:@20466.4]
  reg [31:0] _RAND_112;
  reg  _T_1800; // @[NV_NVDLA_CSC_dl.scala 687:33:@20467.4]
  reg [31:0] _RAND_113;
  reg  _T_1803; // @[NV_NVDLA_CSC_dl.scala 688:34:@20468.4]
  reg [31:0] _RAND_114;
  reg [7:0] _T_1806; // @[NV_NVDLA_CSC_dl.scala 689:33:@20469.4]
  reg [31:0] _RAND_115;
  reg  _T_1809; // @[NV_NVDLA_CSC_dl.scala 690:33:@20470.4]
  reg [31:0] _RAND_116;
  reg [1:0] _T_1812; // @[NV_NVDLA_CSC_dl.scala 691:37:@20471.4]
  reg [31:0] _RAND_117;
  reg  _T_1815; // @[NV_NVDLA_CSC_dl.scala 692:36:@20472.4]
  reg [31:0] _RAND_118;
  reg  _T_1818; // @[NV_NVDLA_CSC_dl.scala 693:31:@20473.4]
  reg [31:0] _RAND_119;
  reg [8:0] _T_1821; // @[NV_NVDLA_CSC_dl.scala 694:32:@20474.4]
  reg [31:0] _RAND_120;
  wire [13:0] _T_1822; // @[NV_NVDLA_CSC_dl.scala 696:29:@20475.4]
  wire [12:0] _T_1823; // @[NV_NVDLA_CSC_dl.scala 696:29:@20476.4]
  wire [13:0] _T_1824; // @[NV_NVDLA_CSC_dl.scala 696:43:@20477.4]
  wire [12:0] _T_1825; // @[NV_NVDLA_CSC_dl.scala 696:43:@20478.4]
  wire [13:0] _T_1826; // @[NV_NVDLA_CSC_dl.scala 696:57:@20479.4]
  wire [12:0] _T_1827; // @[NV_NVDLA_CSC_dl.scala 696:57:@20480.4]
  wire [14:0] _GEN_706; // @[NV_NVDLA_CSC_dl.scala 697:40:@20481.4]
  wire [15:0] _T_1828; // @[NV_NVDLA_CSC_dl.scala 697:40:@20481.4]
  wire [14:0] _T_1829; // @[NV_NVDLA_CSC_dl.scala 697:40:@20482.4]
  wire [14:0] _GEN_707; // @[NV_NVDLA_CSC_dl.scala 697:52:@20483.4]
  wire [15:0] _T_1830; // @[NV_NVDLA_CSC_dl.scala 697:52:@20483.4]
  wire [14:0] _T_1831; // @[NV_NVDLA_CSC_dl.scala 697:52:@20484.4]
  wire [14:0] _GEN_708; // @[NV_NVDLA_CSC_dl.scala 697:64:@20485.4]
  wire [15:0] _T_1832; // @[NV_NVDLA_CSC_dl.scala 697:64:@20485.4]
  wire [14:0] _T_1833; // @[NV_NVDLA_CSC_dl.scala 697:64:@20486.4]
  wire  _T_1840; // @[NV_NVDLA_CSC_dl.scala 698:45:@20489.4]
  wire [15:0] _T_1847; // @[NV_NVDLA_CSC_dl.scala 699:42:@20492.4]
  wire [15:0] _T_1848; // @[NV_NVDLA_CSC_dl.scala 699:42:@20493.4]
  wire [14:0] _T_1849; // @[NV_NVDLA_CSC_dl.scala 699:42:@20494.4]
  wire  _T_1850; // @[NV_NVDLA_CSC_dl.scala 700:35:@20495.4]
  wire [14:0] _T_1856; // @[NV_NVDLA_CSC_dl.scala 701:25:@20497.4]
  wire [14:0] _T_1857; // @[NV_NVDLA_CSC_dl.scala 700:25:@20498.4]
  wire  _T_1881; // @[Mux.scala 46:19:@20508.4]
  wire [12:0] _T_1882; // @[Mux.scala 46:16:@20509.4]
  wire  _T_1883; // @[Mux.scala 46:19:@20510.4]
  wire [12:0] _T_1884; // @[Mux.scala 46:16:@20511.4]
  wire  _T_1885; // @[Mux.scala 46:19:@20512.4]
  wire [12:0] _T_1886; // @[Mux.scala 46:16:@20513.4]
  wire  _T_1887; // @[Mux.scala 46:19:@20514.4]
  wire [12:0] _T_1888; // @[Mux.scala 46:16:@20515.4]
  wire [14:0] _GEN_712; // @[NV_NVDLA_CSC_dl.scala 708:65:@20516.4]
  wire  _T_1889; // @[NV_NVDLA_CSC_dl.scala 708:65:@20516.4]
  wire  _T_1890; // @[NV_NVDLA_CSC_dl.scala 708:85:@20517.4]
  wire  _T_1891; // @[NV_NVDLA_CSC_dl.scala 708:43:@20518.4]
  wire  _T_1892; // @[NV_NVDLA_CSC_dl.scala 710:38:@20519.4]
  wire  _T_1894; // @[NV_NVDLA_CSC_dl.scala 710:78:@20520.4]
  wire  _T_1895; // @[NV_NVDLA_CSC_dl.scala 710:58:@20521.4]
  wire  _T_1896; // @[NV_NVDLA_CSC_dl.scala 710:17:@20522.4]
  wire  _T_1899; // @[NV_NVDLA_CSC_dl.scala 710:78:@20524.4]
  wire  _T_1900; // @[NV_NVDLA_CSC_dl.scala 710:58:@20525.4]
  wire  _T_1901; // @[NV_NVDLA_CSC_dl.scala 710:17:@20526.4]
  wire  _T_1904; // @[NV_NVDLA_CSC_dl.scala 710:78:@20528.4]
  wire  _T_1905; // @[NV_NVDLA_CSC_dl.scala 710:58:@20529.4]
  wire  _T_1906; // @[NV_NVDLA_CSC_dl.scala 710:17:@20530.4]
  wire  _T_1909; // @[NV_NVDLA_CSC_dl.scala 710:78:@20532.4]
  wire  _T_1910; // @[NV_NVDLA_CSC_dl.scala 710:58:@20533.4]
  wire  _T_1911; // @[NV_NVDLA_CSC_dl.scala 710:17:@20534.4]
  wire [14:0] _GEN_96; // @[NV_NVDLA_CSC_dl.scala 717:35:@20540.4]
  wire [14:0] _GEN_97; // @[NV_NVDLA_CSC_dl.scala 717:35:@20543.4]
  wire [14:0] _GEN_98; // @[NV_NVDLA_CSC_dl.scala 717:35:@20546.4]
  wire [14:0] _GEN_99; // @[NV_NVDLA_CSC_dl.scala 717:35:@20549.4]
  wire  _T_1922; // @[NV_NVDLA_CSC_dl.scala 723:14:@20553.4]
  wire [14:0] _GEN_100; // @[NV_NVDLA_CSC_dl.scala 723:34:@20554.4]
  wire [1:0] _GEN_101; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  wire [1:0] _GEN_102; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  wire  _GEN_103; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  wire  _GEN_104; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  wire [7:0] _GEN_105; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  wire  _GEN_106; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  wire [1:0] _GEN_107; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  wire  _GEN_108; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  wire  _GEN_109; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  wire [8:0] _GEN_110; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  wire [6:0] _T_1932; // @[Cat.scala 30:58:@20581.4]
  wire [28:0] _T_1938; // @[Cat.scala 30:58:@20587.4]
  reg  _T_1943; // @[NV_NVDLA_CSC_dl.scala 757:73:@20589.4]
  reg [31:0] _RAND_121;
  reg  _T_1946; // @[NV_NVDLA_CSC_dl.scala 757:73:@20590.4]
  reg [31:0] _RAND_122;
  reg  _T_1949; // @[NV_NVDLA_CSC_dl.scala 757:73:@20591.4]
  reg [31:0] _RAND_123;
  reg  _T_1952; // @[NV_NVDLA_CSC_dl.scala 757:73:@20592.4]
  reg [31:0] _RAND_124;
  reg  _T_1955; // @[NV_NVDLA_CSC_dl.scala 757:73:@20593.4]
  reg [31:0] _RAND_125;
  reg  _T_1958; // @[NV_NVDLA_CSC_dl.scala 757:73:@20594.4]
  reg [31:0] _RAND_126;
  reg [28:0] _T_1963; // @[NV_NVDLA_CSC_dl.scala 759:71:@20596.4]
  reg [31:0] _RAND_127;
  reg [28:0] _T_1966; // @[NV_NVDLA_CSC_dl.scala 759:71:@20597.4]
  reg [31:0] _RAND_128;
  reg [28:0] _T_1969; // @[NV_NVDLA_CSC_dl.scala 759:71:@20598.4]
  reg [31:0] _RAND_129;
  reg [28:0] _T_1972; // @[NV_NVDLA_CSC_dl.scala 759:71:@20599.4]
  reg [31:0] _RAND_130;
  reg [28:0] _T_1975; // @[NV_NVDLA_CSC_dl.scala 759:71:@20600.4]
  reg [31:0] _RAND_131;
  reg [28:0] _T_1978; // @[NV_NVDLA_CSC_dl.scala 759:71:@20601.4]
  reg [31:0] _RAND_132;
  wire [28:0] _GEN_111; // @[NV_NVDLA_CSC_dl.scala 775:33:@20629.4]
  wire [28:0] _GEN_114; // @[NV_NVDLA_CSC_dl.scala 775:33:@20638.4]
  wire [28:0] _GEN_117; // @[NV_NVDLA_CSC_dl.scala 775:33:@20647.4]
  wire [28:0] _GEN_120; // @[NV_NVDLA_CSC_dl.scala 775:33:@20656.4]
  wire [28:0] _GEN_123; // @[NV_NVDLA_CSC_dl.scala 775:33:@20665.4]
  wire [28:0] _GEN_126; // @[NV_NVDLA_CSC_dl.scala 775:33:@20674.4]
  wire [1:0] _T_2039; // @[NV_NVDLA_CSC_dl.scala 792:41:@20682.4]
  wire [1:0] _T_2040; // @[NV_NVDLA_CSC_dl.scala 793:41:@20683.4]
  wire  _T_2041; // @[NV_NVDLA_CSC_dl.scala 794:41:@20684.4]
  wire  _T_2042; // @[NV_NVDLA_CSC_dl.scala 795:42:@20685.4]
  wire [7:0] _T_2043; // @[NV_NVDLA_CSC_dl.scala 796:41:@20686.4]
  wire [1:0] _T_2044; // @[NV_NVDLA_CSC_dl.scala 797:45:@20687.4]
  wire  _T_2047; // @[NV_NVDLA_CSC_dl.scala 800:39:@20690.4]
  wire [8:0] _T_2048; // @[NV_NVDLA_CSC_dl.scala 801:40:@20691.4]
  reg  _T_2051; // @[NV_NVDLA_CSC_dl.scala 806:29:@20692.4]
  reg [31:0] _RAND_133;
  reg  _T_2063; // @[NV_NVDLA_CSC_dl.scala 810:29:@20696.4]
  reg [31:0] _RAND_134;
  reg [511:0] _T_2074; // @[NV_NVDLA_CSC_dl.scala 815:19:@20700.4]
  reg [511:0] _RAND_135;
  reg [511:0] _T_2082; // @[NV_NVDLA_CSC_dl.scala 819:19:@20704.4]
  reg [511:0] _RAND_136;
  wire  _T_2105; // @[NV_NVDLA_CSC_dl.scala 831:69:@20719.4]
  wire  _T_2106; // @[NV_NVDLA_CSC_dl.scala 831:74:@20720.4]
  wire  _T_2107; // @[NV_NVDLA_CSC_dl.scala 831:90:@20721.4]
  wire  _T_2108; // @[NV_NVDLA_CSC_dl.scala 831:88:@20722.4]
  wire  _T_2148; // @[NV_NVDLA_CSC_dl.scala 846:22:@20756.4]
  wire  _T_2162; // @[NV_NVDLA_CSC_dl.scala 850:48:@20767.4]
  wire  _T_2163; // @[NV_NVDLA_CSC_dl.scala 850:22:@20768.4]
  reg [7:0] _T_2182; // @[NV_NVDLA_CSC_dl.scala 867:29:@20809.4]
  reg [31:0] _RAND_137;
  reg [7:0] _T_2185; // @[NV_NVDLA_CSC_dl.scala 868:29:@20810.4]
  reg [31:0] _RAND_138;
  reg [7:0] _T_2188; // @[NV_NVDLA_CSC_dl.scala 869:29:@20811.4]
  reg [31:0] _RAND_139;
  reg [7:0] _T_2191; // @[NV_NVDLA_CSC_dl.scala 870:29:@20812.4]
  reg [31:0] _RAND_140;
  reg [7:0] _T_2194; // @[NV_NVDLA_CSC_dl.scala 871:33:@20813.4]
  reg [31:0] _RAND_141;
  reg [7:0] _T_2197; // @[NV_NVDLA_CSC_dl.scala 872:33:@20814.4]
  reg [31:0] _RAND_142;
  reg [7:0] _T_2200; // @[NV_NVDLA_CSC_dl.scala 873:33:@20815.4]
  reg [31:0] _RAND_143;
  reg [7:0] _T_2203; // @[NV_NVDLA_CSC_dl.scala 874:33:@20816.4]
  reg [31:0] _RAND_144;
  reg  _T_2214; // @[NV_NVDLA_CSC_dl.scala 879:41:@20820.4]
  reg [31:0] _RAND_145;
  reg [26:0] _T_2228; // @[NV_NVDLA_CSC_dl.scala 881:41:@20825.4]
  reg [31:0] _RAND_146;
  wire [26:0] _T_2240; // @[Cat.scala 30:58:@20835.4]
  wire [26:0] _GEN_137; // @[NV_NVDLA_CSC_dl.scala 889:28:@20838.4]
  wire [26:0] _GEN_138; // @[NV_NVDLA_CSC_dl.scala 889:28:@20842.4]
  wire [26:0] _GEN_139; // @[NV_NVDLA_CSC_dl.scala 889:28:@20846.4]
  wire [26:0] _GEN_140; // @[NV_NVDLA_CSC_dl.scala 889:28:@20850.4]
  wire  _T_2269; // @[NV_NVDLA_CSC_dl.scala 907:39:@20876.4]
  wire  _T_2270; // @[NV_NVDLA_CSC_dl.scala 908:39:@20877.4]
  wire  _T_2271; // @[NV_NVDLA_CSC_dl.scala 909:39:@20878.4]
  wire  _T_2272; // @[NV_NVDLA_CSC_dl.scala 910:39:@20879.4]
  wire [8:0] _T_2273; // @[NV_NVDLA_CSC_dl.scala 912:38:@20880.4]
  wire [8:0] _T_2274; // @[NV_NVDLA_CSC_dl.scala 913:38:@20881.4]
  wire [8:0] _T_2275; // @[NV_NVDLA_CSC_dl.scala 914:38:@20882.4]
  wire [8:0] _T_2276; // @[NV_NVDLA_CSC_dl.scala 915:38:@20883.4]
  wire  _T_2277; // @[NV_NVDLA_CSC_dl.scala 917:44:@20884.4]
  wire  _T_2278; // @[NV_NVDLA_CSC_dl.scala 918:44:@20885.4]
  wire  _T_2279; // @[NV_NVDLA_CSC_dl.scala 919:44:@20886.4]
  wire  _T_2280; // @[NV_NVDLA_CSC_dl.scala 920:44:@20887.4]
  wire [1:0] _T_2281; // @[NV_NVDLA_CSC_dl.scala 923:31:@20888.4]
  wire [7:0] _T_2285; // @[NV_NVDLA_CSC_dl.scala 927:31:@20892.4]
  wire [1:0] _T_2286; // @[NV_NVDLA_CSC_dl.scala 928:35:@20893.4]
  wire [7:0] _T_2296; // @[NV_NVDLA_CSC_dl.scala 939:29:@20902.4]
  wire  _T_2307; // @[NV_NVDLA_CSC_dl.scala 944:50:@20906.4]
  wire [7:0] _GEN_713; // @[NV_NVDLA_CSC_dl.scala 944:111:@20907.4]
  wire [8:0] _T_2309; // @[NV_NVDLA_CSC_dl.scala 944:111:@20907.4]
  wire [7:0] _T_2310; // @[NV_NVDLA_CSC_dl.scala 944:111:@20908.4]
  wire [8:0] _T_2311; // @[NV_NVDLA_CSC_dl.scala 944:133:@20909.4]
  wire [8:0] _T_2312; // @[NV_NVDLA_CSC_dl.scala 944:133:@20910.4]
  wire [7:0] _T_2313; // @[NV_NVDLA_CSC_dl.scala 944:133:@20911.4]
  wire [7:0] _T_2314; // @[NV_NVDLA_CSC_dl.scala 944:29:@20912.4]
  wire [8:0] _T_2318; // @[NV_NVDLA_CSC_dl.scala 945:111:@20914.4]
  wire [7:0] _T_2319; // @[NV_NVDLA_CSC_dl.scala 945:111:@20915.4]
  wire [8:0] _T_2320; // @[NV_NVDLA_CSC_dl.scala 945:133:@20916.4]
  wire [8:0] _T_2321; // @[NV_NVDLA_CSC_dl.scala 945:133:@20917.4]
  wire [7:0] _T_2322; // @[NV_NVDLA_CSC_dl.scala 945:133:@20918.4]
  wire [7:0] _T_2323; // @[NV_NVDLA_CSC_dl.scala 945:29:@20919.4]
  wire [8:0] _T_2327; // @[NV_NVDLA_CSC_dl.scala 946:111:@20921.4]
  wire [7:0] _T_2328; // @[NV_NVDLA_CSC_dl.scala 946:111:@20922.4]
  wire [8:0] _T_2329; // @[NV_NVDLA_CSC_dl.scala 946:133:@20923.4]
  wire [8:0] _T_2330; // @[NV_NVDLA_CSC_dl.scala 946:133:@20924.4]
  wire [7:0] _T_2331; // @[NV_NVDLA_CSC_dl.scala 946:133:@20925.4]
  wire [7:0] _T_2332; // @[NV_NVDLA_CSC_dl.scala 946:29:@20926.4]
  wire [8:0] _T_2336; // @[NV_NVDLA_CSC_dl.scala 947:111:@20928.4]
  wire [7:0] _T_2337; // @[NV_NVDLA_CSC_dl.scala 947:111:@20929.4]
  wire [8:0] _T_2338; // @[NV_NVDLA_CSC_dl.scala 947:133:@20930.4]
  wire [8:0] _T_2339; // @[NV_NVDLA_CSC_dl.scala 947:133:@20931.4]
  wire [7:0] _T_2340; // @[NV_NVDLA_CSC_dl.scala 947:133:@20932.4]
  wire [7:0] _T_2341; // @[NV_NVDLA_CSC_dl.scala 947:29:@20933.4]
  wire  _T_2343; // @[NV_NVDLA_CSC_dl.scala 956:52:@20934.4]
  wire  _T_2344; // @[NV_NVDLA_CSC_dl.scala 956:50:@20935.4]
  wire  _T_2345; // @[NV_NVDLA_CSC_dl.scala 957:50:@20936.4]
  wire [7:0] _T_2350; // @[NV_NVDLA_CSC_dl.scala 957:27:@20939.4]
  wire [7:0] _T_2351; // @[NV_NVDLA_CSC_dl.scala 956:27:@20940.4]
  wire [7:0] _T_2352; // @[NV_NVDLA_CSC_dl.scala 955:27:@20941.4]
  wire  _T_2354; // @[NV_NVDLA_CSC_dl.scala 961:52:@20942.4]
  wire  _T_2355; // @[NV_NVDLA_CSC_dl.scala 961:50:@20943.4]
  wire  _T_2356; // @[NV_NVDLA_CSC_dl.scala 962:50:@20944.4]
  wire [7:0] _T_2361; // @[NV_NVDLA_CSC_dl.scala 962:27:@20947.4]
  wire [7:0] _T_2362; // @[NV_NVDLA_CSC_dl.scala 961:27:@20948.4]
  wire [7:0] _T_2363; // @[NV_NVDLA_CSC_dl.scala 960:27:@20949.4]
  wire  _T_2365; // @[NV_NVDLA_CSC_dl.scala 966:52:@20950.4]
  wire  _T_2366; // @[NV_NVDLA_CSC_dl.scala 966:50:@20951.4]
  wire  _T_2367; // @[NV_NVDLA_CSC_dl.scala 967:50:@20952.4]
  wire [7:0] _T_2372; // @[NV_NVDLA_CSC_dl.scala 967:27:@20955.4]
  wire [7:0] _T_2373; // @[NV_NVDLA_CSC_dl.scala 966:27:@20956.4]
  wire [7:0] _T_2374; // @[NV_NVDLA_CSC_dl.scala 965:27:@20957.4]
  wire  _T_2376; // @[NV_NVDLA_CSC_dl.scala 971:52:@20958.4]
  wire  _T_2377; // @[NV_NVDLA_CSC_dl.scala 971:50:@20959.4]
  wire  _T_2378; // @[NV_NVDLA_CSC_dl.scala 972:50:@20960.4]
  wire [7:0] _T_2383; // @[NV_NVDLA_CSC_dl.scala 972:27:@20963.4]
  wire [7:0] _T_2384; // @[NV_NVDLA_CSC_dl.scala 971:27:@20964.4]
  wire [7:0] _T_2385; // @[NV_NVDLA_CSC_dl.scala 970:27:@20965.4]
  wire  _T_2386; // @[NV_NVDLA_CSC_dl.scala 976:46:@20966.4]
  wire  _T_2387; // @[NV_NVDLA_CSC_dl.scala 976:51:@20967.4]
  wire  _T_2388; // @[NV_NVDLA_CSC_dl.scala 976:34:@20968.4]
  wire  _T_2389; // @[NV_NVDLA_CSC_dl.scala 977:46:@20969.4]
  wire  _T_2390; // @[NV_NVDLA_CSC_dl.scala 977:51:@20970.4]
  wire  _T_2392; // @[NV_NVDLA_CSC_dl.scala 977:87:@20971.4]
  wire  _T_2393; // @[NV_NVDLA_CSC_dl.scala 977:69:@20972.4]
  wire  _T_2394; // @[NV_NVDLA_CSC_dl.scala 977:34:@20973.4]
  wire  _T_2395; // @[NV_NVDLA_CSC_dl.scala 978:46:@20974.4]
  wire  _T_2396; // @[NV_NVDLA_CSC_dl.scala 978:51:@20975.4]
  wire  _T_2398; // @[NV_NVDLA_CSC_dl.scala 978:87:@20976.4]
  wire  _T_2399; // @[NV_NVDLA_CSC_dl.scala 978:69:@20977.4]
  wire  _T_2400; // @[NV_NVDLA_CSC_dl.scala 978:34:@20978.4]
  wire  _T_2401; // @[NV_NVDLA_CSC_dl.scala 979:46:@20979.4]
  wire  _T_2402; // @[NV_NVDLA_CSC_dl.scala 979:51:@20980.4]
  wire  _T_2405; // @[NV_NVDLA_CSC_dl.scala 979:69:@20982.4]
  wire  _T_2406; // @[NV_NVDLA_CSC_dl.scala 979:34:@20983.4]
  wire  _T_2407; // @[NV_NVDLA_CSC_dl.scala 981:50:@20984.4]
  wire  _T_2408; // @[NV_NVDLA_CSC_dl.scala 981:55:@20985.4]
  wire  _T_2409; // @[NV_NVDLA_CSC_dl.scala 981:73:@20986.4]
  wire  _T_2410; // @[NV_NVDLA_CSC_dl.scala 981:97:@20987.4]
  wire  _T_2411; // @[NV_NVDLA_CSC_dl.scala 981:38:@20988.4]
  wire  _T_2412; // @[NV_NVDLA_CSC_dl.scala 982:50:@20989.4]
  wire  _T_2413; // @[NV_NVDLA_CSC_dl.scala 982:55:@20990.4]
  wire  _T_2414; // @[NV_NVDLA_CSC_dl.scala 982:73:@20991.4]
  wire  _T_2415; // @[NV_NVDLA_CSC_dl.scala 982:97:@20992.4]
  wire  _T_2417; // @[NV_NVDLA_CSC_dl.scala 982:138:@20993.4]
  wire  _T_2418; // @[NV_NVDLA_CSC_dl.scala 982:120:@20994.4]
  wire  _T_2419; // @[NV_NVDLA_CSC_dl.scala 982:38:@20995.4]
  wire  _T_2420; // @[NV_NVDLA_CSC_dl.scala 983:50:@20996.4]
  wire  _T_2421; // @[NV_NVDLA_CSC_dl.scala 983:55:@20997.4]
  wire  _T_2422; // @[NV_NVDLA_CSC_dl.scala 983:73:@20998.4]
  wire  _T_2423; // @[NV_NVDLA_CSC_dl.scala 983:97:@20999.4]
  wire  _T_2425; // @[NV_NVDLA_CSC_dl.scala 983:138:@21000.4]
  wire  _T_2426; // @[NV_NVDLA_CSC_dl.scala 983:120:@21001.4]
  wire  _T_2427; // @[NV_NVDLA_CSC_dl.scala 983:38:@21002.4]
  wire  _T_2428; // @[NV_NVDLA_CSC_dl.scala 984:50:@21003.4]
  wire  _T_2429; // @[NV_NVDLA_CSC_dl.scala 984:55:@21004.4]
  wire  _T_2430; // @[NV_NVDLA_CSC_dl.scala 984:73:@21005.4]
  wire  _T_2431; // @[NV_NVDLA_CSC_dl.scala 984:97:@21006.4]
  wire  _T_2434; // @[NV_NVDLA_CSC_dl.scala 984:120:@21008.4]
  wire  _T_2435; // @[NV_NVDLA_CSC_dl.scala 984:38:@21009.4]
  wire [7:0] _GEN_141; // @[NV_NVDLA_CSC_dl.scala 986:24:@21010.4]
  wire [7:0] _GEN_142; // @[NV_NVDLA_CSC_dl.scala 987:24:@21013.4]
  wire [7:0] _GEN_143; // @[NV_NVDLA_CSC_dl.scala 988:24:@21016.4]
  wire [7:0] _GEN_144; // @[NV_NVDLA_CSC_dl.scala 989:24:@21019.4]
  wire [7:0] _GEN_145; // @[NV_NVDLA_CSC_dl.scala 990:28:@21022.4]
  wire [7:0] _GEN_146; // @[NV_NVDLA_CSC_dl.scala 991:28:@21025.4]
  wire [7:0] _GEN_147; // @[NV_NVDLA_CSC_dl.scala 992:28:@21028.4]
  wire [7:0] _GEN_148; // @[NV_NVDLA_CSC_dl.scala 993:28:@21031.4]
  wire [7:0] _T_2436; // @[NV_NVDLA_CSC_dl.scala 1002:55:@21034.4]
  wire [63:0] _T_2439; // @[Cat.scala 30:58:@21037.4]
  wire [127:0] _T_2440; // @[Cat.scala 30:58:@21038.4]
  wire [255:0] _T_2441; // @[Cat.scala 30:58:@21039.4]
  wire [511:0] _T_2442; // @[Cat.scala 30:58:@21040.4]
  wire [511:0] _T_2443; // @[NV_NVDLA_CSC_dl.scala 1004:23:@21041.4]
  wire [511:0] _T_2447; // @[NV_NVDLA_CSC_dl.scala 1009:23:@21045.4]
  wire  _T_2453; // @[NV_NVDLA_CSC_dl.scala 1022:37:@21050.4]
  wire  _T_2456; // @[NV_NVDLA_CSC_dl.scala 1023:43:@21051.4]
  wire  _T_2457; // @[NV_NVDLA_CSC_dl.scala 1023:87:@21052.4]
  wire  _T_2459; // @[NV_NVDLA_CSC_dl.scala 1023:91:@21053.4]
  wire  _T_2460; // @[NV_NVDLA_CSC_dl.scala 1023:72:@21054.4]
  wire [255:0] _T_2462; // @[NV_NVDLA_CSC_dl.scala 1023:171:@21055.4]
  wire [511:0] _T_2463; // @[Cat.scala 30:58:@21056.4]
  wire  _T_2469; // @[NV_NVDLA_CSC_dl.scala 1024:72:@21060.4]
  wire [255:0] _T_2471; // @[NV_NVDLA_CSC_dl.scala 1024:171:@21061.4]
  wire [511:0] _T_2472; // @[Cat.scala 30:58:@21062.4]
  wire [511:0] _T_2473; // @[NV_NVDLA_CSC_dl.scala 1024:27:@21063.4]
  wire [511:0] _T_2474; // @[NV_NVDLA_CSC_dl.scala 1023:27:@21064.4]
  wire [511:0] _T_2475; // @[NV_NVDLA_CSC_dl.scala 1022:27:@21065.4]
  wire [7:0] _T_2546; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21068.4]
  wire [7:0] _T_2547; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21070.4]
  wire [7:0] _T_2548; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21072.4]
  wire [7:0] _T_2549; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21074.4]
  wire [7:0] _T_2550; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21076.4]
  wire [7:0] _T_2551; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21078.4]
  wire [7:0] _T_2552; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21080.4]
  wire [7:0] _T_2553; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21082.4]
  wire [7:0] _T_2554; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21084.4]
  wire [7:0] _T_2555; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21086.4]
  wire [7:0] _T_2556; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21088.4]
  wire [7:0] _T_2557; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21090.4]
  wire [7:0] _T_2558; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21092.4]
  wire [7:0] _T_2559; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21094.4]
  wire [7:0] _T_2560; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21096.4]
  wire [7:0] _T_2561; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21098.4]
  wire [7:0] _T_2562; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21100.4]
  wire [7:0] _T_2563; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21102.4]
  wire [7:0] _T_2564; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21104.4]
  wire [7:0] _T_2565; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21106.4]
  wire [7:0] _T_2566; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21108.4]
  wire [7:0] _T_2567; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21110.4]
  wire [7:0] _T_2568; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21112.4]
  wire [7:0] _T_2569; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21114.4]
  wire [7:0] _T_2570; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21116.4]
  wire [7:0] _T_2571; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21118.4]
  wire [7:0] _T_2572; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21120.4]
  wire [7:0] _T_2573; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21122.4]
  wire [7:0] _T_2574; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21124.4]
  wire [7:0] _T_2575; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21126.4]
  wire [7:0] _T_2576; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21128.4]
  wire [7:0] _T_2577; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21130.4]
  wire [7:0] _T_2578; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21132.4]
  wire [7:0] _T_2579; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21134.4]
  wire [7:0] _T_2580; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21136.4]
  wire [7:0] _T_2581; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21138.4]
  wire [7:0] _T_2582; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21140.4]
  wire [7:0] _T_2583; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21142.4]
  wire [7:0] _T_2584; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21144.4]
  wire [7:0] _T_2585; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21146.4]
  wire [7:0] _T_2586; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21148.4]
  wire [7:0] _T_2587; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21150.4]
  wire [7:0] _T_2588; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21152.4]
  wire [7:0] _T_2589; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21154.4]
  wire [7:0] _T_2590; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21156.4]
  wire [7:0] _T_2591; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21158.4]
  wire [7:0] _T_2592; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21160.4]
  wire [7:0] _T_2593; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21162.4]
  wire [7:0] _T_2594; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21164.4]
  wire [7:0] _T_2595; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21166.4]
  wire [7:0] _T_2596; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21168.4]
  wire [7:0] _T_2597; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21170.4]
  wire [7:0] _T_2598; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21172.4]
  wire [7:0] _T_2599; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21174.4]
  wire [7:0] _T_2600; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21176.4]
  wire [7:0] _T_2601; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21178.4]
  wire [7:0] _T_2602; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21180.4]
  wire [7:0] _T_2603; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21182.4]
  wire [7:0] _T_2604; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21184.4]
  wire [7:0] _T_2605; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21186.4]
  wire [7:0] _T_2606; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21188.4]
  wire [7:0] _T_2607; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21190.4]
  wire [7:0] _T_2608; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21192.4]
  wire [7:0] _T_2609; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21194.4]
  reg [255:0] _T_2611; // @[NV_NVDLA_CSC_dl.scala 1044:28:@21196.4]
  reg [255:0] _RAND_147;
  reg [127:0] _T_2613; // @[NV_NVDLA_CSC_dl.scala 1045:28:@21197.4]
  reg [127:0] _RAND_148;
  reg [127:0] _T_2615; // @[NV_NVDLA_CSC_dl.scala 1046:28:@21198.4]
  reg [127:0] _RAND_149;
  reg [127:0] _T_2617; // @[NV_NVDLA_CSC_dl.scala 1048:28:@21199.4]
  reg [127:0] _RAND_150;
  reg [127:0] _T_2619; // @[NV_NVDLA_CSC_dl.scala 1049:28:@21200.4]
  reg [127:0] _RAND_151;
  reg [127:0] _T_2621; // @[NV_NVDLA_CSC_dl.scala 1051:28:@21201.4]
  reg [127:0] _RAND_152;
  wire  _T_2622; // @[NV_NVDLA_CSC_dl.scala 1053:39:@21202.4]
  wire  _T_2623; // @[NV_NVDLA_CSC_dl.scala 1053:29:@21203.4]
  wire [1023:0] _T_2625; // @[Cat.scala 30:58:@21204.4]
  wire [1023:0] _T_2626; // @[NV_NVDLA_CSC_dl.scala 1053:28:@21205.4]
  wire  _T_2627; // @[NV_NVDLA_CSC_dl.scala 1054:39:@21206.4]
  wire  _T_2628; // @[NV_NVDLA_CSC_dl.scala 1054:29:@21207.4]
  wire [1023:0] _T_2630; // @[Cat.scala 30:58:@21208.4]
  wire [1023:0] _T_2631; // @[NV_NVDLA_CSC_dl.scala 1054:28:@21209.4]
  wire  _T_2632; // @[NV_NVDLA_CSC_dl.scala 1055:39:@21210.4]
  wire  _T_2633; // @[NV_NVDLA_CSC_dl.scala 1055:29:@21211.4]
  wire [1023:0] _T_2636; // @[NV_NVDLA_CSC_dl.scala 1055:28:@21213.4]
  wire  _T_2637; // @[NV_NVDLA_CSC_dl.scala 1056:39:@21214.4]
  wire  _T_2638; // @[NV_NVDLA_CSC_dl.scala 1056:29:@21215.4]
  wire [1023:0] _T_2641; // @[NV_NVDLA_CSC_dl.scala 1056:28:@21217.4]
  wire [10:0] _T_2643; // @[Cat.scala 30:58:@21218.4]
  wire [1023:0] _T_2644; // @[NV_NVDLA_CSC_dl.scala 1058:41:@21219.4]
  wire [511:0] _T_2645; // @[NV_NVDLA_CSC_dl.scala 1058:82:@21220.4]
  wire [10:0] _T_2647; // @[Cat.scala 30:58:@21221.4]
  wire [1023:0] _T_2648; // @[NV_NVDLA_CSC_dl.scala 1059:41:@21222.4]
  wire [511:0] _T_2649; // @[NV_NVDLA_CSC_dl.scala 1059:82:@21223.4]
  wire [10:0] _T_2651; // @[Cat.scala 30:58:@21224.4]
  wire [1023:0] _T_2652; // @[NV_NVDLA_CSC_dl.scala 1060:41:@21225.4]
  wire [511:0] _T_2653; // @[NV_NVDLA_CSC_dl.scala 1060:82:@21226.4]
  wire [10:0] _T_2655; // @[Cat.scala 30:58:@21227.4]
  wire [1023:0] _T_2656; // @[NV_NVDLA_CSC_dl.scala 1061:41:@21228.4]
  wire [511:0] _T_2657; // @[NV_NVDLA_CSC_dl.scala 1061:82:@21229.4]
  wire  _T_2658; // @[NV_NVDLA_CSC_dl.scala 1063:36:@21230.4]
  wire  _T_2659; // @[NV_NVDLA_CSC_dl.scala 1063:26:@21231.4]
  wire  _T_2662; // @[NV_NVDLA_CSC_dl.scala 1064:41:@21232.4]
  wire [127:0] _T_2663; // @[NV_NVDLA_CSC_dl.scala 1064:81:@21233.4]
  wire [511:0] _T_2669; // @[Cat.scala 30:58:@21239.4]
  wire  _T_2671; // @[NV_NVDLA_CSC_dl.scala 1065:41:@21240.4]
  wire [255:0] _T_2672; // @[NV_NVDLA_CSC_dl.scala 1065:81:@21241.4]
  wire [511:0] _T_2674; // @[Cat.scala 30:58:@21243.4]
  wire [511:0] _T_2676; // @[NV_NVDLA_CSC_dl.scala 1065:25:@21245.4]
  wire [511:0] _T_2677; // @[NV_NVDLA_CSC_dl.scala 1064:25:@21246.4]
  wire [511:0] _T_2678; // @[NV_NVDLA_CSC_dl.scala 1063:25:@21247.4]
  wire [7:0] _T_2749; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21249.4]
  wire [7:0] _T_2750; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21251.4]
  wire [7:0] _T_2751; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21253.4]
  wire [7:0] _T_2752; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21255.4]
  wire [7:0] _T_2753; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21257.4]
  wire [7:0] _T_2754; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21259.4]
  wire [7:0] _T_2755; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21261.4]
  wire [7:0] _T_2756; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21263.4]
  wire [7:0] _T_2757; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21265.4]
  wire [7:0] _T_2758; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21267.4]
  wire [7:0] _T_2759; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21269.4]
  wire [7:0] _T_2760; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21271.4]
  wire [7:0] _T_2761; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21273.4]
  wire [7:0] _T_2762; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21275.4]
  wire [7:0] _T_2763; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21277.4]
  wire [7:0] _T_2764; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21279.4]
  wire [7:0] _T_2765; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21281.4]
  wire [7:0] _T_2766; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21283.4]
  wire [7:0] _T_2767; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21285.4]
  wire [7:0] _T_2768; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21287.4]
  wire [7:0] _T_2769; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21289.4]
  wire [7:0] _T_2770; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21291.4]
  wire [7:0] _T_2771; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21293.4]
  wire [7:0] _T_2772; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21295.4]
  wire [7:0] _T_2773; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21297.4]
  wire [7:0] _T_2774; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21299.4]
  wire [7:0] _T_2775; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21301.4]
  wire [7:0] _T_2776; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21303.4]
  wire [7:0] _T_2777; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21305.4]
  wire [7:0] _T_2778; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21307.4]
  wire [7:0] _T_2779; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21309.4]
  wire [7:0] _T_2780; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21311.4]
  wire [7:0] _T_2781; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21313.4]
  wire [7:0] _T_2782; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21315.4]
  wire [7:0] _T_2783; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21317.4]
  wire [7:0] _T_2784; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21319.4]
  wire [7:0] _T_2785; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21321.4]
  wire [7:0] _T_2786; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21323.4]
  wire [7:0] _T_2787; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21325.4]
  wire [7:0] _T_2788; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21327.4]
  wire [7:0] _T_2789; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21329.4]
  wire [7:0] _T_2790; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21331.4]
  wire [7:0] _T_2791; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21333.4]
  wire [7:0] _T_2792; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21335.4]
  wire [7:0] _T_2793; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21337.4]
  wire [7:0] _T_2794; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21339.4]
  wire [7:0] _T_2795; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21341.4]
  wire [7:0] _T_2796; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21343.4]
  wire [7:0] _T_2797; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21345.4]
  wire [7:0] _T_2798; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21347.4]
  wire [7:0] _T_2799; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21349.4]
  wire [7:0] _T_2800; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21351.4]
  wire [7:0] _T_2801; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21353.4]
  wire [7:0] _T_2802; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21355.4]
  wire [7:0] _T_2803; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21357.4]
  wire [7:0] _T_2804; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21359.4]
  wire [7:0] _T_2805; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21361.4]
  wire [7:0] _T_2806; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21363.4]
  wire [7:0] _T_2807; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21365.4]
  wire [7:0] _T_2808; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21367.4]
  wire [7:0] _T_2809; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21369.4]
  wire [7:0] _T_2810; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21371.4]
  wire [7:0] _T_2811; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21373.4]
  wire [7:0] _T_2812; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21375.4]
  wire  _T_2814; // @[NV_NVDLA_CSC_dl.scala 1074:59:@21377.4]
  wire  _T_2815; // @[NV_NVDLA_CSC_dl.scala 1074:41:@21378.4]
  wire  _T_2817; // @[NV_NVDLA_CSC_dl.scala 1075:59:@21379.4]
  wire  _T_2818; // @[NV_NVDLA_CSC_dl.scala 1075:41:@21380.4]
  wire  _T_2821; // @[NV_NVDLA_CSC_dl.scala 1076:41:@21382.4]
  wire [511:0] _GEN_149; // @[NV_NVDLA_CSC_dl.scala 1078:24:@21383.4]
  wire [255:0] _GEN_150; // @[NV_NVDLA_CSC_dl.scala 1081:24:@21386.4]
  wire [511:0] _GEN_151; // @[NV_NVDLA_CSC_dl.scala 1081:24:@21386.4]
  wire [511:0] _GEN_154; // @[NV_NVDLA_CSC_dl.scala 1085:24:@21390.4]
  wire [318:0] _T_2827; // @[NV_NVDLA_CSC_dl.scala 1094:56:@21396.4]
  wire [63:0] _T_2828; // @[NV_NVDLA_CSC_dl.scala 1094:73:@21397.4]
  wire [63:0] _T_2829; // @[NV_NVDLA_CSC_dl.scala 1094:24:@21398.4]
  wire  _T_2831; // @[NV_NVDLA_CSC_dl.scala 1096:51:@21399.4]
  wire [63:0] _T_2838; // @[NV_NVDLA_CSC_dl.scala 1096:32:@21401.4]
  wire  _T_2840; // @[NV_NVDLA_CSC_dl.scala 1097:51:@21402.4]
  wire [31:0] _T_2847; // @[NV_NVDLA_CSC_dl.scala 1097:32:@21404.4]
  wire  _T_2849; // @[NV_NVDLA_CSC_dl.scala 1098:51:@21405.4]
  wire [31:0] _T_2856; // @[NV_NVDLA_CSC_dl.scala 1098:32:@21407.4]
  wire [31:0] _T_2857; // @[NV_NVDLA_CSC_dl.scala 1100:57:@21408.4]
  wire [63:0] _T_2863; // @[Cat.scala 30:58:@21410.4]
  wire [15:0] _T_2864; // @[NV_NVDLA_CSC_dl.scala 1101:57:@21411.4]
  wire [15:0] _T_2865; // @[NV_NVDLA_CSC_dl.scala 1101:106:@21412.4]
  wire [15:0] _T_2866; // @[NV_NVDLA_CSC_dl.scala 1101:155:@21413.4]
  wire [63:0] _T_2874; // @[Cat.scala 30:58:@21417.4]
  wire  _T_2876; // @[NV_NVDLA_CSC_dl.scala 1103:43:@21418.4]
  wire [15:0] _T_2877; // @[NV_NVDLA_CSC_dl.scala 1103:89:@21419.4]
  wire [63:0] _T_2879; // @[Cat.scala 30:58:@21421.4]
  wire [63:0] _T_2880; // @[NV_NVDLA_CSC_dl.scala 1103:116:@21422.4]
  wire  _T_2882; // @[NV_NVDLA_CSC_dl.scala 1104:43:@21423.4]
  wire [31:0] _T_2883; // @[NV_NVDLA_CSC_dl.scala 1104:89:@21424.4]
  wire [63:0] _T_2884; // @[Cat.scala 30:58:@21425.4]
  wire [63:0] _T_2885; // @[NV_NVDLA_CSC_dl.scala 1104:116:@21426.4]
  wire [63:0] _T_2886; // @[NV_NVDLA_CSC_dl.scala 1104:26:@21427.4]
  wire [63:0] _T_2887; // @[NV_NVDLA_CSC_dl.scala 1103:26:@21428.4]
  wire  _T_2888; // @[NV_NVDLA_CSC_dl.scala 1108:35:@21429.4]
  wire [7:0] _T_2889_0; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_1; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_2; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_3; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_4; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_5; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_6; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_7; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_8; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_9; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_10; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_11; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_12; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_13; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_14; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_15; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_16; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_17; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_18; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_19; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_20; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_21; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_22; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_23; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_24; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_25; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_26; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_27; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_28; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_29; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_30; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_31; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_32; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_33; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_34; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_35; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_36; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_37; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_38; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_39; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_40; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_41; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_42; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_43; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_44; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_45; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_46; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_47; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_48; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_49; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_50; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_51; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_52; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_53; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_54; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_55; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_56; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_57; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_58; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_59; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_60; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_61; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_62; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire [7:0] _T_2889_63; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  wire  _T_3022; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21431.4]
  wire  _T_3024; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21432.4]
  wire  _T_3026; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21433.4]
  wire  _T_3028; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21434.4]
  wire  _T_3030; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21435.4]
  wire  _T_3032; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21436.4]
  wire  _T_3034; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21437.4]
  wire  _T_3036; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21438.4]
  wire  _T_3038; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21439.4]
  wire  _T_3040; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21440.4]
  wire  _T_3042; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21441.4]
  wire  _T_3044; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21442.4]
  wire  _T_3046; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21443.4]
  wire  _T_3048; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21444.4]
  wire  _T_3050; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21445.4]
  wire  _T_3052; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21446.4]
  wire  _T_3054; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21447.4]
  wire  _T_3056; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21448.4]
  wire  _T_3058; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21449.4]
  wire  _T_3060; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21450.4]
  wire  _T_3062; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21451.4]
  wire  _T_3064; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21452.4]
  wire  _T_3066; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21453.4]
  wire  _T_3068; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21454.4]
  wire  _T_3070; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21455.4]
  wire  _T_3072; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21456.4]
  wire  _T_3074; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21457.4]
  wire  _T_3076; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21458.4]
  wire  _T_3078; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21459.4]
  wire  _T_3080; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21460.4]
  wire  _T_3082; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21461.4]
  wire  _T_3084; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21462.4]
  wire  _T_3086; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21463.4]
  wire  _T_3088; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21464.4]
  wire  _T_3090; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21465.4]
  wire  _T_3092; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21466.4]
  wire  _T_3094; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21467.4]
  wire  _T_3096; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21468.4]
  wire  _T_3098; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21469.4]
  wire  _T_3100; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21470.4]
  wire  _T_3102; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21471.4]
  wire  _T_3104; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21472.4]
  wire  _T_3106; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21473.4]
  wire  _T_3108; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21474.4]
  wire  _T_3110; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21475.4]
  wire  _T_3112; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21476.4]
  wire  _T_3114; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21477.4]
  wire  _T_3116; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21478.4]
  wire  _T_3118; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21479.4]
  wire  _T_3120; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21480.4]
  wire  _T_3122; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21481.4]
  wire  _T_3124; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21482.4]
  wire  _T_3126; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21483.4]
  wire  _T_3128; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21484.4]
  wire  _T_3130; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21485.4]
  wire  _T_3132; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21486.4]
  wire  _T_3134; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21487.4]
  wire  _T_3136; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21488.4]
  wire  _T_3138; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21489.4]
  wire  _T_3140; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21490.4]
  wire  _T_3142; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21491.4]
  wire  _T_3144; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21492.4]
  wire  _T_3146; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21493.4]
  wire  _T_3148; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21494.4]
  wire  _T_3219; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21560.4]
  wire  _T_3220; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21561.4]
  wire  _T_3221; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21562.4]
  wire  _T_3222; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21563.4]
  wire  _T_3223; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21564.4]
  wire  _T_3224; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21565.4]
  wire  _T_3225; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21566.4]
  wire  _T_3226; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21567.4]
  wire  _T_3227; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21568.4]
  wire  _T_3228; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21569.4]
  wire  _T_3229; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21570.4]
  wire  _T_3230; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21571.4]
  wire  _T_3231; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21572.4]
  wire  _T_3232; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21573.4]
  wire  _T_3233; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21574.4]
  wire  _T_3234; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21575.4]
  wire  _T_3235; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21576.4]
  wire  _T_3236; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21577.4]
  wire  _T_3237; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21578.4]
  wire  _T_3238; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21579.4]
  wire  _T_3239; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21580.4]
  wire  _T_3240; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21581.4]
  wire  _T_3241; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21582.4]
  wire  _T_3242; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21583.4]
  wire  _T_3243; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21584.4]
  wire  _T_3244; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21585.4]
  wire  _T_3245; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21586.4]
  wire  _T_3246; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21587.4]
  wire  _T_3247; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21588.4]
  wire  _T_3248; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21589.4]
  wire  _T_3249; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21590.4]
  wire  _T_3250; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21591.4]
  wire  _T_3251; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21592.4]
  wire  _T_3252; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21593.4]
  wire  _T_3253; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21594.4]
  wire  _T_3254; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21595.4]
  wire  _T_3255; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21596.4]
  wire  _T_3256; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21597.4]
  wire  _T_3257; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21598.4]
  wire  _T_3258; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21599.4]
  wire  _T_3259; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21600.4]
  wire  _T_3260; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21601.4]
  wire  _T_3261; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21602.4]
  wire  _T_3262; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21603.4]
  wire  _T_3263; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21604.4]
  wire  _T_3264; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21605.4]
  wire  _T_3265; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21606.4]
  wire  _T_3266; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21607.4]
  wire  _T_3267; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21608.4]
  wire  _T_3268; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21609.4]
  wire  _T_3269; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21610.4]
  wire  _T_3270; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21611.4]
  wire  _T_3271; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21612.4]
  wire  _T_3272; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21613.4]
  wire  _T_3273; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21614.4]
  wire  _T_3274; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21615.4]
  wire  _T_3275; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21616.4]
  wire  _T_3276; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21617.4]
  wire  _T_3277; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21618.4]
  wire  _T_3278; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21619.4]
  wire  _T_3279; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21620.4]
  wire  _T_3280; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21621.4]
  wire  _T_3281; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21622.4]
  wire  _T_3282; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21623.4]
  wire  _T_3283; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21624.4]
  wire  _T_3284; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21625.4]
  wire  _T_3285; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21626.4]
  wire  _T_3286; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21627.4]
  wire  _T_3287; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21628.4]
  wire  _T_3288; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21629.4]
  wire  _T_3289; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21630.4]
  wire  _T_3290; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21631.4]
  wire  _T_3291; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21632.4]
  wire  _T_3292; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21633.4]
  wire  _T_3293; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21634.4]
  wire  _T_3294; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21635.4]
  wire  _T_3295; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21636.4]
  wire  _T_3296; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21637.4]
  wire  _T_3297; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21638.4]
  wire  _T_3298; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21639.4]
  wire  _T_3299; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21640.4]
  wire  _T_3300; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21641.4]
  wire  _T_3301; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21642.4]
  wire  _T_3302; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21643.4]
  wire  _T_3303; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21644.4]
  wire  _T_3304; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21645.4]
  wire  _T_3305; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21646.4]
  wire  _T_3306; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21647.4]
  wire  _T_3307; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21648.4]
  wire  _T_3308; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21649.4]
  wire  _T_3309; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21650.4]
  wire  _T_3310; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21651.4]
  wire  _T_3311; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21652.4]
  wire  _T_3312; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21653.4]
  wire  _T_3313; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21654.4]
  wire  _T_3314; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21655.4]
  wire  _T_3315; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21656.4]
  wire  _T_3316; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21657.4]
  wire  _T_3317; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21658.4]
  wire  _T_3318; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21659.4]
  wire  _T_3319; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21660.4]
  wire  _T_3320; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21661.4]
  wire  _T_3321; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21662.4]
  wire  _T_3322; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21663.4]
  wire  _T_3323; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21664.4]
  wire  _T_3324; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21665.4]
  wire  _T_3325; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21666.4]
  wire  _T_3326; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21667.4]
  wire  _T_3327; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21668.4]
  wire  _T_3328; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21669.4]
  wire  _T_3329; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21670.4]
  wire  _T_3330; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21671.4]
  wire  _T_3331; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21672.4]
  wire  _T_3332; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21673.4]
  wire  _T_3333; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21674.4]
  wire  _T_3334; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21675.4]
  wire  _T_3335; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21676.4]
  wire  _T_3336; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21677.4]
  wire  _T_3337; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21678.4]
  wire  _T_3338; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21679.4]
  wire  _T_3339; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21680.4]
  wire  _T_3340; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21681.4]
  wire  _T_3341; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21682.4]
  wire  _T_3342; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21683.4]
  wire  _T_3343; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21684.4]
  wire  _T_3344; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21685.4]
  wire  _T_3345; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21686.4]
  wire  _T_3346; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21687.4]
  reg  _T_3419; // @[NV_NVDLA_CSC_dl.scala 1117:27:@21753.4]
  reg [31:0] _RAND_153;
  reg  _T_3689_0; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_154;
  reg  _T_3689_1; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_155;
  reg  _T_3689_2; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_156;
  reg  _T_3689_3; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_157;
  reg  _T_3689_4; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_158;
  reg  _T_3689_5; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_159;
  reg  _T_3689_6; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_160;
  reg  _T_3689_7; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_161;
  reg  _T_3689_8; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_162;
  reg  _T_3689_9; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_163;
  reg  _T_3689_10; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_164;
  reg  _T_3689_11; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_165;
  reg  _T_3689_12; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_166;
  reg  _T_3689_13; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_167;
  reg  _T_3689_14; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_168;
  reg  _T_3689_15; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_169;
  reg  _T_3689_16; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_170;
  reg  _T_3689_17; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_171;
  reg  _T_3689_18; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_172;
  reg  _T_3689_19; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_173;
  reg  _T_3689_20; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_174;
  reg  _T_3689_21; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_175;
  reg  _T_3689_22; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_176;
  reg  _T_3689_23; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_177;
  reg  _T_3689_24; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_178;
  reg  _T_3689_25; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_179;
  reg  _T_3689_26; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_180;
  reg  _T_3689_27; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_181;
  reg  _T_3689_28; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_182;
  reg  _T_3689_29; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_183;
  reg  _T_3689_30; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_184;
  reg  _T_3689_31; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_185;
  reg  _T_3689_32; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_186;
  reg  _T_3689_33; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_187;
  reg  _T_3689_34; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_188;
  reg  _T_3689_35; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_189;
  reg  _T_3689_36; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_190;
  reg  _T_3689_37; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_191;
  reg  _T_3689_38; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_192;
  reg  _T_3689_39; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_193;
  reg  _T_3689_40; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_194;
  reg  _T_3689_41; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_195;
  reg  _T_3689_42; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_196;
  reg  _T_3689_43; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_197;
  reg  _T_3689_44; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_198;
  reg  _T_3689_45; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_199;
  reg  _T_3689_46; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_200;
  reg  _T_3689_47; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_201;
  reg  _T_3689_48; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_202;
  reg  _T_3689_49; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_203;
  reg  _T_3689_50; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_204;
  reg  _T_3689_51; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_205;
  reg  _T_3689_52; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_206;
  reg  _T_3689_53; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_207;
  reg  _T_3689_54; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_208;
  reg  _T_3689_55; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_209;
  reg  _T_3689_56; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_210;
  reg  _T_3689_57; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_211;
  reg  _T_3689_58; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_212;
  reg  _T_3689_59; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_213;
  reg  _T_3689_60; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_214;
  reg  _T_3689_61; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_215;
  reg  _T_3689_62; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_216;
  reg  _T_3689_63; // @[NV_NVDLA_CSC_dl.scala 1119:34:@21820.4]
  reg [31:0] _RAND_217;
  reg [7:0] _T_3889_0; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_218;
  reg [7:0] _T_3889_1; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_219;
  reg [7:0] _T_3889_2; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_220;
  reg [7:0] _T_3889_3; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_221;
  reg [7:0] _T_3889_4; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_222;
  reg [7:0] _T_3889_5; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_223;
  reg [7:0] _T_3889_6; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_224;
  reg [7:0] _T_3889_7; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_225;
  reg [7:0] _T_3889_8; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_226;
  reg [7:0] _T_3889_9; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_227;
  reg [7:0] _T_3889_10; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_228;
  reg [7:0] _T_3889_11; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_229;
  reg [7:0] _T_3889_12; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_230;
  reg [7:0] _T_3889_13; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_231;
  reg [7:0] _T_3889_14; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_232;
  reg [7:0] _T_3889_15; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_233;
  reg [7:0] _T_3889_16; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_234;
  reg [7:0] _T_3889_17; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_235;
  reg [7:0] _T_3889_18; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_236;
  reg [7:0] _T_3889_19; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_237;
  reg [7:0] _T_3889_20; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_238;
  reg [7:0] _T_3889_21; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_239;
  reg [7:0] _T_3889_22; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_240;
  reg [7:0] _T_3889_23; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_241;
  reg [7:0] _T_3889_24; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_242;
  reg [7:0] _T_3889_25; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_243;
  reg [7:0] _T_3889_26; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_244;
  reg [7:0] _T_3889_27; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_245;
  reg [7:0] _T_3889_28; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_246;
  reg [7:0] _T_3889_29; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_247;
  reg [7:0] _T_3889_30; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_248;
  reg [7:0] _T_3889_31; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_249;
  reg [7:0] _T_3889_32; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_250;
  reg [7:0] _T_3889_33; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_251;
  reg [7:0] _T_3889_34; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_252;
  reg [7:0] _T_3889_35; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_253;
  reg [7:0] _T_3889_36; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_254;
  reg [7:0] _T_3889_37; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_255;
  reg [7:0] _T_3889_38; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_256;
  reg [7:0] _T_3889_39; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_257;
  reg [7:0] _T_3889_40; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_258;
  reg [7:0] _T_3889_41; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_259;
  reg [7:0] _T_3889_42; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_260;
  reg [7:0] _T_3889_43; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_261;
  reg [7:0] _T_3889_44; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_262;
  reg [7:0] _T_3889_45; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_263;
  reg [7:0] _T_3889_46; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_264;
  reg [7:0] _T_3889_47; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_265;
  reg [7:0] _T_3889_48; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_266;
  reg [7:0] _T_3889_49; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_267;
  reg [7:0] _T_3889_50; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_268;
  reg [7:0] _T_3889_51; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_269;
  reg [7:0] _T_3889_52; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_270;
  reg [7:0] _T_3889_53; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_271;
  reg [7:0] _T_3889_54; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_272;
  reg [7:0] _T_3889_55; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_273;
  reg [7:0] _T_3889_56; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_274;
  reg [7:0] _T_3889_57; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_275;
  reg [7:0] _T_3889_58; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_276;
  reg [7:0] _T_3889_59; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_277;
  reg [7:0] _T_3889_60; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_278;
  reg [7:0] _T_3889_61; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_279;
  reg [7:0] _T_3889_62; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_280;
  reg [7:0] _T_3889_63; // @[NV_NVDLA_CSC_dl.scala 1120:30:@21821.4]
  reg [31:0] _RAND_281;
  wire  _GEN_156; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_157; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_158; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_159; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_160; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_161; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_162; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_163; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_164; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_165; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_166; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_167; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_168; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_169; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_170; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_171; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_172; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_173; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_174; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_175; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_176; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_177; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_178; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_179; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_180; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_181; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_182; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_183; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_184; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_185; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_186; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_187; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_188; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_189; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_190; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_191; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_192; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_193; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_194; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_195; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_196; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_197; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_198; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_199; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_200; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_201; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_202; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_203; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_204; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_205; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_206; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_207; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_208; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_209; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_210; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_211; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_212; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_213; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_214; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_215; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_216; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_217; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_218; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _GEN_219; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  wire  _T_3956; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21892.4]
  wire  _T_3957; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21896.4]
  wire  _T_3958; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21900.4]
  wire  _T_3959; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21904.4]
  wire  _T_3960; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21908.4]
  wire  _T_3961; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21912.4]
  wire  _T_3962; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21916.4]
  wire  _T_3963; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21920.4]
  wire  _T_3964; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21924.4]
  wire  _T_3965; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21928.4]
  wire  _T_3966; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21932.4]
  wire  _T_3967; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21936.4]
  wire  _T_3968; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21940.4]
  wire  _T_3969; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21944.4]
  wire  _T_3970; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21948.4]
  wire  _T_3971; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21952.4]
  wire  _T_3972; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21956.4]
  wire  _T_3973; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21960.4]
  wire  _T_3974; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21964.4]
  wire  _T_3975; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21968.4]
  wire  _T_3976; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21972.4]
  wire  _T_3977; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21976.4]
  wire  _T_3978; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21980.4]
  wire  _T_3979; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21984.4]
  wire  _T_3980; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21988.4]
  wire  _T_3981; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21992.4]
  wire  _T_3982; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21996.4]
  wire  _T_3983; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22000.4]
  wire  _T_3984; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22004.4]
  wire  _T_3985; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22008.4]
  wire  _T_3986; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22012.4]
  wire  _T_3987; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22016.4]
  wire  _T_3988; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22020.4]
  wire  _T_3989; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22024.4]
  wire  _T_3990; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22028.4]
  wire  _T_3991; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22032.4]
  wire  _T_3992; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22036.4]
  wire  _T_3993; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22040.4]
  wire  _T_3994; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22044.4]
  wire  _T_3995; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22048.4]
  wire  _T_3996; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22052.4]
  wire  _T_3997; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22056.4]
  wire  _T_3998; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22060.4]
  wire  _T_3999; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22064.4]
  wire  _T_4000; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22068.4]
  wire  _T_4001; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22072.4]
  wire  _T_4002; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22076.4]
  wire  _T_4003; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22080.4]
  wire  _T_4004; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22084.4]
  wire  _T_4005; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22088.4]
  wire  _T_4006; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22092.4]
  wire  _T_4007; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22096.4]
  wire  _T_4008; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22100.4]
  wire  _T_4009; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22104.4]
  wire  _T_4010; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22108.4]
  wire  _T_4011; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22112.4]
  wire  _T_4012; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22116.4]
  wire  _T_4013; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22120.4]
  wire  _T_4014; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22124.4]
  wire  _T_4015; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22128.4]
  wire  _T_4016; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22132.4]
  wire  _T_4017; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22136.4]
  wire  _T_4018; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22140.4]
  wire  _T_4019; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22144.4]
  reg  _T_4022; // @[NV_NVDLA_CSC_dl.scala 1145:26:@22148.4]
  reg [31:0] _RAND_282;
  reg  _T_4289_0; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_283;
  reg  _T_4289_1; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_284;
  reg  _T_4289_2; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_285;
  reg  _T_4289_3; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_286;
  reg  _T_4289_4; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_287;
  reg  _T_4289_5; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_288;
  reg  _T_4289_6; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_289;
  reg  _T_4289_7; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_290;
  reg  _T_4289_8; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_291;
  reg  _T_4289_9; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_292;
  reg  _T_4289_10; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_293;
  reg  _T_4289_11; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_294;
  reg  _T_4289_12; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_295;
  reg  _T_4289_13; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_296;
  reg  _T_4289_14; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_297;
  reg  _T_4289_15; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_298;
  reg  _T_4289_16; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_299;
  reg  _T_4289_17; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_300;
  reg  _T_4289_18; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_301;
  reg  _T_4289_19; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_302;
  reg  _T_4289_20; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_303;
  reg  _T_4289_21; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_304;
  reg  _T_4289_22; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_305;
  reg  _T_4289_23; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_306;
  reg  _T_4289_24; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_307;
  reg  _T_4289_25; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_308;
  reg  _T_4289_26; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_309;
  reg  _T_4289_27; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_310;
  reg  _T_4289_28; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_311;
  reg  _T_4289_29; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_312;
  reg  _T_4289_30; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_313;
  reg  _T_4289_31; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_314;
  reg  _T_4289_32; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_315;
  reg  _T_4289_33; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_316;
  reg  _T_4289_34; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_317;
  reg  _T_4289_35; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_318;
  reg  _T_4289_36; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_319;
  reg  _T_4289_37; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_320;
  reg  _T_4289_38; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_321;
  reg  _T_4289_39; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_322;
  reg  _T_4289_40; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_323;
  reg  _T_4289_41; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_324;
  reg  _T_4289_42; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_325;
  reg  _T_4289_43; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_326;
  reg  _T_4289_44; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_327;
  reg  _T_4289_45; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_328;
  reg  _T_4289_46; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_329;
  reg  _T_4289_47; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_330;
  reg  _T_4289_48; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_331;
  reg  _T_4289_49; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_332;
  reg  _T_4289_50; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_333;
  reg  _T_4289_51; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_334;
  reg  _T_4289_52; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_335;
  reg  _T_4289_53; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_336;
  reg  _T_4289_54; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_337;
  reg  _T_4289_55; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_338;
  reg  _T_4289_56; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_339;
  reg  _T_4289_57; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_340;
  reg  _T_4289_58; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_341;
  reg  _T_4289_59; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_342;
  reg  _T_4289_60; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_343;
  reg  _T_4289_61; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_344;
  reg  _T_4289_62; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_345;
  reg  _T_4289_63; // @[NV_NVDLA_CSC_dl.scala 1146:26:@22214.4]
  reg [31:0] _RAND_346;
  reg [8:0] _T_4488; // @[NV_NVDLA_CSC_dl.scala 1147:26:@22215.4]
  reg [31:0] _RAND_347;
  reg [7:0] _T_4492_0; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_348;
  reg [7:0] _T_4492_1; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_349;
  reg [7:0] _T_4492_2; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_350;
  reg [7:0] _T_4492_3; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_351;
  reg [7:0] _T_4492_4; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_352;
  reg [7:0] _T_4492_5; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_353;
  reg [7:0] _T_4492_6; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_354;
  reg [7:0] _T_4492_7; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_355;
  reg [7:0] _T_4492_8; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_356;
  reg [7:0] _T_4492_9; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_357;
  reg [7:0] _T_4492_10; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_358;
  reg [7:0] _T_4492_11; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_359;
  reg [7:0] _T_4492_12; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_360;
  reg [7:0] _T_4492_13; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_361;
  reg [7:0] _T_4492_14; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_362;
  reg [7:0] _T_4492_15; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_363;
  reg [7:0] _T_4492_16; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_364;
  reg [7:0] _T_4492_17; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_365;
  reg [7:0] _T_4492_18; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_366;
  reg [7:0] _T_4492_19; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_367;
  reg [7:0] _T_4492_20; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_368;
  reg [7:0] _T_4492_21; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_369;
  reg [7:0] _T_4492_22; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_370;
  reg [7:0] _T_4492_23; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_371;
  reg [7:0] _T_4492_24; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_372;
  reg [7:0] _T_4492_25; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_373;
  reg [7:0] _T_4492_26; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_374;
  reg [7:0] _T_4492_27; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_375;
  reg [7:0] _T_4492_28; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_376;
  reg [7:0] _T_4492_29; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_377;
  reg [7:0] _T_4492_30; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_378;
  reg [7:0] _T_4492_31; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_379;
  reg [7:0] _T_4492_32; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_380;
  reg [7:0] _T_4492_33; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_381;
  reg [7:0] _T_4492_34; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_382;
  reg [7:0] _T_4492_35; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_383;
  reg [7:0] _T_4492_36; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_384;
  reg [7:0] _T_4492_37; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_385;
  reg [7:0] _T_4492_38; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_386;
  reg [7:0] _T_4492_39; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_387;
  reg [7:0] _T_4492_40; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_388;
  reg [7:0] _T_4492_41; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_389;
  reg [7:0] _T_4492_42; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_390;
  reg [7:0] _T_4492_43; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_391;
  reg [7:0] _T_4492_44; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_392;
  reg [7:0] _T_4492_45; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_393;
  reg [7:0] _T_4492_46; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_394;
  reg [7:0] _T_4492_47; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_395;
  reg [7:0] _T_4492_48; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_396;
  reg [7:0] _T_4492_49; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_397;
  reg [7:0] _T_4492_50; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_398;
  reg [7:0] _T_4492_51; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_399;
  reg [7:0] _T_4492_52; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_400;
  reg [7:0] _T_4492_53; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_401;
  reg [7:0] _T_4492_54; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_402;
  reg [7:0] _T_4492_55; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_403;
  reg [7:0] _T_4492_56; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_404;
  reg [7:0] _T_4492_57; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_405;
  reg [7:0] _T_4492_58; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_406;
  reg [7:0] _T_4492_59; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_407;
  reg [7:0] _T_4492_60; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_408;
  reg [7:0] _T_4492_61; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_409;
  reg [7:0] _T_4492_62; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_410;
  reg [7:0] _T_4492_63; // @[NV_NVDLA_CSC_dl.scala 1148:22:@22216.4]
  reg [31:0] _RAND_411;
  wire  _T_4559; // @[NV_NVDLA_CSC_dl.scala 1151:24:@22217.4]
  wire  _T_4694_0; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_1; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_2; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_3; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_4; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_5; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_6; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_7; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_8; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_9; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_10; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_11; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_12; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_13; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_14; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_15; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_16; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_17; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_18; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_19; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_20; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_21; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_22; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_23; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_24; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_25; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_26; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_27; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_28; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_29; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_30; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_31; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_32; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_33; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_34; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_35; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_36; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_37; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_38; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_39; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_40; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_41; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_42; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_43; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_44; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_45; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_46; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_47; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_48; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_49; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_50; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_51; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_52; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_53; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_54; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_55; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_56; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_57; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_58; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_59; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_60; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_61; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_62; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4694_63; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  wire  _T_4826; // @[NV_NVDLA_CSC_dl.scala 1155:19:@22285.4]
  wire  _GEN_284; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_285; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_286; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_287; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_288; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_289; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_290; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_291; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_292; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_293; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_294; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_295; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_296; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_297; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_298; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_299; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_300; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_301; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_302; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_303; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_304; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_305; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_306; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_307; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_308; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_309; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_310; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_311; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_312; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_313; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_314; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_315; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_316; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_317; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_318; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_319; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_320; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_321; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_322; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_323; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_324; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_325; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_326; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_327; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_328; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_329; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_330; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_331; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_332; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_333; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_334; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_335; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_336; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_337; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_338; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_339; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_340; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_341; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_342; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_343; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_344; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_345; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_346; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire  _GEN_347; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  wire [8:0] _GEN_348; // @[NV_NVDLA_CSC_dl.scala 1158:19:@22352.4]
  reg  _T_4829; // @[NV_NVDLA_CSC_dl.scala 1171:29:@22547.4]
  reg [31:0] _RAND_412;
  wire  _T_4830; // @[NV_NVDLA_CSC_dl.scala 1172:27:@22549.4]
  wire [8:0] _T_4832; // @[NV_NVDLA_CSC_dl.scala 1172:26:@22550.4]
  reg  _T_4835; // @[NV_NVDLA_CSC_dl.scala 1174:33:@22551.4]
  reg [31:0] _RAND_413;
  reg  _T_4838; // @[NV_NVDLA_CSC_dl.scala 1175:33:@22554.4]
  reg [31:0] _RAND_414;
  wire  _T_4840; // @[NV_NVDLA_CSC_dl.scala 1176:85:@22557.4]
  reg [8:0] _T_4842; // @[Reg.scala 19:20:@22558.4]
  reg [31:0] _RAND_415;
  wire [8:0] _GEN_413; // @[Reg.scala 20:19:@22559.4]
  reg [8:0] _T_4846; // @[Reg.scala 19:20:@22564.4]
  reg [31:0] _RAND_416;
  wire [8:0] _GEN_414; // @[Reg.scala 20:19:@22565.4]
  reg  _T_5114_0; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_417;
  reg  _T_5114_1; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_418;
  reg  _T_5114_2; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_419;
  reg  _T_5114_3; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_420;
  reg  _T_5114_4; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_421;
  reg  _T_5114_5; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_422;
  reg  _T_5114_6; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_423;
  reg  _T_5114_7; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_424;
  reg  _T_5114_8; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_425;
  reg  _T_5114_9; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_426;
  reg  _T_5114_10; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_427;
  reg  _T_5114_11; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_428;
  reg  _T_5114_12; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_429;
  reg  _T_5114_13; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_430;
  reg  _T_5114_14; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_431;
  reg  _T_5114_15; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_432;
  reg  _T_5114_16; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_433;
  reg  _T_5114_17; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_434;
  reg  _T_5114_18; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_435;
  reg  _T_5114_19; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_436;
  reg  _T_5114_20; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_437;
  reg  _T_5114_21; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_438;
  reg  _T_5114_22; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_439;
  reg  _T_5114_23; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_440;
  reg  _T_5114_24; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_441;
  reg  _T_5114_25; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_442;
  reg  _T_5114_26; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_443;
  reg  _T_5114_27; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_444;
  reg  _T_5114_28; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_445;
  reg  _T_5114_29; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_446;
  reg  _T_5114_30; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_447;
  reg  _T_5114_31; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_448;
  reg  _T_5114_32; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_449;
  reg  _T_5114_33; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_450;
  reg  _T_5114_34; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_451;
  reg  _T_5114_35; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_452;
  reg  _T_5114_36; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_453;
  reg  _T_5114_37; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_454;
  reg  _T_5114_38; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_455;
  reg  _T_5114_39; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_456;
  reg  _T_5114_40; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_457;
  reg  _T_5114_41; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_458;
  reg  _T_5114_42; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_459;
  reg  _T_5114_43; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_460;
  reg  _T_5114_44; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_461;
  reg  _T_5114_45; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_462;
  reg  _T_5114_46; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_463;
  reg  _T_5114_47; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_464;
  reg  _T_5114_48; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_465;
  reg  _T_5114_49; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_466;
  reg  _T_5114_50; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_467;
  reg  _T_5114_51; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_468;
  reg  _T_5114_52; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_469;
  reg  _T_5114_53; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_470;
  reg  _T_5114_54; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_471;
  reg  _T_5114_55; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_472;
  reg  _T_5114_56; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_473;
  reg  _T_5114_57; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_474;
  reg  _T_5114_58; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_475;
  reg  _T_5114_59; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_476;
  reg  _T_5114_60; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_477;
  reg  _T_5114_61; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_478;
  reg  _T_5114_62; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_479;
  reg  _T_5114_63; // @[Reg.scala 19:20:@22635.4]
  reg [31:0] _RAND_480;
  wire  _GEN_415; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_416; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_417; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_418; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_419; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_420; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_421; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_422; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_423; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_424; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_425; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_426; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_427; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_428; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_429; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_430; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_431; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_432; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_433; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_434; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_435; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_436; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_437; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_438; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_439; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_440; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_441; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_442; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_443; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_444; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_445; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_446; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_447; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_448; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_449; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_450; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_451; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_452; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_453; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_454; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_455; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_456; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_457; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_458; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_459; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_460; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_461; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_462; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_463; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_464; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_465; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_466; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_467; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_468; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_469; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_470; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_471; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_472; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_473; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_474; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_475; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_476; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_477; // @[Reg.scala 20:19:@22636.4]
  wire  _GEN_478; // @[Reg.scala 20:19:@22636.4]
  reg  _T_5578_0; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_481;
  reg  _T_5578_1; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_482;
  reg  _T_5578_2; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_483;
  reg  _T_5578_3; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_484;
  reg  _T_5578_4; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_485;
  reg  _T_5578_5; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_486;
  reg  _T_5578_6; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_487;
  reg  _T_5578_7; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_488;
  reg  _T_5578_8; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_489;
  reg  _T_5578_9; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_490;
  reg  _T_5578_10; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_491;
  reg  _T_5578_11; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_492;
  reg  _T_5578_12; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_493;
  reg  _T_5578_13; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_494;
  reg  _T_5578_14; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_495;
  reg  _T_5578_15; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_496;
  reg  _T_5578_16; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_497;
  reg  _T_5578_17; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_498;
  reg  _T_5578_18; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_499;
  reg  _T_5578_19; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_500;
  reg  _T_5578_20; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_501;
  reg  _T_5578_21; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_502;
  reg  _T_5578_22; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_503;
  reg  _T_5578_23; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_504;
  reg  _T_5578_24; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_505;
  reg  _T_5578_25; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_506;
  reg  _T_5578_26; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_507;
  reg  _T_5578_27; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_508;
  reg  _T_5578_28; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_509;
  reg  _T_5578_29; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_510;
  reg  _T_5578_30; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_511;
  reg  _T_5578_31; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_512;
  reg  _T_5578_32; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_513;
  reg  _T_5578_33; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_514;
  reg  _T_5578_34; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_515;
  reg  _T_5578_35; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_516;
  reg  _T_5578_36; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_517;
  reg  _T_5578_37; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_518;
  reg  _T_5578_38; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_519;
  reg  _T_5578_39; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_520;
  reg  _T_5578_40; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_521;
  reg  _T_5578_41; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_522;
  reg  _T_5578_42; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_523;
  reg  _T_5578_43; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_524;
  reg  _T_5578_44; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_525;
  reg  _T_5578_45; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_526;
  reg  _T_5578_46; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_527;
  reg  _T_5578_47; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_528;
  reg  _T_5578_48; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_529;
  reg  _T_5578_49; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_530;
  reg  _T_5578_50; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_531;
  reg  _T_5578_51; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_532;
  reg  _T_5578_52; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_533;
  reg  _T_5578_53; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_534;
  reg  _T_5578_54; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_535;
  reg  _T_5578_55; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_536;
  reg  _T_5578_56; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_537;
  reg  _T_5578_57; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_538;
  reg  _T_5578_58; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_539;
  reg  _T_5578_59; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_540;
  reg  _T_5578_60; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_541;
  reg  _T_5578_61; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_542;
  reg  _T_5578_62; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_543;
  reg  _T_5578_63; // @[Reg.scala 19:20:@22832.4]
  reg [31:0] _RAND_544;
  wire  _GEN_479; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_480; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_481; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_482; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_483; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_484; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_485; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_486; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_487; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_488; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_489; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_490; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_491; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_492; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_493; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_494; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_495; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_496; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_497; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_498; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_499; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_500; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_501; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_502; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_503; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_504; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_505; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_506; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_507; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_508; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_509; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_510; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_511; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_512; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_513; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_514; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_515; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_516; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_517; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_518; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_519; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_520; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_521; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_522; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_523; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_524; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_525; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_526; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_527; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_528; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_529; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_530; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_531; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_532; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_533; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_534; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_535; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_536; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_537; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_538; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_539; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_540; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_541; // @[Reg.scala 20:19:@22833.4]
  wire  _GEN_542; // @[Reg.scala 20:19:@22833.4]
  reg [7:0] _T_5776; // @[Reg.scala 11:16:@22963.4]
  reg [31:0] _RAND_545;
  reg [7:0] _T_5778; // @[Reg.scala 11:16:@22968.4]
  reg [31:0] _RAND_546;
  reg [7:0] _T_5780; // @[Reg.scala 11:16:@22973.4]
  reg [31:0] _RAND_547;
  reg [7:0] _T_5782; // @[Reg.scala 11:16:@22978.4]
  reg [31:0] _RAND_548;
  reg [7:0] _T_5784; // @[Reg.scala 11:16:@22983.4]
  reg [31:0] _RAND_549;
  reg [7:0] _T_5786; // @[Reg.scala 11:16:@22988.4]
  reg [31:0] _RAND_550;
  reg [7:0] _T_5788; // @[Reg.scala 11:16:@22993.4]
  reg [31:0] _RAND_551;
  reg [7:0] _T_5790; // @[Reg.scala 11:16:@22998.4]
  reg [31:0] _RAND_552;
  reg [7:0] _T_5792; // @[Reg.scala 11:16:@23003.4]
  reg [31:0] _RAND_553;
  reg [7:0] _T_5794; // @[Reg.scala 11:16:@23008.4]
  reg [31:0] _RAND_554;
  reg [7:0] _T_5796; // @[Reg.scala 11:16:@23013.4]
  reg [31:0] _RAND_555;
  reg [7:0] _T_5798; // @[Reg.scala 11:16:@23018.4]
  reg [31:0] _RAND_556;
  reg [7:0] _T_5800; // @[Reg.scala 11:16:@23023.4]
  reg [31:0] _RAND_557;
  reg [7:0] _T_5802; // @[Reg.scala 11:16:@23028.4]
  reg [31:0] _RAND_558;
  reg [7:0] _T_5804; // @[Reg.scala 11:16:@23033.4]
  reg [31:0] _RAND_559;
  reg [7:0] _T_5806; // @[Reg.scala 11:16:@23038.4]
  reg [31:0] _RAND_560;
  reg [7:0] _T_5808; // @[Reg.scala 11:16:@23043.4]
  reg [31:0] _RAND_561;
  reg [7:0] _T_5810; // @[Reg.scala 11:16:@23048.4]
  reg [31:0] _RAND_562;
  reg [7:0] _T_5812; // @[Reg.scala 11:16:@23053.4]
  reg [31:0] _RAND_563;
  reg [7:0] _T_5814; // @[Reg.scala 11:16:@23058.4]
  reg [31:0] _RAND_564;
  reg [7:0] _T_5816; // @[Reg.scala 11:16:@23063.4]
  reg [31:0] _RAND_565;
  reg [7:0] _T_5818; // @[Reg.scala 11:16:@23068.4]
  reg [31:0] _RAND_566;
  reg [7:0] _T_5820; // @[Reg.scala 11:16:@23073.4]
  reg [31:0] _RAND_567;
  reg [7:0] _T_5822; // @[Reg.scala 11:16:@23078.4]
  reg [31:0] _RAND_568;
  reg [7:0] _T_5824; // @[Reg.scala 11:16:@23083.4]
  reg [31:0] _RAND_569;
  reg [7:0] _T_5826; // @[Reg.scala 11:16:@23088.4]
  reg [31:0] _RAND_570;
  reg [7:0] _T_5828; // @[Reg.scala 11:16:@23093.4]
  reg [31:0] _RAND_571;
  reg [7:0] _T_5830; // @[Reg.scala 11:16:@23098.4]
  reg [31:0] _RAND_572;
  reg [7:0] _T_5832; // @[Reg.scala 11:16:@23103.4]
  reg [31:0] _RAND_573;
  reg [7:0] _T_5834; // @[Reg.scala 11:16:@23108.4]
  reg [31:0] _RAND_574;
  reg [7:0] _T_5836; // @[Reg.scala 11:16:@23113.4]
  reg [31:0] _RAND_575;
  reg [7:0] _T_5838; // @[Reg.scala 11:16:@23118.4]
  reg [31:0] _RAND_576;
  reg [7:0] _T_5840; // @[Reg.scala 11:16:@23123.4]
  reg [31:0] _RAND_577;
  reg [7:0] _T_5842; // @[Reg.scala 11:16:@23128.4]
  reg [31:0] _RAND_578;
  reg [7:0] _T_5844; // @[Reg.scala 11:16:@23133.4]
  reg [31:0] _RAND_579;
  reg [7:0] _T_5846; // @[Reg.scala 11:16:@23138.4]
  reg [31:0] _RAND_580;
  reg [7:0] _T_5848; // @[Reg.scala 11:16:@23143.4]
  reg [31:0] _RAND_581;
  reg [7:0] _T_5850; // @[Reg.scala 11:16:@23148.4]
  reg [31:0] _RAND_582;
  reg [7:0] _T_5852; // @[Reg.scala 11:16:@23153.4]
  reg [31:0] _RAND_583;
  reg [7:0] _T_5854; // @[Reg.scala 11:16:@23158.4]
  reg [31:0] _RAND_584;
  reg [7:0] _T_5856; // @[Reg.scala 11:16:@23163.4]
  reg [31:0] _RAND_585;
  reg [7:0] _T_5858; // @[Reg.scala 11:16:@23168.4]
  reg [31:0] _RAND_586;
  reg [7:0] _T_5860; // @[Reg.scala 11:16:@23173.4]
  reg [31:0] _RAND_587;
  reg [7:0] _T_5862; // @[Reg.scala 11:16:@23178.4]
  reg [31:0] _RAND_588;
  reg [7:0] _T_5864; // @[Reg.scala 11:16:@23183.4]
  reg [31:0] _RAND_589;
  reg [7:0] _T_5866; // @[Reg.scala 11:16:@23188.4]
  reg [31:0] _RAND_590;
  reg [7:0] _T_5868; // @[Reg.scala 11:16:@23193.4]
  reg [31:0] _RAND_591;
  reg [7:0] _T_5870; // @[Reg.scala 11:16:@23198.4]
  reg [31:0] _RAND_592;
  reg [7:0] _T_5872; // @[Reg.scala 11:16:@23203.4]
  reg [31:0] _RAND_593;
  reg [7:0] _T_5874; // @[Reg.scala 11:16:@23208.4]
  reg [31:0] _RAND_594;
  reg [7:0] _T_5876; // @[Reg.scala 11:16:@23213.4]
  reg [31:0] _RAND_595;
  reg [7:0] _T_5878; // @[Reg.scala 11:16:@23218.4]
  reg [31:0] _RAND_596;
  reg [7:0] _T_5880; // @[Reg.scala 11:16:@23223.4]
  reg [31:0] _RAND_597;
  reg [7:0] _T_5882; // @[Reg.scala 11:16:@23228.4]
  reg [31:0] _RAND_598;
  reg [7:0] _T_5884; // @[Reg.scala 11:16:@23233.4]
  reg [31:0] _RAND_599;
  reg [7:0] _T_5886; // @[Reg.scala 11:16:@23238.4]
  reg [31:0] _RAND_600;
  reg [7:0] _T_5888; // @[Reg.scala 11:16:@23243.4]
  reg [31:0] _RAND_601;
  reg [7:0] _T_5890; // @[Reg.scala 11:16:@23248.4]
  reg [31:0] _RAND_602;
  reg [7:0] _T_5892; // @[Reg.scala 11:16:@23253.4]
  reg [31:0] _RAND_603;
  reg [7:0] _T_5894; // @[Reg.scala 11:16:@23258.4]
  reg [31:0] _RAND_604;
  reg [7:0] _T_5896; // @[Reg.scala 11:16:@23263.4]
  reg [31:0] _RAND_605;
  reg [7:0] _T_5898; // @[Reg.scala 11:16:@23268.4]
  reg [31:0] _RAND_606;
  reg [7:0] _T_5900; // @[Reg.scala 11:16:@23273.4]
  reg [31:0] _RAND_607;
  reg [7:0] _T_5902; // @[Reg.scala 11:16:@23278.4]
  reg [31:0] _RAND_608;
  reg [7:0] _T_5904; // @[Reg.scala 11:16:@23283.4]
  reg [31:0] _RAND_609;
  reg [7:0] _T_5906; // @[Reg.scala 11:16:@23288.4]
  reg [31:0] _RAND_610;
  reg [7:0] _T_5908; // @[Reg.scala 11:16:@23293.4]
  reg [31:0] _RAND_611;
  reg [7:0] _T_5910; // @[Reg.scala 11:16:@23298.4]
  reg [31:0] _RAND_612;
  reg [7:0] _T_5912; // @[Reg.scala 11:16:@23303.4]
  reg [31:0] _RAND_613;
  reg [7:0] _T_5914; // @[Reg.scala 11:16:@23308.4]
  reg [31:0] _RAND_614;
  reg [7:0] _T_5916; // @[Reg.scala 11:16:@23313.4]
  reg [31:0] _RAND_615;
  reg [7:0] _T_5918; // @[Reg.scala 11:16:@23318.4]
  reg [31:0] _RAND_616;
  reg [7:0] _T_5920; // @[Reg.scala 11:16:@23323.4]
  reg [31:0] _RAND_617;
  reg [7:0] _T_5922; // @[Reg.scala 11:16:@23328.4]
  reg [31:0] _RAND_618;
  reg [7:0] _T_5924; // @[Reg.scala 11:16:@23333.4]
  reg [31:0] _RAND_619;
  reg [7:0] _T_5926; // @[Reg.scala 11:16:@23338.4]
  reg [31:0] _RAND_620;
  reg [7:0] _T_5928; // @[Reg.scala 11:16:@23343.4]
  reg [31:0] _RAND_621;
  reg [7:0] _T_5930; // @[Reg.scala 11:16:@23348.4]
  reg [31:0] _RAND_622;
  reg [7:0] _T_5932; // @[Reg.scala 11:16:@23353.4]
  reg [31:0] _RAND_623;
  reg [7:0] _T_5934; // @[Reg.scala 11:16:@23358.4]
  reg [31:0] _RAND_624;
  reg [7:0] _T_5936; // @[Reg.scala 11:16:@23363.4]
  reg [31:0] _RAND_625;
  reg [7:0] _T_5938; // @[Reg.scala 11:16:@23368.4]
  reg [31:0] _RAND_626;
  reg [7:0] _T_5940; // @[Reg.scala 11:16:@23373.4]
  reg [31:0] _RAND_627;
  reg [7:0] _T_5942; // @[Reg.scala 11:16:@23378.4]
  reg [31:0] _RAND_628;
  reg [7:0] _T_5944; // @[Reg.scala 11:16:@23383.4]
  reg [31:0] _RAND_629;
  reg [7:0] _T_5946; // @[Reg.scala 11:16:@23388.4]
  reg [31:0] _RAND_630;
  reg [7:0] _T_5948; // @[Reg.scala 11:16:@23393.4]
  reg [31:0] _RAND_631;
  reg [7:0] _T_5950; // @[Reg.scala 11:16:@23398.4]
  reg [31:0] _RAND_632;
  reg [7:0] _T_5952; // @[Reg.scala 11:16:@23403.4]
  reg [31:0] _RAND_633;
  reg [7:0] _T_5954; // @[Reg.scala 11:16:@23408.4]
  reg [31:0] _RAND_634;
  reg [7:0] _T_5956; // @[Reg.scala 11:16:@23413.4]
  reg [31:0] _RAND_635;
  reg [7:0] _T_5958; // @[Reg.scala 11:16:@23418.4]
  reg [31:0] _RAND_636;
  reg [7:0] _T_5960; // @[Reg.scala 11:16:@23423.4]
  reg [31:0] _RAND_637;
  reg [7:0] _T_5962; // @[Reg.scala 11:16:@23428.4]
  reg [31:0] _RAND_638;
  reg [7:0] _T_5964; // @[Reg.scala 11:16:@23433.4]
  reg [31:0] _RAND_639;
  reg [7:0] _T_5966; // @[Reg.scala 11:16:@23438.4]
  reg [31:0] _RAND_640;
  reg [7:0] _T_5968; // @[Reg.scala 11:16:@23443.4]
  reg [31:0] _RAND_641;
  reg [7:0] _T_5970; // @[Reg.scala 11:16:@23448.4]
  reg [31:0] _RAND_642;
  reg [7:0] _T_5972; // @[Reg.scala 11:16:@23453.4]
  reg [31:0] _RAND_643;
  reg [7:0] _T_5974; // @[Reg.scala 11:16:@23458.4]
  reg [31:0] _RAND_644;
  reg [7:0] _T_5976; // @[Reg.scala 11:16:@23463.4]
  reg [31:0] _RAND_645;
  reg [7:0] _T_5978; // @[Reg.scala 11:16:@23468.4]
  reg [31:0] _RAND_646;
  reg [7:0] _T_5980; // @[Reg.scala 11:16:@23473.4]
  reg [31:0] _RAND_647;
  reg [7:0] _T_5982; // @[Reg.scala 11:16:@23478.4]
  reg [31:0] _RAND_648;
  reg [7:0] _T_5984; // @[Reg.scala 11:16:@23483.4]
  reg [31:0] _RAND_649;
  reg [7:0] _T_5986; // @[Reg.scala 11:16:@23488.4]
  reg [31:0] _RAND_650;
  reg [7:0] _T_5988; // @[Reg.scala 11:16:@23493.4]
  reg [31:0] _RAND_651;
  reg [7:0] _T_5990; // @[Reg.scala 11:16:@23498.4]
  reg [31:0] _RAND_652;
  reg [7:0] _T_5992; // @[Reg.scala 11:16:@23503.4]
  reg [31:0] _RAND_653;
  reg [7:0] _T_5994; // @[Reg.scala 11:16:@23508.4]
  reg [31:0] _RAND_654;
  reg [7:0] _T_5996; // @[Reg.scala 11:16:@23513.4]
  reg [31:0] _RAND_655;
  reg [7:0] _T_5998; // @[Reg.scala 11:16:@23518.4]
  reg [31:0] _RAND_656;
  reg [7:0] _T_6000; // @[Reg.scala 11:16:@23523.4]
  reg [31:0] _RAND_657;
  reg [7:0] _T_6002; // @[Reg.scala 11:16:@23528.4]
  reg [31:0] _RAND_658;
  reg [7:0] _T_6004; // @[Reg.scala 11:16:@23533.4]
  reg [31:0] _RAND_659;
  reg [7:0] _T_6006; // @[Reg.scala 11:16:@23538.4]
  reg [31:0] _RAND_660;
  reg [7:0] _T_6008; // @[Reg.scala 11:16:@23543.4]
  reg [31:0] _RAND_661;
  reg [7:0] _T_6010; // @[Reg.scala 11:16:@23548.4]
  reg [31:0] _RAND_662;
  reg [7:0] _T_6012; // @[Reg.scala 11:16:@23553.4]
  reg [31:0] _RAND_663;
  reg [7:0] _T_6014; // @[Reg.scala 11:16:@23558.4]
  reg [31:0] _RAND_664;
  reg [7:0] _T_6016; // @[Reg.scala 11:16:@23563.4]
  reg [31:0] _RAND_665;
  reg [7:0] _T_6018; // @[Reg.scala 11:16:@23568.4]
  reg [31:0] _RAND_666;
  reg [7:0] _T_6020; // @[Reg.scala 11:16:@23573.4]
  reg [31:0] _RAND_667;
  reg [7:0] _T_6022; // @[Reg.scala 11:16:@23578.4]
  reg [31:0] _RAND_668;
  reg [7:0] _T_6024; // @[Reg.scala 11:16:@23583.4]
  reg [31:0] _RAND_669;
  reg [7:0] _T_6026; // @[Reg.scala 11:16:@23588.4]
  reg [31:0] _RAND_670;
  reg [7:0] _T_6028; // @[Reg.scala 11:16:@23593.4]
  reg [31:0] _RAND_671;
  reg [7:0] _T_6030; // @[Reg.scala 11:16:@23598.4]
  reg [31:0] _RAND_672;
  assign _T_622 = io_sc_state == 2'h0; // @[NV_NVDLA_CSC_dl.scala 75:31:@19633.4]
  assign _T_626 = io_sc_state == 2'h3; // @[NV_NVDLA_CSC_dl.scala 77:31:@19635.4]
  assign _T_630 = io_reg2dp_op_en & _T_622; // @[NV_NVDLA_CSC_dl.scala 84:32:@19638.4]
  assign _T_634 = io_reg2dp_conv_mode == 1'h0; // @[NV_NVDLA_CSC_dl.scala 86:35:@19640.4]
  assign _T_635 = _T_634 & io_reg2dp_datain_format; // @[NV_NVDLA_CSC_dl.scala 87:22:@19641.4]
  assign _T_640 = 7'h9 << io_reg2dp_y_extension; // @[NV_NVDLA_CSC_dl.scala 94:53:@19642.4]
  assign _T_642 = _T_635 ? _T_640 : 7'h8; // @[NV_NVDLA_CSC_dl.scala 94:24:@19643.4]
  assign _T_643 = _T_642[5:3]; // @[NV_NVDLA_CSC_dl.scala 94:100:@19644.4]
  assign _T_645 = _T_635 ? _T_643 : 3'h1; // @[NV_NVDLA_CSC_dl.scala 95:22:@19645.4]
  assign _T_647 = _T_645 - 3'h1; // @[NV_NVDLA_CSC_dl.scala 96:34:@19646.4]
  assign _T_648 = $unsigned(_T_647); // @[NV_NVDLA_CSC_dl.scala 96:34:@19647.4]
  assign _T_650 = io_reg2dp_conv_x_stride_ext + 3'h1; // @[NV_NVDLA_CSC_dl.scala 97:51:@19648.4]
  assign _T_651 = io_reg2dp_datain_channel_ext[1:0]; // @[NV_NVDLA_CSC_dl.scala 98:62:@19649.4]
  assign _T_654 = {_T_650,2'h0}; // @[Cat.scala 30:58:@19650.4]
  assign _T_657 = {_T_650,1'h0}; // @[Cat.scala 30:58:@19651.4]
  assign _GEN_671 = {{1'd0}, _T_650}; // @[NV_NVDLA_CSC_dl.scala 100:74:@19652.4]
  assign _T_658 = _T_657 + _GEN_671; // @[NV_NVDLA_CSC_dl.scala 100:74:@19652.4]
  assign _T_659 = 2'h2 == _T_651; // @[Mux.scala 46:19:@19653.4]
  assign _T_660 = _T_659 ? _T_658 : {{2'd0}, _T_650}; // @[Mux.scala 46:16:@19654.4]
  assign _T_661 = 2'h3 == _T_651; // @[Mux.scala 46:19:@19655.4]
  assign _T_662 = _T_661 ? _T_654 : _T_660; // @[Mux.scala 46:16:@19656.4]
  assign _T_664 = io_reg2dp_weight_channel_ext >= 13'h40; // @[NV_NVDLA_CSC_dl.scala 102:88:@19657.4]
  assign _T_670 = io_reg2dp_weight_channel_ext[5:0]; // @[NV_NVDLA_CSC_dl.scala 102:172:@19659.4]
  assign _T_671 = _T_664 ? 6'h3f : _T_670; // @[NV_NVDLA_CSC_dl.scala 102:58:@19660.4]
  assign _T_674 = {_T_662,1'h0}; // @[Cat.scala 30:58:@19661.4]
  assign _GEN_672 = {{1'd0}, _T_662}; // @[NV_NVDLA_CSC_dl.scala 103:81:@19662.4]
  assign _T_675 = _T_674 + _GEN_672; // @[NV_NVDLA_CSC_dl.scala 103:81:@19662.4]
  assign _T_676 = _T_674 + _GEN_672; // @[NV_NVDLA_CSC_dl.scala 103:81:@19663.4]
  assign _GEN_673 = {{1'd0}, _T_670}; // @[NV_NVDLA_CSC_dl.scala 103:100:@19665.4]
  assign _T_678 = _T_676 + _GEN_673; // @[NV_NVDLA_CSC_dl.scala 103:100:@19665.4]
  assign _T_679 = _T_676 + _GEN_673; // @[NV_NVDLA_CSC_dl.scala 103:100:@19666.4]
  assign _T_682 = _T_662 + _T_670; // @[NV_NVDLA_CSC_dl.scala 104:58:@19668.4]
  assign _T_683 = _T_662 + _T_670; // @[NV_NVDLA_CSC_dl.scala 104:58:@19669.4]
  assign _T_684 = 2'h1 == io_reg2dp_y_extension; // @[Mux.scala 46:19:@19670.4]
  assign _T_685 = _T_684 ? _T_683 : _T_671; // @[Mux.scala 46:16:@19671.4]
  assign _T_686 = 2'h2 == io_reg2dp_y_extension; // @[Mux.scala 46:19:@19672.4]
  assign _T_687 = _T_686 ? _T_679 : {{1'd0}, _T_685}; // @[Mux.scala 46:16:@19673.4]
  assign _T_690 = _T_670 + 6'h1; // @[NV_NVDLA_CSC_dl.scala 105:80:@19675.4]
  assign _T_693 = {_T_662,2'h0}; // @[Cat.scala 30:58:@19676.4]
  assign _T_698 = _T_684 ? _T_674 : {{1'd0}, _T_662}; // @[Mux.scala 46:16:@19679.4]
  assign _T_700 = _T_686 ? _T_693 : {{1'd0}, _T_698}; // @[Mux.scala 46:16:@19681.4]
  assign _T_702 = {_T_662,6'h0}; // @[Cat.scala 30:58:@19682.4]
  assign _T_704 = io_reg2dp_conv_y_stride_ext + 3'h1; // @[NV_NVDLA_CSC_dl.scala 115:52:@19683.4]
  assign _T_707 = io_reg2dp_x_dilation_ext + 5'h1; // @[NV_NVDLA_CSC_dl.scala 116:60:@19684.4]
  assign _T_708 = _T_635 ? 6'h1 : _T_707; // @[NV_NVDLA_CSC_dl.scala 116:21:@19685.4]
  assign _T_711 = io_reg2dp_y_dilation_ext + 5'h1; // @[NV_NVDLA_CSC_dl.scala 117:60:@19686.4]
  assign _T_712 = _T_635 ? 6'h1 : _T_711; // @[NV_NVDLA_CSC_dl.scala 117:21:@19687.4]
  assign _T_794 = io_reg2dp_entries + 14'h1; // @[NV_NVDLA_CSC_dl.scala 133:43:@19711.4]
  assign _T_796 = _T_794 * 15'h1; // @[NV_NVDLA_CSC_dl.scala 134:41:@19713.4]
  assign _T_797 = _T_796[14:0]; // @[NV_NVDLA_CSC_dl.scala 134:56:@19714.4]
  assign _T_798 = 6'h1 * _T_712; // @[NV_NVDLA_CSC_dl.scala 136:37:@19715.4]
  assign _GEN_674 = {{9'd0}, _T_722}; // @[NV_NVDLA_CSC_dl.scala 137:34:@19716.4]
  assign _T_799 = _T_743 * _GEN_674; // @[NV_NVDLA_CSC_dl.scala 137:34:@19716.4]
  assign _T_800 = _T_799[11:0]; // @[NV_NVDLA_CSC_dl.scala 137:47:@19717.4]
  assign _GEN_675 = {{1'd0}, _T_736}; // @[NV_NVDLA_CSC_dl.scala 138:34:@19718.4]
  assign _T_801 = _T_743 * _GEN_675; // @[NV_NVDLA_CSC_dl.scala 138:34:@19718.4]
  assign _T_802 = _T_801[11:0]; // @[NV_NVDLA_CSC_dl.scala 138:51:@19719.4]
  assign _T_804 = io_reg2dp_rls_slices + 12'h1; // @[NV_NVDLA_CSC_dl.scala 139:41:@19720.4]
  assign _T_805 = io_reg2dp_rls_slices + 12'h1; // @[NV_NVDLA_CSC_dl.scala 139:41:@19721.4]
  assign _T_807 = io_reg2dp_datain_height_ext + 13'h1; // @[NV_NVDLA_CSC_dl.scala 140:77:@19722.4]
  assign _GEN_676 = {{1'd0}, io_reg2dp_rls_slices}; // @[NV_NVDLA_CSC_dl.scala 140:113:@19723.4]
  assign _T_808 = io_reg2dp_datain_height_ext - _GEN_676; // @[NV_NVDLA_CSC_dl.scala 140:113:@19723.4]
  assign _T_809 = $unsigned(_T_808); // @[NV_NVDLA_CSC_dl.scala 140:113:@19724.4]
  assign _T_810 = io_reg2dp_skip_data_rls ? _T_807 : _T_809; // @[NV_NVDLA_CSC_dl.scala 140:23:@19725.4]
  assign _T_811 = _T_715 ? _T_729 : _T_792; // @[NV_NVDLA_CSC_dl.scala 141:24:@19726.4]
  assign _GEN_677 = {{1'd0}, _T_811}; // @[NV_NVDLA_CSC_dl.scala 142:38:@19727.4]
  assign _T_812 = _T_750 * _GEN_677; // @[NV_NVDLA_CSC_dl.scala 142:38:@19727.4]
  assign _T_813 = _T_812[14:0]; // @[NV_NVDLA_CSC_dl.scala 142:54:@19728.4]
  assign _T_1038 = _T_635 ? 34'h3ffffffff : 34'h0; // @[Bitwise.scala 72:12:@19799.6]
  assign _T_1040 = io_reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CSC_dl.scala 191:38:@19801.6]
  assign _T_1041 = io_reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CSC_dl.scala 191:38:@19802.6]
  assign _T_1043 = io_reg2dp_datain_width_ext + 13'h1; // @[NV_NVDLA_CSC_dl.scala 192:48:@19804.6]
  assign _T_1049 = io_reg2dp_weight_channel_ext[12:6]; // @[NV_NVDLA_CSC_dl.scala 195:93:@19809.6]
  assign _T_1050 = {4'h0,_T_1049}; // @[Cat.scala 30:58:@19810.6]
  assign _T_1054 = {1'h0,io_reg2dp_entries}; // @[Cat.scala 30:58:@19843.6]
  assign _GEN_1 = _T_630 ? _T_1038 : _T_831; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_2 = _T_630 ? _T_1041 : _T_838; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_3 = _T_630 ? _T_1043 : _T_845; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_4 = _T_630 ? io_reg2dp_datain_width_ext : _T_852; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_5 = _T_630 ? io_reg2dp_datain_height_ext : _T_859; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_6 = _T_630 ? _T_1050 : _T_866; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_7 = _T_630 ? _T_643 : _T_869; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_8 = _T_630 ? _T_643 : _T_872; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_10 = _T_630 ? _T_643 : _T_878; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_11 = _T_630 ? _T_643 : _T_881; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_12 = _T_630 ? _T_643 : _T_884; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_13 = _T_630 ? _T_643 : _T_887; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_15 = _T_630 ? _T_643 : _T_893; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_16 = _T_630 ? _T_643 : _T_896; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_18 = _T_630 ? _T_643 : _T_902; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_19 = _T_630 ? _T_645 : _T_905; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_20 = _T_630 ? _T_645 : _T_908; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_21 = _T_630 ? _T_650 : _T_915; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_22 = _T_630 ? _T_704 : _T_922; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_24 = _T_630 ? 6'h1 : _T_722; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_25 = _T_630 ? 5'h0 : _T_932; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_26 = _T_630 ? _T_687 : _T_939; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_27 = _T_630 ? _T_690 : _T_946; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_28 = _T_630 ? _T_700 : _T_953; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_29 = _T_630 ? {{1'd0}, _T_662} : _T_960; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_30 = _T_630 ? _T_702 : _T_967; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_31 = _T_630 ? _T_708 : _T_974; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_32 = _T_630 ? _T_712 : _T_981; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_33 = _T_630 ? io_reg2dp_pad_value : _T_988; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_34 = _T_630 ? _T_794 : _T_743; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_35 = _T_630 ? _T_797 : _T_750; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_36 = _T_630 ? _T_1054 : _T_995; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_37 = _T_630 ? {{2'd0}, _T_798} : _T_736; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_38 = _T_630 ? {{2'd0}, _T_805} : _T_729; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_39 = _T_630 ? _T_810 : _T_792; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_40 = _T_630 ? io_reg2dp_dataout_width : _T_757; // @[NV_NVDLA_CSC_dl.scala 188:15:@19795.4]
  assign _GEN_43 = _T_715 ? _T_800 : _T_778; // @[NV_NVDLA_CSC_dl.scala 233:18:@19856.4]
  assign _GEN_44 = _T_715 ? _T_802 : _T_785; // @[NV_NVDLA_CSC_dl.scala 233:18:@19856.4]
  assign _GEN_45 = _T_715 ? _T_743 : _T_1002; // @[NV_NVDLA_CSC_dl.scala 233:18:@19856.4]
  assign _GEN_46 = _T_715 ? _T_743 : _T_1009; // @[NV_NVDLA_CSC_dl.scala 233:18:@19856.4]
  assign _GEN_47 = _T_715 ? _T_813 : _T_771; // @[NV_NVDLA_CSC_dl.scala 233:18:@19856.4]
  assign _GEN_48 = _T_626 ? _T_792 : _T_1016; // @[NV_NVDLA_CSC_dl.scala 240:17:@19863.4]
  assign _GEN_49 = _T_626 ? _T_813 : _T_1023; // @[NV_NVDLA_CSC_dl.scala 240:17:@19863.4]
  assign _T_1156 = _T_1016 != 14'h0; // @[NV_NVDLA_CSC_dl.scala 304:37:@19938.4]
  assign _T_1157 = io_sg2dl_reuse_rls & _T_1156; // @[NV_NVDLA_CSC_dl.scala 304:23:@19939.4]
  assign _T_2241 = _T_878[2]; // @[NV_NVDLA_CSC_dl.scala 894:32:@20853.4]
  assign _T_2242 = _T_2241 & _T_2217; // @[NV_NVDLA_CSC_dl.scala 894:36:@20854.4]
  assign _T_2243 = _T_878[1]; // @[NV_NVDLA_CSC_dl.scala 895:35:@20855.4]
  assign _T_2244 = _T_2243 & _T_2211; // @[NV_NVDLA_CSC_dl.scala 895:39:@20856.4]
  assign _T_2245 = _T_2242 | _T_2244; // @[NV_NVDLA_CSC_dl.scala 894:57:@20857.4]
  assign _T_2246 = _T_878[0]; // @[NV_NVDLA_CSC_dl.scala 896:35:@20858.4]
  assign _T_2247 = _T_2246 & _T_2208; // @[NV_NVDLA_CSC_dl.scala 896:39:@20859.4]
  assign _T_2248 = _T_2245 | _T_2247; // @[NV_NVDLA_CSC_dl.scala 895:60:@20860.4]
  assign _T_2249 = _T_881[2]; // @[NV_NVDLA_CSC_dl.scala 903:42:@20862.4]
  assign _T_2253 = _T_2249 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@20864.4]
  assign _T_2254 = _T_2253 & _T_2231; // @[NV_NVDLA_CSC_dl.scala 903:47:@20865.4]
  assign _T_2255 = _T_881[1]; // @[NV_NVDLA_CSC_dl.scala 904:42:@20866.4]
  assign _T_2259 = _T_2255 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@20868.4]
  assign _T_2260 = _T_2259 & _T_2225; // @[NV_NVDLA_CSC_dl.scala 904:47:@20869.4]
  assign _T_2261 = _T_2254 | _T_2260; // @[NV_NVDLA_CSC_dl.scala 903:66:@20870.4]
  assign _T_2262 = _T_881[0]; // @[NV_NVDLA_CSC_dl.scala 905:42:@20871.4]
  assign _T_2266 = _T_2262 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@20873.4]
  assign _T_2267 = _T_2266 & _T_2222; // @[NV_NVDLA_CSC_dl.scala 905:47:@20874.4]
  assign _T_2268 = _T_2261 | _T_2267; // @[NV_NVDLA_CSC_dl.scala 904:66:@20875.4]
  assign _T_2287 = _T_2268[17]; // @[NV_NVDLA_CSC_dl.scala 929:26:@20894.4]
  assign _T_1154 = _T_2248 & _T_2287; // @[NV_NVDLA_CSC_dl.scala 301:29:@19937.4]
  assign _T_1159 = _T_729 != 14'h0; // @[NV_NVDLA_CSC_dl.scala 304:66:@19940.4]
  assign _T_1160 = _T_1154 & _T_1159; // @[NV_NVDLA_CSC_dl.scala 304:53:@19941.4]
  assign _T_1161 = _T_1157 | _T_1160; // @[NV_NVDLA_CSC_dl.scala 304:42:@19942.4]
  assign _T_1162 = _T_1154 ? _T_729 : _T_1016; // @[NV_NVDLA_CSC_dl.scala 305:28:@19944.4]
  assign _T_1163 = _T_1154 ? _T_771 : _T_1023; // @[NV_NVDLA_CSC_dl.scala 306:29:@19946.4]
  assign _T_1094 = _T_1161 ? _T_1163 : 15'h0; // @[NV_NVDLA_CSC_dl.scala 273:28:@19886.4]
  assign _T_1102 = _T_1076 + _T_1094; // @[NV_NVDLA_CSC_dl.scala 278:37:@19893.4]
  assign _T_1103 = _T_1076 + _T_1094; // @[NV_NVDLA_CSC_dl.scala 278:37:@19894.4]
  assign _T_1109 = {_T_838,9'h0}; // @[Cat.scala 30:58:@19896.4]
  assign _GEN_678 = {{1'd0}, _T_1109}; // @[NV_NVDLA_CSC_dl.scala 279:46:@19897.4]
  assign _T_1110 = _T_1103 - _GEN_678; // @[NV_NVDLA_CSC_dl.scala 279:46:@19897.4]
  assign _T_1111 = $unsigned(_T_1110); // @[NV_NVDLA_CSC_dl.scala 279:46:@19898.4]
  assign _T_1112 = _T_1111[14:0]; // @[NV_NVDLA_CSC_dl.scala 279:46:@19899.4]
  assign _T_1119 = _T_1103 >= _GEN_678; // @[NV_NVDLA_CSC_dl.scala 280:45:@19902.4]
  assign _T_1121 = _T_1119 ? _T_1112 : _T_1103; // @[NV_NVDLA_CSC_dl.scala 281:83:@19903.4]
  assign _T_1122 = io_sc2cdma_dat_pending_req ? 15'h0 : _T_1121; // @[NV_NVDLA_CSC_dl.scala 281:25:@19904.4]
  assign _T_1148 = _T_1161 | io_sc2cdma_dat_pending_req; // @[NV_NVDLA_CSC_dl.scala 292:13:@19927.4]
  assign _GEN_52 = _T_1148 ? _T_1122 : _T_1076; // @[NV_NVDLA_CSC_dl.scala 292:25:@19928.4]
  assign _GEN_54 = _T_1161 ? _T_1162 : _T_1169; // @[Reg.scala 20:19:@19952.4]
  assign _GEN_55 = _T_1161 ? _T_1163 : _T_1172; // @[Reg.scala 20:19:@19957.4]
  assign _T_1222 = {{30'd0}, _T_1189}; // @[NV_NVDLA_CSC_dl.scala 341:19:@20000.4 NV_NVDLA_CSC_dl.scala 345:12:@20006.4]
  assign _GEN_61 = _T_1189 ? _T_1222 : _T_1225; // @[NV_NVDLA_CSC_dl.scala 349:23:@20008.4]
  assign _GEN_62 = _T_1211 ? _T_1225 : _T_1228; // @[NV_NVDLA_CSC_dl.scala 349:23:@20012.4]
  assign _GEN_63 = _T_1214 ? _T_1228 : _T_1231; // @[NV_NVDLA_CSC_dl.scala 349:23:@20016.4]
  assign _GEN_64 = _T_1217 ? _T_1231 : _T_1234; // @[NV_NVDLA_CSC_dl.scala 349:23:@20020.4]
  assign _T_1235 = _T_869[2]; // @[NV_NVDLA_CSC_dl.scala 354:30:@20023.4]
  assign _T_1236 = _T_1235 & _T_1211; // @[NV_NVDLA_CSC_dl.scala 354:34:@20024.4]
  assign _T_1237 = _T_869[1]; // @[NV_NVDLA_CSC_dl.scala 355:30:@20025.4]
  assign _T_1238 = _T_1237 & _T_1217; // @[NV_NVDLA_CSC_dl.scala 355:34:@20026.4]
  assign _T_1239 = _T_1236 | _T_1238; // @[NV_NVDLA_CSC_dl.scala 354:50:@20027.4]
  assign _T_1240 = _T_869[0]; // @[NV_NVDLA_CSC_dl.scala 356:30:@20028.4]
  assign _T_1241 = _T_1240 & _T_1220; // @[NV_NVDLA_CSC_dl.scala 356:34:@20029.4]
  assign _T_1242 = _T_1239 | _T_1241; // @[NV_NVDLA_CSC_dl.scala 355:50:@20030.4]
  assign _T_1243 = _T_872[2]; // @[NV_NVDLA_CSC_dl.scala 358:37:@20031.4]
  assign _T_1247 = _T_1243 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@20033.4]
  assign _T_1248 = _T_1247 & _T_1225; // @[NV_NVDLA_CSC_dl.scala 358:42:@20034.4]
  assign _T_1249 = _T_872[1]; // @[NV_NVDLA_CSC_dl.scala 359:37:@20035.4]
  assign _T_1253 = _T_1249 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@20037.4]
  assign _T_1254 = _T_1253 & _T_1231; // @[NV_NVDLA_CSC_dl.scala 359:42:@20038.4]
  assign _T_1255 = _T_1248 | _T_1254; // @[NV_NVDLA_CSC_dl.scala 358:56:@20039.4]
  assign _T_1256 = _T_872[0]; // @[NV_NVDLA_CSC_dl.scala 360:37:@20040.4]
  assign _T_1260 = _T_1256 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@20042.4]
  assign _T_1261 = _T_1260 & _T_1234; // @[NV_NVDLA_CSC_dl.scala 360:42:@20043.4]
  assign _T_1262 = _T_1255 | _T_1261; // @[NV_NVDLA_CSC_dl.scala 359:56:@20044.4]
  assign _T_1263 = _T_1262[4:0]; // @[NV_NVDLA_CSC_dl.scala 363:24:@20045.4]
  assign _T_1264 = _T_1262[9:5]; // @[NV_NVDLA_CSC_dl.scala 364:24:@20046.4]
  assign _T_1265 = _T_1262[16:10]; // @[NV_NVDLA_CSC_dl.scala 365:28:@20047.4]
  assign _T_1266 = _T_1262[23:17]; // @[NV_NVDLA_CSC_dl.scala 366:29:@20048.4]
  assign _T_1267 = _T_1262[25:24]; // @[NV_NVDLA_CSC_dl.scala 367:25:@20049.4]
  assign _T_1268 = _T_1262[26]; // @[NV_NVDLA_CSC_dl.scala 368:25:@20050.4]
  assign _T_1269 = _T_1262[27]; // @[NV_NVDLA_CSC_dl.scala 369:27:@20051.4]
  assign _T_1270 = _T_1262[28]; // @[NV_NVDLA_CSC_dl.scala 370:25:@20052.4]
  assign _T_1271 = _T_1262[29]; // @[NV_NVDLA_CSC_dl.scala 371:25:@20053.4]
  assign _T_1272 = _T_1262[30]; // @[NV_NVDLA_CSC_dl.scala 372:27:@20054.4]
  assign _T_1283 = _T_1279 + 5'h1; // @[NV_NVDLA_CSC_dl.scala 381:24:@20058.4]
  assign _T_1284 = _T_1279 + 5'h1; // @[NV_NVDLA_CSC_dl.scala 381:24:@20059.4]
  assign _T_1287 = _T_1279 == _T_932; // @[NV_NVDLA_CSC_dl.scala 383:27:@20063.4]
  assign _T_1285 = _T_1287 ? 5'h0 : _T_1284; // @[NV_NVDLA_CSC_dl.scala 380:17:@20060.4]
  assign _T_1286 = _T_630 ? 5'h0 : _T_1285; // @[NV_NVDLA_CSC_dl.scala 379:17:@20061.4]
  assign _T_1294 = _T_1290 + 2'h1; // @[NV_NVDLA_CSC_dl.scala 389:31:@20067.4]
  assign _T_1295 = _T_1290 + 2'h1; // @[NV_NVDLA_CSC_dl.scala 389:31:@20068.4]
  assign _GEN_682 = {{1'd0}, _T_1295}; // @[NV_NVDLA_CSC_dl.scala 390:32:@20069.4]
  assign _T_1296 = _GEN_682 == _T_905; // @[NV_NVDLA_CSC_dl.scala 390:32:@20069.4]
  assign _T_1298 = io_reg2dp_y_extension != 2'h0; // @[NV_NVDLA_CSC_dl.scala 391:61:@20071.4]
  assign _T_1346 = _T_1306 != 7'h0; // @[NV_NVDLA_CSC_dl.scala 424:37:@20108.4]
  assign _T_1347 = ~ _T_1346; // @[NV_NVDLA_CSC_dl.scala 424:24:@20109.4]
  assign _T_1349 = _T_1290 != 2'h0; // @[NV_NVDLA_CSC_dl.scala 424:56:@20110.4]
  assign _T_1350 = ~ _T_1349; // @[NV_NVDLA_CSC_dl.scala 424:44:@20111.4]
  assign _T_1351 = _T_1347 & _T_1350; // @[NV_NVDLA_CSC_dl.scala 424:42:@20112.4]
  assign _T_1353 = _T_1279 != 5'h0; // @[NV_NVDLA_CSC_dl.scala 424:75:@20113.4]
  assign _T_1354 = ~ _T_1353; // @[NV_NVDLA_CSC_dl.scala 424:63:@20114.4]
  assign _T_1355 = _T_1351 & _T_1354; // @[NV_NVDLA_CSC_dl.scala 424:61:@20115.4]
  assign _T_1357 = _T_1355 ? 1'h0 : _T_1335; // @[NV_NVDLA_CSC_dl.scala 424:22:@20116.4]
  assign _T_1358 = _T_1242 ? 1'h1 : _T_1357; // @[NV_NVDLA_CSC_dl.scala 423:22:@20117.4]
  assign _T_1299 = _T_1298 & _T_1358; // @[NV_NVDLA_CSC_dl.scala 391:66:@20072.4]
  assign _T_1300 = _T_630 | _T_1299; // @[NV_NVDLA_CSC_dl.scala 391:33:@20073.4]
  assign _T_1301 = _T_630 | _T_1296; // @[NV_NVDLA_CSC_dl.scala 393:31:@20075.6]
  assign _T_1303 = _T_1301 ? 2'h0 : _T_1295; // @[NV_NVDLA_CSC_dl.scala 393:21:@20076.6]
  assign _GEN_65 = _T_1300 ? _T_1303 : _T_1290; // @[NV_NVDLA_CSC_dl.scala 392:23:@20074.4]
  assign _T_1312 = _T_1306 + 7'h1; // @[NV_NVDLA_CSC_dl.scala 401:33:@20082.4]
  assign _T_1313 = _T_1306 + 7'h1; // @[NV_NVDLA_CSC_dl.scala 401:33:@20083.4]
  assign _T_1314 = _T_1313 == _T_1266; // @[NV_NVDLA_CSC_dl.scala 402:51:@20084.4]
  assign _T_1315 = _T_1287 & _T_1314; // @[NV_NVDLA_CSC_dl.scala 402:33:@20085.4]
  assign _T_1316 = _T_1315 & _T_1296; // @[NV_NVDLA_CSC_dl.scala 403:34:@20087.4]
  assign _T_1317 = _T_1358 & _T_1287; // @[NV_NVDLA_CSC_dl.scala 404:52:@20089.4]
  assign _T_1318 = _T_630 | _T_1317; // @[NV_NVDLA_CSC_dl.scala 404:34:@20090.4]
  assign _T_1320 = ~ _T_1296; // @[NV_NVDLA_CSC_dl.scala 408:41:@20092.6]
  assign _T_1321 = _T_1315 & _T_1320; // @[NV_NVDLA_CSC_dl.scala 408:39:@20093.6]
  assign _T_1324 = _T_1316 ? 7'h0 : _T_1313; // @[NV_NVDLA_CSC_dl.scala 409:22:@20094.6]
  assign _T_1325 = _T_1321 ? 7'h0 : _T_1324; // @[NV_NVDLA_CSC_dl.scala 408:22:@20095.6]
  assign _T_1326 = _T_630 ? 7'h0 : _T_1325; // @[NV_NVDLA_CSC_dl.scala 407:22:@20096.6]
  assign _GEN_66 = _T_1318 ? _T_1326 : _T_1306; // @[NV_NVDLA_CSC_dl.scala 406:24:@20091.4]
  assign _T_1343 = _T_1242 | _T_1329; // @[NV_NVDLA_CSC_dl.scala 422:27:@20106.4]
  assign _T_1338 = _T_1343 & _T_1315; // @[NV_NVDLA_CSC_dl.scala 419:49:@20103.4]
  assign _T_1341 = _T_1242 ? 1'h1 : _T_1329; // @[NV_NVDLA_CSC_dl.scala 420:32:@20104.4]
  assign _T_1342 = _T_1338 ? 1'h0 : _T_1341; // @[NV_NVDLA_CSC_dl.scala 419:33:@20105.4]
  assign _T_1363 = {1'h0,_T_1265}; // @[Cat.scala 30:58:@20123.4]
  assign _GEN_67 = _T_1358 ? _T_1363 : _T_1361; // @[NV_NVDLA_CSC_dl.scala 434:21:@20124.4]
  assign _GEN_683 = {{10'd0}, _T_908}; // @[NV_NVDLA_CSC_dl.scala 444:39:@20129.4]
  assign _T_1370 = _T_1366 + _GEN_683; // @[NV_NVDLA_CSC_dl.scala 444:39:@20129.4]
  assign _T_1371 = _T_1366 + _GEN_683; // @[NV_NVDLA_CSC_dl.scala 444:39:@20130.4]
  assign _T_1372 = _T_1287 & _T_1296; // @[NV_NVDLA_CSC_dl.scala 445:29:@20131.4]
  assign _T_1373 = _T_1366 >= _T_757; // @[NV_NVDLA_CSC_dl.scala 445:61:@20132.4]
  assign _T_1374 = _T_1372 & _T_1373; // @[NV_NVDLA_CSC_dl.scala 445:44:@20133.4]
  assign _T_1377 = ~ _T_1269; // @[NV_NVDLA_CSC_dl.scala 448:43:@20136.4]
  assign _T_1378 = _T_1316 & _T_1377; // @[NV_NVDLA_CSC_dl.scala 448:41:@20137.4]
  assign _T_1379 = _T_1374 ? {{9'd0}, _T_648} : _T_1371; // @[NV_NVDLA_CSC_dl.scala 449:26:@20138.4]
  assign _T_1380 = _T_1378 ? _T_1369 : _T_1379; // @[NV_NVDLA_CSC_dl.scala 448:26:@20139.4]
  assign _T_1381 = _T_630 ? {{9'd0}, _T_648} : _T_1380; // @[NV_NVDLA_CSC_dl.scala 447:26:@20140.4]
  assign _T_1383 = _T_1317 & _T_1296; // @[NV_NVDLA_CSC_dl.scala 450:70:@20142.4]
  assign _T_1384 = _T_630 | _T_1383; // @[NV_NVDLA_CSC_dl.scala 450:37:@20143.4]
  assign _T_1385 = _T_1358 & _T_1316; // @[NV_NVDLA_CSC_dl.scala 451:55:@20144.4]
  assign _T_1386 = _T_1385 & _T_1269; // @[NV_NVDLA_CSC_dl.scala 451:71:@20145.4]
  assign _T_1387 = _T_630 | _T_1386; // @[NV_NVDLA_CSC_dl.scala 451:37:@20146.4]
  assign _GEN_68 = _T_1384 ? _T_1381 : _T_1366; // @[NV_NVDLA_CSC_dl.scala 453:27:@20147.4]
  assign _GEN_69 = _T_1387 ? _T_1381 : _T_1369; // @[NV_NVDLA_CSC_dl.scala 456:27:@20150.4]
  assign _T_1391 = _T_1390 == _T_866; // @[NV_NVDLA_CSC_dl.scala 463:37:@20154.4]
  assign _T_1393 = _T_1385 & _T_1268; // @[NV_NVDLA_CSC_dl.scala 464:70:@20156.4]
  assign _T_1394 = _T_630 | _T_1393; // @[NV_NVDLA_CSC_dl.scala 464:36:@20157.4]
  assign _T_1398 = _T_1390 + 11'h1; // @[NV_NVDLA_CSC_dl.scala 469:34:@20159.6]
  assign _T_1399 = _T_1390 + 11'h1; // @[NV_NVDLA_CSC_dl.scala 469:34:@20160.6]
  assign _T_1400 = _T_1269 ? 11'h0 : _T_1399; // @[NV_NVDLA_CSC_dl.scala 468:24:@20161.6]
  assign _T_1401 = _T_630 ? 11'h0 : _T_1400; // @[NV_NVDLA_CSC_dl.scala 467:24:@20162.6]
  assign _GEN_70 = _T_1394 ? _T_1401 : _T_1390; // @[NV_NVDLA_CSC_dl.scala 466:26:@20158.4]
  assign _GEN_684 = {{8'd0}, io_reg2dp_pad_left}; // @[NV_NVDLA_CSC_dl.scala 484:41:@20174.4]
  assign _T_1430 = 13'h0 - _GEN_684; // @[NV_NVDLA_CSC_dl.scala 484:41:@20174.4]
  assign _T_1431 = $unsigned(_T_1430); // @[NV_NVDLA_CSC_dl.scala 484:41:@20175.4]
  assign _T_1432 = _T_635 ? 14'h0 : _T_1431; // @[NV_NVDLA_CSC_dl.scala 483:26:@20176.4]
  assign _GEN_685 = {{10'd0}, _T_915}; // @[NV_NVDLA_CSC_dl.scala 485:37:@20177.4]
  assign _T_1433 = _T_1404 + _GEN_685; // @[NV_NVDLA_CSC_dl.scala 485:37:@20177.4]
  assign _T_1434 = _T_1404 + _GEN_685; // @[NV_NVDLA_CSC_dl.scala 485:37:@20178.4]
  assign _T_1437 = _T_1374 ? _T_1432 : _T_1434; // @[NV_NVDLA_CSC_dl.scala 490:25:@20181.4]
  assign _T_1438 = _T_1378 ? _T_1407 : _T_1437; // @[NV_NVDLA_CSC_dl.scala 489:25:@20182.4]
  assign _T_1439 = _T_630 ? _T_1432 : _T_1438; // @[NV_NVDLA_CSC_dl.scala 488:25:@20183.4]
  assign _GEN_686 = {{1'd0}, _T_1263}; // @[NV_NVDLA_CSC_dl.scala 492:35:@20184.4]
  assign _T_1440 = _GEN_686 * _T_974; // @[NV_NVDLA_CSC_dl.scala 492:35:@20184.4]
  assign _GEN_687 = {{3'd0}, _T_1440}; // @[NV_NVDLA_CSC_dl.scala 493:33:@20185.4]
  assign _T_1441 = _T_1404 + _GEN_687; // @[NV_NVDLA_CSC_dl.scala 493:33:@20185.4]
  assign _T_1442 = _T_1404 + _GEN_687; // @[NV_NVDLA_CSC_dl.scala 493:33:@20186.4]
  assign _T_1445 = _T_831[0]; // @[NV_NVDLA_CSC_dl.scala 494:96:@20189.4]
  assign _T_1446 = ~ _T_1445; // @[NV_NVDLA_CSC_dl.scala 494:86:@20190.4]
  assign _T_1447 = _T_1383 & _T_1446; // @[NV_NVDLA_CSC_dl.scala 494:84:@20191.4]
  assign _T_1448 = _T_630 | _T_1447; // @[NV_NVDLA_CSC_dl.scala 494:36:@20192.4]
  assign _T_1451 = _T_831[1]; // @[NV_NVDLA_CSC_dl.scala 495:99:@20195.4]
  assign _T_1452 = ~ _T_1451; // @[NV_NVDLA_CSC_dl.scala 495:89:@20196.4]
  assign _T_1453 = _T_1386 & _T_1452; // @[NV_NVDLA_CSC_dl.scala 495:87:@20197.4]
  assign _T_1454 = _T_630 | _T_1453; // @[NV_NVDLA_CSC_dl.scala 495:36:@20198.4]
  assign _T_1456 = _T_1296 ? _T_953 : 8'h0; // @[NV_NVDLA_CSC_dl.scala 498:26:@20199.4]
  assign _T_1459 = _T_670 == 6'h0; // @[NV_NVDLA_CSC_dl.scala 500:79:@20201.4]
  assign _T_1463 = _T_1049 + 7'h1; // @[NV_NVDLA_CSC_dl.scala 501:74:@20204.4]
  assign _T_1464 = _T_1049 + 7'h1; // @[NV_NVDLA_CSC_dl.scala 501:74:@20205.4]
  assign _T_1465 = _T_1459 ? _T_1049 : _T_1464; // @[NV_NVDLA_CSC_dl.scala 500:27:@20206.4]
  assign _T_1466 = _T_1269 & _T_1316; // @[NV_NVDLA_CSC_dl.scala 502:37:@20207.4]
  assign _T_1468 = _T_1268 & _T_1316; // @[NV_NVDLA_CSC_dl.scala 503:35:@20208.4]
  assign _T_1470 = _T_1419 + 13'h1; // @[NV_NVDLA_CSC_dl.scala 503:66:@20209.4]
  assign _T_1471 = _T_1419 + 13'h1; // @[NV_NVDLA_CSC_dl.scala 503:66:@20210.4]
  assign _T_1472 = _T_1468 ? _T_1471 : _T_1419; // @[NV_NVDLA_CSC_dl.scala 503:22:@20211.4]
  assign _T_1473 = _T_1466 ? 13'h2 : _T_1472; // @[NV_NVDLA_CSC_dl.scala 502:22:@20212.4]
  assign _GEN_688 = {{6'd0}, _T_1465}; // @[NV_NVDLA_CSC_dl.scala 505:44:@20214.4]
  assign _T_1474 = _T_1419 >= _GEN_688; // @[NV_NVDLA_CSC_dl.scala 505:44:@20214.4]
  assign _T_1475 = _T_1316 & _T_1268; // @[NV_NVDLA_CSC_dl.scala 509:39:@20215.4]
  assign _T_1476 = _T_1475 & _T_1269; // @[NV_NVDLA_CSC_dl.scala 509:54:@20216.4]
  assign _T_1477 = _T_1476 & _T_1374; // @[NV_NVDLA_CSC_dl.scala 509:71:@20217.4]
  assign _T_1480 = ~ _T_1374; // @[NV_NVDLA_CSC_dl.scala 510:73:@20220.4]
  assign _T_1481 = _T_1476 & _T_1480; // @[NV_NVDLA_CSC_dl.scala 510:71:@20221.4]
  assign _GEN_689 = {{4'd0}, _T_967}; // @[NV_NVDLA_CSC_dl.scala 510:99:@20222.4]
  assign _T_1482 = _T_1416 + _GEN_689; // @[NV_NVDLA_CSC_dl.scala 510:99:@20222.4]
  assign _T_1483 = _T_1416 + _GEN_689; // @[NV_NVDLA_CSC_dl.scala 510:99:@20223.4]
  assign _T_1485 = _T_1475 & _T_1474; // @[NV_NVDLA_CSC_dl.scala 511:54:@20225.4]
  assign _GEN_690 = {{9'd0}, _T_946}; // @[NV_NVDLA_CSC_dl.scala 511:90:@20226.4]
  assign _T_1486 = _T_1413 + _GEN_690; // @[NV_NVDLA_CSC_dl.scala 511:90:@20226.4]
  assign _T_1487 = _T_1413 + _GEN_690; // @[NV_NVDLA_CSC_dl.scala 511:90:@20227.4]
  assign _T_1489 = ~ _T_1474; // @[NV_NVDLA_CSC_dl.scala 512:56:@20229.4]
  assign _T_1490 = _T_1475 & _T_1489; // @[NV_NVDLA_CSC_dl.scala 512:54:@20230.4]
  assign _T_1492 = _T_1413 + 16'h40; // @[NV_NVDLA_CSC_dl.scala 512:91:@20231.4]
  assign _T_1493 = _T_1413 + 16'h40; // @[NV_NVDLA_CSC_dl.scala 512:91:@20232.4]
  assign _T_1494 = ~ _T_1268; // @[NV_NVDLA_CSC_dl.scala 513:41:@20233.4]
  assign _T_1495 = _T_1316 & _T_1494; // @[NV_NVDLA_CSC_dl.scala 513:39:@20234.4]
  assign _GEN_691 = {{8'd0}, _T_1456}; // @[NV_NVDLA_CSC_dl.scala 513:81:@20235.4]
  assign _T_1496 = _T_1410 + _GEN_691; // @[NV_NVDLA_CSC_dl.scala 513:81:@20235.4]
  assign _T_1497 = _T_1410 + _GEN_691; // @[NV_NVDLA_CSC_dl.scala 513:81:@20236.4]
  assign _T_1498 = _T_1495 ? _T_1413 : _T_1497; // @[NV_NVDLA_CSC_dl.scala 513:24:@20237.4]
  assign _T_1499 = _T_1490 ? _T_1493 : _T_1498; // @[NV_NVDLA_CSC_dl.scala 512:24:@20238.4]
  assign _T_1500 = _T_1485 ? _T_1487 : _T_1499; // @[NV_NVDLA_CSC_dl.scala 511:24:@20239.4]
  assign _T_1501 = _T_1481 ? _T_1483 : _T_1500; // @[NV_NVDLA_CSC_dl.scala 510:24:@20240.4]
  assign _T_1502 = _T_1477 ? {{9'd0}, _T_939} : _T_1501; // @[NV_NVDLA_CSC_dl.scala 509:24:@20241.4]
  assign _T_1503 = _T_715 ? {{9'd0}, _T_939} : _T_1502; // @[NV_NVDLA_CSC_dl.scala 508:24:@20242.4]
  assign _T_1509 = _T_1410[15:6]; // @[NV_NVDLA_CSC_dl.scala 515:68:@20244.4]
  assign _T_1510 = {5'h0,_T_1509}; // @[Cat.scala 30:58:@20245.4]
  assign _T_1521 = _T_831[4]; // @[NV_NVDLA_CSC_dl.scala 518:68:@20256.4]
  assign _T_1522 = _T_1358 & _T_1521; // @[NV_NVDLA_CSC_dl.scala 518:57:@20257.4]
  assign _T_1523 = _T_1522 & _T_1316; // @[NV_NVDLA_CSC_dl.scala 518:72:@20258.4]
  assign _T_1524 = _T_1523 & _T_1268; // @[NV_NVDLA_CSC_dl.scala 518:88:@20259.4]
  assign _T_1525 = _T_1524 & _T_1269; // @[NV_NVDLA_CSC_dl.scala 518:103:@20260.4]
  assign _T_1526 = _T_715 | _T_1525; // @[NV_NVDLA_CSC_dl.scala 518:39:@20261.4]
  assign _T_1528 = _T_1445 & _T_1242; // @[NV_NVDLA_CSC_dl.scala 520:42:@20263.4]
  assign _T_1531 = _T_1424 ? 1'h0 : _T_1427; // @[NV_NVDLA_CSC_dl.scala 520:74:@20264.4]
  assign _T_1532 = _T_1528 ? 1'h1 : _T_1531; // @[NV_NVDLA_CSC_dl.scala 520:28:@20265.4]
  assign _T_1534 = _T_1445 & _T_1296; // @[NV_NVDLA_CSC_dl.scala 521:36:@20267.4]
  assign _T_1535 = _T_1532 | _T_1427; // @[NV_NVDLA_CSC_dl.scala 521:72:@20268.4]
  assign _T_1536 = _T_1534 & _T_1535; // @[NV_NVDLA_CSC_dl.scala 521:51:@20269.4]
  assign _GEN_71 = _T_1448 ? _T_1439 : _T_1404; // @[NV_NVDLA_CSC_dl.scala 523:26:@20270.4]
  assign _GEN_72 = _T_1448 ? _T_1503 : _T_1410; // @[NV_NVDLA_CSC_dl.scala 523:26:@20270.4]
  assign _GEN_73 = _T_1454 ? _T_1439 : _T_1407; // @[NV_NVDLA_CSC_dl.scala 527:26:@20274.4]
  assign _GEN_74 = _T_1454 ? _T_1503 : _T_1413; // @[NV_NVDLA_CSC_dl.scala 527:26:@20274.4]
  assign _GEN_75 = _T_1526 ? _T_1503 : _T_1416; // @[NV_NVDLA_CSC_dl.scala 531:26:@20278.4]
  assign _GEN_692 = {{9'd0}, io_reg2dp_pad_top}; // @[NV_NVDLA_CSC_dl.scala 540:41:@20283.4]
  assign _T_1544 = 14'h0 - _GEN_692; // @[NV_NVDLA_CSC_dl.scala 540:41:@20283.4]
  assign _T_1545 = $unsigned(_T_1544); // @[NV_NVDLA_CSC_dl.scala 540:41:@20284.4]
  assign _T_1546 = _T_1545[13:0]; // @[NV_NVDLA_CSC_dl.scala 540:41:@20285.4]
  assign _GEN_693 = {{10'd0}, _T_922}; // @[NV_NVDLA_CSC_dl.scala 541:37:@20286.4]
  assign _T_1547 = _T_1539 + _GEN_693; // @[NV_NVDLA_CSC_dl.scala 541:37:@20286.4]
  assign _T_1548 = _T_1539 + _GEN_693; // @[NV_NVDLA_CSC_dl.scala 541:37:@20287.4]
  assign _T_1549 = _T_1316 & _T_1270; // @[NV_NVDLA_CSC_dl.scala 542:52:@20288.4]
  assign _T_1550 = _T_630 | _T_1549; // @[NV_NVDLA_CSC_dl.scala 542:35:@20289.4]
  assign _T_1553 = _T_1374 ? _T_1548 : _T_1539; // @[NV_NVDLA_CSC_dl.scala 544:25:@20292.4]
  assign _T_1554 = _T_1378 ? _T_1542 : _T_1553; // @[NV_NVDLA_CSC_dl.scala 543:25:@20293.4]
  assign _T_1555 = _T_1550 ? _T_1546 : _T_1554; // @[NV_NVDLA_CSC_dl.scala 542:25:@20294.4]
  assign _T_1558 = _T_1378 | _T_1374; // @[NV_NVDLA_CSC_dl.scala 545:91:@20297.4]
  assign _T_1559 = _T_1358 & _T_1558; // @[NV_NVDLA_CSC_dl.scala 545:54:@20298.4]
  assign _T_1560 = _T_630 | _T_1559; // @[NV_NVDLA_CSC_dl.scala 545:36:@20299.4]
  assign _GEN_694 = {{1'd0}, _T_1264}; // @[NV_NVDLA_CSC_dl.scala 547:35:@20303.4]
  assign _T_1564 = _GEN_694 * _T_981; // @[NV_NVDLA_CSC_dl.scala 547:35:@20303.4]
  assign _GEN_695 = {{3'd0}, _T_1564}; // @[NV_NVDLA_CSC_dl.scala 548:33:@20304.4]
  assign _T_1565 = _T_1539 + _GEN_695; // @[NV_NVDLA_CSC_dl.scala 548:33:@20304.4]
  assign _T_1566 = _T_1539 + _GEN_695; // @[NV_NVDLA_CSC_dl.scala 548:33:@20305.4]
  assign _GEN_696 = {{12'd0}, _T_1290}; // @[NV_NVDLA_CSC_dl.scala 548:51:@20306.4]
  assign _T_1567 = _T_1566 + _GEN_696; // @[NV_NVDLA_CSC_dl.scala 548:51:@20306.4]
  assign _T_1568 = _T_1566 + _GEN_696; // @[NV_NVDLA_CSC_dl.scala 548:51:@20307.4]
  assign _GEN_76 = _T_1560 ? _T_1555 : _T_1539; // @[NV_NVDLA_CSC_dl.scala 550:26:@20308.4]
  assign _GEN_77 = _T_1387 ? _T_1555 : _T_1542; // @[NV_NVDLA_CSC_dl.scala 551:26:@20311.4]
  assign _T_1569 = _T_1442[13]; // @[NV_NVDLA_CSC_dl.scala 554:39:@20314.4]
  assign _GEN_697 = {{1'd0}, _T_852}; // @[NV_NVDLA_CSC_dl.scala 554:59:@20315.4]
  assign _T_1570 = _T_1442 > _GEN_697; // @[NV_NVDLA_CSC_dl.scala 554:59:@20315.4]
  assign _T_1571 = _T_1569 | _T_1570; // @[NV_NVDLA_CSC_dl.scala 554:44:@20316.4]
  assign _T_1572 = _T_1568[13]; // @[NV_NVDLA_CSC_dl.scala 554:92:@20317.4]
  assign _T_1573 = _T_1571 | _T_1572; // @[NV_NVDLA_CSC_dl.scala 554:78:@20318.4]
  assign _GEN_698 = {{1'd0}, _T_859}; // @[NV_NVDLA_CSC_dl.scala 554:112:@20319.4]
  assign _T_1574 = _T_1568 > _GEN_698; // @[NV_NVDLA_CSC_dl.scala 554:112:@20319.4]
  assign _T_1575 = _T_1573 | _T_1574; // @[NV_NVDLA_CSC_dl.scala 554:97:@20320.4]
  assign _T_1588 = _T_1572 | _T_1574; // @[NV_NVDLA_CSC_dl.scala 557:42:@20330.4]
  assign _T_1698 = _T_831[10]; // @[NV_NVDLA_CSC_dl.scala 642:33:@20416.4]
  assign _T_1699 = ~ _T_1391; // @[NV_NVDLA_CSC_dl.scala 643:24:@20417.4]
  assign _T_1701 = _T_1442[12:0]; // @[NV_NVDLA_CSC_dl.scala 643:77:@20418.4]
  assign _T_1702 = {2'h0,_T_1701}; // @[Cat.scala 30:58:@20419.4]
  assign _T_1704 = _T_1363 > 8'h20; // @[NV_NVDLA_CSC_dl.scala 644:38:@20420.4]
  assign _T_1709 = _T_1442[12:1]; // @[NV_NVDLA_CSC_dl.scala 645:54:@20423.4]
  assign _T_1710 = {3'h0,_T_1709}; // @[Cat.scala 30:58:@20424.4]
  assign _T_1711 = _T_1704 ? _T_1702 : _T_1710; // @[NV_NVDLA_CSC_dl.scala 644:23:@20425.4]
  assign _T_1712 = _T_1699 ? _T_1702 : _T_1711; // @[NV_NVDLA_CSC_dl.scala 643:23:@20426.4]
  assign _T_1713 = _T_1698 ? _T_1510 : _T_1712; // @[NV_NVDLA_CSC_dl.scala 642:23:@20427.4]
  assign _T_1714 = _T_1713[13:0]; // @[NV_NVDLA_CSC_dl.scala 654:24:@20429.4]
  assign _T_1591 = _T_1714[13:2]; // @[NV_NVDLA_CSC_dl.scala 561:32:@20332.4]
  assign _GEN_700 = {{3'd0}, _T_1591}; // @[NV_NVDLA_CSC_dl.scala 561:40:@20333.4]
  assign _T_1592 = _GEN_700 > _T_995; // @[NV_NVDLA_CSC_dl.scala 561:40:@20333.4]
  assign _T_1593 = _T_831[5]; // @[NV_NVDLA_CSC_dl.scala 562:34:@20334.4]
  assign _T_1594 = _T_1593 ? _T_1588 : _T_1575; // @[NV_NVDLA_CSC_dl.scala 562:24:@20335.4]
  assign _T_1595 = _T_831[6]; // @[NV_NVDLA_CSC_dl.scala 563:29:@20336.4]
  assign _T_1596 = _T_1595 & _T_1592; // @[NV_NVDLA_CSC_dl.scala 563:33:@20337.4]
  assign _T_1597 = ~ _T_1594; // @[NV_NVDLA_CSC_dl.scala 564:39:@20338.4]
  assign _T_1598 = _T_1358 & _T_1597; // @[NV_NVDLA_CSC_dl.scala 564:37:@20339.4]
  assign _T_1599 = ~ _T_1596; // @[NV_NVDLA_CSC_dl.scala 564:56:@20340.4]
  assign _T_1600 = _T_1598 & _T_1599; // @[NV_NVDLA_CSC_dl.scala 564:54:@20341.4]
  assign _T_1601 = _T_831[7]; // @[NV_NVDLA_CSC_dl.scala 567:37:@20342.4]
  assign _T_1602 = ~ _T_1601; // @[NV_NVDLA_CSC_dl.scala 567:27:@20343.4]
  assign _T_1603 = _T_1390[0]; // @[NV_NVDLA_CSC_dl.scala 567:54:@20344.4]
  assign _T_1604 = _T_1602 ? _T_1603 : _T_1268; // @[NV_NVDLA_CSC_dl.scala 567:26:@20345.4]
  assign _T_1605 = _T_1442[1:0]; // @[NV_NVDLA_CSC_dl.scala 568:35:@20346.4]
  assign _T_1607 = _T_1290 == 2'h0; // @[NV_NVDLA_CSC_dl.scala 569:55:@20347.4]
  assign _T_1608 = _T_1358 & _T_1607; // @[NV_NVDLA_CSC_dl.scala 569:42:@20348.4]
  assign _T_1609 = _T_1315 & _T_1343; // @[NV_NVDLA_CSC_dl.scala 572:42:@20350.4]
  assign _T_1613 = {_T_1271,_T_1269,_T_1609,_T_1242,_T_1279}; // @[Cat.scala 30:58:@20354.4]
  assign _T_1644 = _T_1272 & _T_1315; // @[NV_NVDLA_CSC_dl.scala 599:38:@20374.6]
  assign _T_1645 = _T_1644 & _T_1343; // @[NV_NVDLA_CSC_dl.scala 599:56:@20375.6]
  assign _GEN_78 = _T_1358 ? _T_1605 : _T_1619; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  assign _GEN_79 = _T_1358 ? _T_1290 : _T_1622; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  assign _GEN_80 = _T_1358 ? _T_1604 : _T_1625; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  assign _GEN_81 = _T_1358 ? _T_1391 : _T_1628; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  assign _GEN_82 = _T_1358 ? _T_1358 : _T_1631; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  assign _GEN_83 = _T_1358 ? _T_1267 : _T_1634; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  assign _GEN_84 = _T_1358 ? _T_1613 : _T_1640; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  assign _GEN_85 = _T_1358 ? _T_1645 : _T_1643; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  assign _GEN_86 = _T_1358 ? _T_1532 : _T_1427; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  assign _GEN_87 = _T_1358 ? _T_1536 : _T_1424; // @[NV_NVDLA_CSC_dl.scala 591:21:@20366.4]
  assign _GEN_88 = _T_1608 ? _T_1242 : _T_1637; // @[NV_NVDLA_CSC_dl.scala 603:26:@20380.4]
  assign _T_1667 = _T_831[8]; // @[NV_NVDLA_CSC_dl.scala 620:32:@20390.4]
  assign _T_1668 = ~ _T_1667; // @[NV_NVDLA_CSC_dl.scala 620:22:@20391.4]
  assign _T_1669 = _T_845[11:0]; // @[NV_NVDLA_CSC_dl.scala 620:49:@20392.4]
  assign _T_1671 = _T_1668 ? _T_1669 : 12'h0; // @[NV_NVDLA_CSC_dl.scala 620:21:@20393.4]
  assign _T_1673 = _T_1316 & _T_1269; // @[NV_NVDLA_CSC_dl.scala 622:34:@20394.4]
  assign _GEN_701 = {{1'd0}, _T_1671}; // @[NV_NVDLA_CSC_dl.scala 622:64:@20395.4]
  assign _T_1675 = _T_1648 + _GEN_701; // @[NV_NVDLA_CSC_dl.scala 622:64:@20395.4]
  assign _T_1676 = _T_1648 + _GEN_701; // @[NV_NVDLA_CSC_dl.scala 622:64:@20396.4]
  assign _T_1677 = _T_1673 ? 13'h0 : _T_1676; // @[NV_NVDLA_CSC_dl.scala 622:19:@20397.4]
  assign _T_1678 = _T_630 ? 13'h0 : _T_1677; // @[NV_NVDLA_CSC_dl.scala 621:19:@20398.4]
  assign _T_1682 = _T_1648 != _T_1651; // @[NV_NVDLA_CSC_dl.scala 624:31:@20402.4]
  assign _GEN_702 = {{2'd0}, _T_778}; // @[NV_NVDLA_CSC_dl.scala 627:32:@20403.4]
  assign _T_1683 = _T_1539 * _GEN_702; // @[NV_NVDLA_CSC_dl.scala 627:32:@20403.4]
  assign _T_1684 = _T_1683[12:0]; // @[NV_NVDLA_CSC_dl.scala 627:50:@20404.4]
  assign _GEN_703 = {{7'd0}, _T_1264}; // @[NV_NVDLA_CSC_dl.scala 628:31:@20405.4]
  assign _T_1685 = _GEN_703 * _T_785; // @[NV_NVDLA_CSC_dl.scala 628:31:@20405.4]
  assign _T_1686 = _T_1685[12:0]; // @[NV_NVDLA_CSC_dl.scala 628:49:@20406.4]
  assign _GEN_704 = {{10'd0}, _T_1279}; // @[NV_NVDLA_CSC_dl.scala 629:29:@20407.4]
  assign _T_1687 = _GEN_704 * _T_1002; // @[NV_NVDLA_CSC_dl.scala 629:29:@20407.4]
  assign _T_1688 = _T_1687[12:0]; // @[NV_NVDLA_CSC_dl.scala 629:47:@20408.4]
  assign _GEN_705 = {{13'd0}, _T_1290}; // @[NV_NVDLA_CSC_dl.scala 630:47:@20409.4]
  assign _T_1690 = _GEN_705 * _T_1009; // @[NV_NVDLA_CSC_dl.scala 630:47:@20409.4]
  assign _T_1691 = _T_630 ? 17'h0 : _T_1690; // @[NV_NVDLA_CSC_dl.scala 630:21:@20410.4]
  assign _T_1692 = _T_1691[12:0]; // @[NV_NVDLA_CSC_dl.scala 630:65:@20411.4]
  assign _T_1693 = _T_831[9]; // @[NV_NVDLA_CSC_dl.scala 631:45:@20412.4]
  assign _T_1694 = _T_630 | _T_1693; // @[NV_NVDLA_CSC_dl.scala 631:34:@20413.4]
  assign _T_1695 = {_T_1694,_T_1358}; // @[Cat.scala 30:58:@20414.4]
  assign _GEN_89 = _T_1394 ? _T_1678 : _T_1648; // @[NV_NVDLA_CSC_dl.scala 658:20:@20431.4]
  assign _GEN_90 = _T_1682 ? _T_1648 : _T_1651; // @[NV_NVDLA_CSC_dl.scala 661:23:@20434.4]
  assign _T_1715 = _T_1695[0]; // @[NV_NVDLA_CSC_dl.scala 664:19:@20437.4]
  assign _GEN_91 = _T_1715 ? _T_1684 : _T_1654; // @[NV_NVDLA_CSC_dl.scala 664:23:@20438.4]
  assign _GEN_92 = _T_1715 ? _T_1686 : _T_1657; // @[NV_NVDLA_CSC_dl.scala 664:23:@20438.4]
  assign _GEN_93 = _T_1715 ? _T_1688 : _T_1660; // @[NV_NVDLA_CSC_dl.scala 664:23:@20438.4]
  assign _T_1716 = _T_1695[1]; // @[NV_NVDLA_CSC_dl.scala 669:19:@20443.4]
  assign _GEN_94 = _T_1716 ? _T_1692 : _T_1663; // @[NV_NVDLA_CSC_dl.scala 669:23:@20444.4]
  assign _GEN_95 = _T_1358 ? _T_1714 : {{1'd0}, _T_1666}; // @[NV_NVDLA_CSC_dl.scala 672:20:@20447.4]
  assign _T_1822 = _T_1654 + _T_1657; // @[NV_NVDLA_CSC_dl.scala 696:29:@20475.4]
  assign _T_1823 = _T_1654 + _T_1657; // @[NV_NVDLA_CSC_dl.scala 696:29:@20476.4]
  assign _T_1824 = _T_1823 + _T_1660; // @[NV_NVDLA_CSC_dl.scala 696:43:@20477.4]
  assign _T_1825 = _T_1823 + _T_1660; // @[NV_NVDLA_CSC_dl.scala 696:43:@20478.4]
  assign _T_1826 = _T_1825 + _T_1663; // @[NV_NVDLA_CSC_dl.scala 696:57:@20479.4]
  assign _T_1827 = _T_1825 + _T_1663; // @[NV_NVDLA_CSC_dl.scala 696:57:@20480.4]
  assign _GEN_706 = {{2'd0}, _T_1651}; // @[NV_NVDLA_CSC_dl.scala 697:40:@20481.4]
  assign _T_1828 = _T_1076 + _GEN_706; // @[NV_NVDLA_CSC_dl.scala 697:40:@20481.4]
  assign _T_1829 = _T_1076 + _GEN_706; // @[NV_NVDLA_CSC_dl.scala 697:40:@20482.4]
  assign _GEN_707 = {{2'd0}, _T_1827}; // @[NV_NVDLA_CSC_dl.scala 697:52:@20483.4]
  assign _T_1830 = _T_1829 + _GEN_707; // @[NV_NVDLA_CSC_dl.scala 697:52:@20483.4]
  assign _T_1831 = _T_1829 + _GEN_707; // @[NV_NVDLA_CSC_dl.scala 697:52:@20484.4]
  assign _GEN_708 = {{2'd0}, _T_1666}; // @[NV_NVDLA_CSC_dl.scala 697:64:@20485.4]
  assign _T_1832 = _T_1831 + _GEN_708; // @[NV_NVDLA_CSC_dl.scala 697:64:@20485.4]
  assign _T_1833 = _T_1831 + _GEN_708; // @[NV_NVDLA_CSC_dl.scala 697:64:@20486.4]
  assign _T_1840 = _T_1833 >= _GEN_678; // @[NV_NVDLA_CSC_dl.scala 698:45:@20489.4]
  assign _T_1847 = _T_1833 - _GEN_678; // @[NV_NVDLA_CSC_dl.scala 699:42:@20492.4]
  assign _T_1848 = $unsigned(_T_1847); // @[NV_NVDLA_CSC_dl.scala 699:42:@20493.4]
  assign _T_1849 = _T_1848[14:0]; // @[NV_NVDLA_CSC_dl.scala 699:42:@20494.4]
  assign _T_1850 = _T_630 | _T_1631; // @[NV_NVDLA_CSC_dl.scala 700:35:@20495.4]
  assign _T_1856 = _T_1840 ? _T_1849 : _T_1833; // @[NV_NVDLA_CSC_dl.scala 701:25:@20497.4]
  assign _T_1857 = _T_1850 ? 15'h1fff : _T_1856; // @[NV_NVDLA_CSC_dl.scala 700:25:@20498.4]
  assign _T_1881 = 2'h3 == _T_1622; // @[Mux.scala 46:19:@20508.4]
  assign _T_1882 = _T_1881 ? _T_1759_3 : 13'h0; // @[Mux.scala 46:16:@20509.4]
  assign _T_1883 = 2'h2 == _T_1622; // @[Mux.scala 46:19:@20510.4]
  assign _T_1884 = _T_1883 ? _T_1759_2 : _T_1882; // @[Mux.scala 46:16:@20511.4]
  assign _T_1885 = 2'h1 == _T_1622; // @[Mux.scala 46:19:@20512.4]
  assign _T_1886 = _T_1885 ? _T_1759_1 : _T_1884; // @[Mux.scala 46:16:@20513.4]
  assign _T_1887 = 2'h0 == _T_1622; // @[Mux.scala 46:19:@20514.4]
  assign _T_1888 = _T_1887 ? _T_1759_0 : _T_1886; // @[Mux.scala 46:16:@20515.4]
  assign _GEN_712 = {{2'd0}, _T_1888}; // @[NV_NVDLA_CSC_dl.scala 708:65:@20516.4]
  assign _T_1889 = _GEN_712 != _T_1857; // @[NV_NVDLA_CSC_dl.scala 708:65:@20516.4]
  assign _T_1890 = _T_1889 | _T_1427; // @[NV_NVDLA_CSC_dl.scala 708:85:@20517.4]
  assign _T_1891 = _T_1616 & _T_1890; // @[NV_NVDLA_CSC_dl.scala 708:43:@20518.4]
  assign _T_1892 = _T_1616 | _T_1631; // @[NV_NVDLA_CSC_dl.scala 710:38:@20519.4]
  assign _T_1894 = _T_1622 == 2'h0; // @[NV_NVDLA_CSC_dl.scala 710:78:@20520.4]
  assign _T_1895 = _T_1892 & _T_1894; // @[NV_NVDLA_CSC_dl.scala 710:58:@20521.4]
  assign _T_1896 = _T_630 | _T_1895; // @[NV_NVDLA_CSC_dl.scala 710:17:@20522.4]
  assign _T_1899 = _T_1622 == 2'h1; // @[NV_NVDLA_CSC_dl.scala 710:78:@20524.4]
  assign _T_1900 = _T_1892 & _T_1899; // @[NV_NVDLA_CSC_dl.scala 710:58:@20525.4]
  assign _T_1901 = _T_630 | _T_1900; // @[NV_NVDLA_CSC_dl.scala 710:17:@20526.4]
  assign _T_1904 = _T_1622 == 2'h2; // @[NV_NVDLA_CSC_dl.scala 710:78:@20528.4]
  assign _T_1905 = _T_1892 & _T_1904; // @[NV_NVDLA_CSC_dl.scala 710:58:@20529.4]
  assign _T_1906 = _T_630 | _T_1905; // @[NV_NVDLA_CSC_dl.scala 710:17:@20530.4]
  assign _T_1909 = _T_1622 == 2'h3; // @[NV_NVDLA_CSC_dl.scala 710:78:@20532.4]
  assign _T_1910 = _T_1892 & _T_1909; // @[NV_NVDLA_CSC_dl.scala 710:58:@20533.4]
  assign _T_1911 = _T_630 | _T_1910; // @[NV_NVDLA_CSC_dl.scala 710:17:@20534.4]
  assign _GEN_96 = _T_1896 ? _T_1857 : {{2'd0}, _T_1759_0}; // @[NV_NVDLA_CSC_dl.scala 717:35:@20540.4]
  assign _GEN_97 = _T_1901 ? _T_1857 : {{2'd0}, _T_1759_1}; // @[NV_NVDLA_CSC_dl.scala 717:35:@20543.4]
  assign _GEN_98 = _T_1906 ? _T_1857 : {{2'd0}, _T_1759_2}; // @[NV_NVDLA_CSC_dl.scala 717:35:@20546.4]
  assign _GEN_99 = _T_1911 ? _T_1857 : {{2'd0}, _T_1759_3}; // @[NV_NVDLA_CSC_dl.scala 717:35:@20549.4]
  assign _T_1922 = _T_630 | _T_1891; // @[NV_NVDLA_CSC_dl.scala 723:14:@20553.4]
  assign _GEN_100 = _T_1922 ? _T_1857 : _T_1785; // @[NV_NVDLA_CSC_dl.scala 723:34:@20554.4]
  assign _GEN_101 = _T_1335 ? _T_1619 : _T_1794; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  assign _GEN_102 = _T_1335 ? _T_1622 : _T_1797; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  assign _GEN_103 = _T_1335 ? _T_1625 : _T_1800; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  assign _GEN_104 = _T_1335 ? _T_1628 : _T_1803; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  assign _GEN_105 = _T_1335 ? _T_1361 : _T_1806; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  assign _GEN_106 = _T_1335 ? _T_1631 : _T_1809; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  assign _GEN_107 = _T_1335 ? _T_1634 : _T_1812; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  assign _GEN_108 = _T_1335 ? _T_1637 : _T_1815; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  assign _GEN_109 = _T_1335 ? _T_1643 : _T_1818; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  assign _GEN_110 = _T_1335 ? _T_1640 : {{8'd0}, _T_1335}; // @[NV_NVDLA_CSC_dl.scala 730:24:@20561.4]
  assign _T_1932 = {1'h0,_T_1803,_T_1800,_T_1797,_T_1794}; // @[Cat.scala 30:58:@20581.4]
  assign _T_1938 = {_T_1821,_T_1818,_T_1815,_T_1809,_T_1812,_T_1806,_T_1932}; // @[Cat.scala 30:58:@20587.4]
  assign _GEN_111 = _T_1788 ? _T_1938 : _T_1963; // @[NV_NVDLA_CSC_dl.scala 775:33:@20629.4]
  assign _GEN_114 = _T_1943 ? _T_1963 : _T_1966; // @[NV_NVDLA_CSC_dl.scala 775:33:@20638.4]
  assign _GEN_117 = _T_1946 ? _T_1966 : _T_1969; // @[NV_NVDLA_CSC_dl.scala 775:33:@20647.4]
  assign _GEN_120 = _T_1949 ? _T_1969 : _T_1972; // @[NV_NVDLA_CSC_dl.scala 775:33:@20656.4]
  assign _GEN_123 = _T_1952 ? _T_1972 : _T_1975; // @[NV_NVDLA_CSC_dl.scala 775:33:@20665.4]
  assign _GEN_126 = _T_1955 ? _T_1975 : _T_1978; // @[NV_NVDLA_CSC_dl.scala 775:33:@20674.4]
  assign _T_2039 = _T_1978[1:0]; // @[NV_NVDLA_CSC_dl.scala 792:41:@20682.4]
  assign _T_2040 = _T_1978[3:2]; // @[NV_NVDLA_CSC_dl.scala 793:41:@20683.4]
  assign _T_2041 = _T_1978[4]; // @[NV_NVDLA_CSC_dl.scala 794:41:@20684.4]
  assign _T_2042 = _T_1978[5]; // @[NV_NVDLA_CSC_dl.scala 795:42:@20685.4]
  assign _T_2043 = _T_1978[14:7]; // @[NV_NVDLA_CSC_dl.scala 796:41:@20686.4]
  assign _T_2044 = _T_1978[16:15]; // @[NV_NVDLA_CSC_dl.scala 797:45:@20687.4]
  assign _T_2047 = _T_1978[19]; // @[NV_NVDLA_CSC_dl.scala 800:39:@20690.4]
  assign _T_2048 = _T_1978[28:20]; // @[NV_NVDLA_CSC_dl.scala 801:40:@20691.4]
  assign _T_2105 = _T_831[12]; // @[NV_NVDLA_CSC_dl.scala 831:69:@20719.4]
  assign _T_2106 = _T_2105 & io_sc2buf_dat_rd_data_valid; // @[NV_NVDLA_CSC_dl.scala 831:74:@20720.4]
  assign _T_2107 = ~ _T_2051; // @[NV_NVDLA_CSC_dl.scala 831:90:@20721.4]
  assign _T_2108 = _T_2106 & _T_2107; // @[NV_NVDLA_CSC_dl.scala 831:88:@20722.4]
  assign _T_2148 = io_sc2buf_dat_rd_data_valid ? 1'h0 : _T_2051; // @[NV_NVDLA_CSC_dl.scala 846:22:@20756.4]
  assign _T_2162 = io_sc2buf_dat_rd_data_valid ? _T_2051 : _T_2063; // @[NV_NVDLA_CSC_dl.scala 850:48:@20767.4]
  assign _T_2163 = _T_2108 ? 1'h0 : _T_2162; // @[NV_NVDLA_CSC_dl.scala 850:22:@20768.4]
  assign _T_2240 = {_T_2048,_T_2047,_T_2044,_T_2043,1'h0,_T_2042,_T_2041,_T_2040,_T_2039}; // @[Cat.scala 30:58:@20835.4]
  assign _GEN_137 = _T_1958 ? _T_2240 : _T_2222; // @[NV_NVDLA_CSC_dl.scala 889:28:@20838.4]
  assign _GEN_138 = _T_2208 ? _T_2222 : _T_2225; // @[NV_NVDLA_CSC_dl.scala 889:28:@20842.4]
  assign _GEN_139 = _T_2211 ? _T_2225 : _T_2228; // @[NV_NVDLA_CSC_dl.scala 889:28:@20846.4]
  assign _GEN_140 = _T_2214 ? _T_2228 : _T_2231; // @[NV_NVDLA_CSC_dl.scala 889:28:@20850.4]
  assign _T_2269 = _T_2222[4]; // @[NV_NVDLA_CSC_dl.scala 907:39:@20876.4]
  assign _T_2270 = _T_2225[4]; // @[NV_NVDLA_CSC_dl.scala 908:39:@20877.4]
  assign _T_2271 = _T_2228[4]; // @[NV_NVDLA_CSC_dl.scala 909:39:@20878.4]
  assign _T_2272 = _T_2231[4]; // @[NV_NVDLA_CSC_dl.scala 910:39:@20879.4]
  assign _T_2273 = _T_2222[26:18]; // @[NV_NVDLA_CSC_dl.scala 912:38:@20880.4]
  assign _T_2274 = _T_2225[26:18]; // @[NV_NVDLA_CSC_dl.scala 913:38:@20881.4]
  assign _T_2275 = _T_2228[26:18]; // @[NV_NVDLA_CSC_dl.scala 914:38:@20882.4]
  assign _T_2276 = _T_2231[26:18]; // @[NV_NVDLA_CSC_dl.scala 915:38:@20883.4]
  assign _T_2277 = _T_2273[6]; // @[NV_NVDLA_CSC_dl.scala 917:44:@20884.4]
  assign _T_2278 = _T_2274[6]; // @[NV_NVDLA_CSC_dl.scala 918:44:@20885.4]
  assign _T_2279 = _T_2275[6]; // @[NV_NVDLA_CSC_dl.scala 919:44:@20886.4]
  assign _T_2280 = _T_2276[6]; // @[NV_NVDLA_CSC_dl.scala 920:44:@20887.4]
  assign _T_2281 = _T_2268[1:0]; // @[NV_NVDLA_CSC_dl.scala 923:31:@20888.4]
  assign _T_2285 = _T_2268[14:7]; // @[NV_NVDLA_CSC_dl.scala 927:31:@20892.4]
  assign _T_2286 = _T_2268[16:15]; // @[NV_NVDLA_CSC_dl.scala 928:35:@20893.4]
  assign _T_2296 = io_sc2buf_dat_rd_data_valid ? 8'h40 : 8'h0; // @[NV_NVDLA_CSC_dl.scala 939:29:@20902.4]
  assign _T_2307 = _T_960 > 7'h40; // @[NV_NVDLA_CSC_dl.scala 944:50:@20906.4]
  assign _GEN_713 = {{1'd0}, _T_960}; // @[NV_NVDLA_CSC_dl.scala 944:111:@20907.4]
  assign _T_2309 = _T_2182 + _GEN_713; // @[NV_NVDLA_CSC_dl.scala 944:111:@20907.4]
  assign _T_2310 = _T_2182 + _GEN_713; // @[NV_NVDLA_CSC_dl.scala 944:111:@20908.4]
  assign _T_2311 = _T_2310 - _T_2296; // @[NV_NVDLA_CSC_dl.scala 944:133:@20909.4]
  assign _T_2312 = $unsigned(_T_2311); // @[NV_NVDLA_CSC_dl.scala 944:133:@20910.4]
  assign _T_2313 = _T_2312[7:0]; // @[NV_NVDLA_CSC_dl.scala 944:133:@20911.4]
  assign _T_2314 = _T_2307 ? 8'h40 : _T_2313; // @[NV_NVDLA_CSC_dl.scala 944:29:@20912.4]
  assign _T_2318 = _T_2185 + _GEN_713; // @[NV_NVDLA_CSC_dl.scala 945:111:@20914.4]
  assign _T_2319 = _T_2185 + _GEN_713; // @[NV_NVDLA_CSC_dl.scala 945:111:@20915.4]
  assign _T_2320 = _T_2319 - 8'h0; // @[NV_NVDLA_CSC_dl.scala 945:133:@20916.4]
  assign _T_2321 = $unsigned(_T_2320); // @[NV_NVDLA_CSC_dl.scala 945:133:@20917.4]
  assign _T_2322 = _T_2321[7:0]; // @[NV_NVDLA_CSC_dl.scala 945:133:@20918.4]
  assign _T_2323 = _T_2307 ? 8'h40 : _T_2322; // @[NV_NVDLA_CSC_dl.scala 945:29:@20919.4]
  assign _T_2327 = _T_2188 + _GEN_713; // @[NV_NVDLA_CSC_dl.scala 946:111:@20921.4]
  assign _T_2328 = _T_2188 + _GEN_713; // @[NV_NVDLA_CSC_dl.scala 946:111:@20922.4]
  assign _T_2329 = _T_2328 - 8'h0; // @[NV_NVDLA_CSC_dl.scala 946:133:@20923.4]
  assign _T_2330 = $unsigned(_T_2329); // @[NV_NVDLA_CSC_dl.scala 946:133:@20924.4]
  assign _T_2331 = _T_2330[7:0]; // @[NV_NVDLA_CSC_dl.scala 946:133:@20925.4]
  assign _T_2332 = _T_2307 ? 8'h40 : _T_2331; // @[NV_NVDLA_CSC_dl.scala 946:29:@20926.4]
  assign _T_2336 = _T_2191 + _GEN_713; // @[NV_NVDLA_CSC_dl.scala 947:111:@20928.4]
  assign _T_2337 = _T_2191 + _GEN_713; // @[NV_NVDLA_CSC_dl.scala 947:111:@20929.4]
  assign _T_2338 = _T_2337 - 8'h0; // @[NV_NVDLA_CSC_dl.scala 947:133:@20930.4]
  assign _T_2339 = $unsigned(_T_2338); // @[NV_NVDLA_CSC_dl.scala 947:133:@20931.4]
  assign _T_2340 = _T_2339[7:0]; // @[NV_NVDLA_CSC_dl.scala 947:133:@20932.4]
  assign _T_2341 = _T_2307 ? 8'h40 : _T_2340; // @[NV_NVDLA_CSC_dl.scala 947:29:@20933.4]
  assign _T_2343 = ~ _T_2269; // @[NV_NVDLA_CSC_dl.scala 956:52:@20934.4]
  assign _T_2344 = _T_2277 & _T_2343; // @[NV_NVDLA_CSC_dl.scala 956:50:@20935.4]
  assign _T_2345 = _T_2277 & _T_2269; // @[NV_NVDLA_CSC_dl.scala 957:50:@20936.4]
  assign _T_2350 = _T_2345 ? 8'h40 : _T_2314; // @[NV_NVDLA_CSC_dl.scala 957:27:@20939.4]
  assign _T_2351 = _T_2344 ? _T_2194 : _T_2350; // @[NV_NVDLA_CSC_dl.scala 956:27:@20940.4]
  assign _T_2352 = _T_630 ? 8'h40 : _T_2351; // @[NV_NVDLA_CSC_dl.scala 955:27:@20941.4]
  assign _T_2354 = ~ _T_2270; // @[NV_NVDLA_CSC_dl.scala 961:52:@20942.4]
  assign _T_2355 = _T_2278 & _T_2354; // @[NV_NVDLA_CSC_dl.scala 961:50:@20943.4]
  assign _T_2356 = _T_2278 & _T_2270; // @[NV_NVDLA_CSC_dl.scala 962:50:@20944.4]
  assign _T_2361 = _T_2356 ? 8'h40 : _T_2323; // @[NV_NVDLA_CSC_dl.scala 962:27:@20947.4]
  assign _T_2362 = _T_2355 ? _T_2197 : _T_2361; // @[NV_NVDLA_CSC_dl.scala 961:27:@20948.4]
  assign _T_2363 = _T_630 ? 8'h40 : _T_2362; // @[NV_NVDLA_CSC_dl.scala 960:27:@20949.4]
  assign _T_2365 = ~ _T_2271; // @[NV_NVDLA_CSC_dl.scala 966:52:@20950.4]
  assign _T_2366 = _T_2279 & _T_2365; // @[NV_NVDLA_CSC_dl.scala 966:50:@20951.4]
  assign _T_2367 = _T_2279 & _T_2271; // @[NV_NVDLA_CSC_dl.scala 967:50:@20952.4]
  assign _T_2372 = _T_2367 ? 8'h40 : _T_2332; // @[NV_NVDLA_CSC_dl.scala 967:27:@20955.4]
  assign _T_2373 = _T_2366 ? _T_2200 : _T_2372; // @[NV_NVDLA_CSC_dl.scala 966:27:@20956.4]
  assign _T_2374 = _T_630 ? 8'h40 : _T_2373; // @[NV_NVDLA_CSC_dl.scala 965:27:@20957.4]
  assign _T_2376 = ~ _T_2272; // @[NV_NVDLA_CSC_dl.scala 971:52:@20958.4]
  assign _T_2377 = _T_2280 & _T_2376; // @[NV_NVDLA_CSC_dl.scala 971:50:@20959.4]
  assign _T_2378 = _T_2280 & _T_2272; // @[NV_NVDLA_CSC_dl.scala 972:50:@20960.4]
  assign _T_2383 = _T_2378 ? 8'h40 : _T_2341; // @[NV_NVDLA_CSC_dl.scala 972:27:@20963.4]
  assign _T_2384 = _T_2377 ? _T_2203 : _T_2383; // @[NV_NVDLA_CSC_dl.scala 971:27:@20964.4]
  assign _T_2385 = _T_630 ? 8'h40 : _T_2384; // @[NV_NVDLA_CSC_dl.scala 970:27:@20965.4]
  assign _T_2386 = _T_831[17]; // @[NV_NVDLA_CSC_dl.scala 976:46:@20966.4]
  assign _T_2387 = _T_2386 & _T_2208; // @[NV_NVDLA_CSC_dl.scala 976:51:@20967.4]
  assign _T_2388 = _T_630 | _T_2387; // @[NV_NVDLA_CSC_dl.scala 976:34:@20968.4]
  assign _T_2389 = _T_831[18]; // @[NV_NVDLA_CSC_dl.scala 977:46:@20969.4]
  assign _T_2390 = _T_2389 & _T_2211; // @[NV_NVDLA_CSC_dl.scala 977:51:@20970.4]
  assign _T_2392 = _T_884 != 3'h1; // @[NV_NVDLA_CSC_dl.scala 977:87:@20971.4]
  assign _T_2393 = _T_2390 & _T_2392; // @[NV_NVDLA_CSC_dl.scala 977:69:@20972.4]
  assign _T_2394 = _T_630 | _T_2393; // @[NV_NVDLA_CSC_dl.scala 977:34:@20973.4]
  assign _T_2395 = _T_831[19]; // @[NV_NVDLA_CSC_dl.scala 978:46:@20974.4]
  assign _T_2396 = _T_2395 & _T_2214; // @[NV_NVDLA_CSC_dl.scala 978:51:@20975.4]
  assign _T_2398 = _T_884 == 3'h4; // @[NV_NVDLA_CSC_dl.scala 978:87:@20976.4]
  assign _T_2399 = _T_2396 & _T_2398; // @[NV_NVDLA_CSC_dl.scala 978:69:@20977.4]
  assign _T_2400 = _T_630 | _T_2399; // @[NV_NVDLA_CSC_dl.scala 978:34:@20978.4]
  assign _T_2401 = _T_831[20]; // @[NV_NVDLA_CSC_dl.scala 979:46:@20979.4]
  assign _T_2402 = _T_2401 & _T_2217; // @[NV_NVDLA_CSC_dl.scala 979:51:@20980.4]
  assign _T_2405 = _T_2402 & _T_2398; // @[NV_NVDLA_CSC_dl.scala 979:69:@20982.4]
  assign _T_2406 = _T_630 | _T_2405; // @[NV_NVDLA_CSC_dl.scala 979:34:@20983.4]
  assign _T_2407 = _T_831[21]; // @[NV_NVDLA_CSC_dl.scala 981:50:@20984.4]
  assign _T_2408 = _T_2407 & _T_2208; // @[NV_NVDLA_CSC_dl.scala 981:55:@20985.4]
  assign _T_2409 = _T_2408 & _T_2277; // @[NV_NVDLA_CSC_dl.scala 981:73:@20986.4]
  assign _T_2410 = _T_2409 & _T_2269; // @[NV_NVDLA_CSC_dl.scala 981:97:@20987.4]
  assign _T_2411 = _T_630 | _T_2410; // @[NV_NVDLA_CSC_dl.scala 981:38:@20988.4]
  assign _T_2412 = _T_831[22]; // @[NV_NVDLA_CSC_dl.scala 982:50:@20989.4]
  assign _T_2413 = _T_2412 & _T_2211; // @[NV_NVDLA_CSC_dl.scala 982:55:@20990.4]
  assign _T_2414 = _T_2413 & _T_2278; // @[NV_NVDLA_CSC_dl.scala 982:73:@20991.4]
  assign _T_2415 = _T_2414 & _T_2270; // @[NV_NVDLA_CSC_dl.scala 982:97:@20992.4]
  assign _T_2417 = _T_887 != 3'h1; // @[NV_NVDLA_CSC_dl.scala 982:138:@20993.4]
  assign _T_2418 = _T_2415 & _T_2417; // @[NV_NVDLA_CSC_dl.scala 982:120:@20994.4]
  assign _T_2419 = _T_630 | _T_2418; // @[NV_NVDLA_CSC_dl.scala 982:38:@20995.4]
  assign _T_2420 = _T_831[23]; // @[NV_NVDLA_CSC_dl.scala 983:50:@20996.4]
  assign _T_2421 = _T_2420 & _T_2214; // @[NV_NVDLA_CSC_dl.scala 983:55:@20997.4]
  assign _T_2422 = _T_2421 & _T_2279; // @[NV_NVDLA_CSC_dl.scala 983:73:@20998.4]
  assign _T_2423 = _T_2422 & _T_2271; // @[NV_NVDLA_CSC_dl.scala 983:97:@20999.4]
  assign _T_2425 = _T_887 == 3'h4; // @[NV_NVDLA_CSC_dl.scala 983:138:@21000.4]
  assign _T_2426 = _T_2423 & _T_2425; // @[NV_NVDLA_CSC_dl.scala 983:120:@21001.4]
  assign _T_2427 = _T_630 | _T_2426; // @[NV_NVDLA_CSC_dl.scala 983:38:@21002.4]
  assign _T_2428 = _T_831[24]; // @[NV_NVDLA_CSC_dl.scala 984:50:@21003.4]
  assign _T_2429 = _T_2428 & _T_2217; // @[NV_NVDLA_CSC_dl.scala 984:55:@21004.4]
  assign _T_2430 = _T_2429 & _T_2280; // @[NV_NVDLA_CSC_dl.scala 984:73:@21005.4]
  assign _T_2431 = _T_2430 & _T_2272; // @[NV_NVDLA_CSC_dl.scala 984:97:@21006.4]
  assign _T_2434 = _T_2431 & _T_2425; // @[NV_NVDLA_CSC_dl.scala 984:120:@21008.4]
  assign _T_2435 = _T_630 | _T_2434; // @[NV_NVDLA_CSC_dl.scala 984:38:@21009.4]
  assign _GEN_141 = _T_2388 ? _T_2352 : _T_2182; // @[NV_NVDLA_CSC_dl.scala 986:24:@21010.4]
  assign _GEN_142 = _T_2394 ? _T_2363 : _T_2185; // @[NV_NVDLA_CSC_dl.scala 987:24:@21013.4]
  assign _GEN_143 = _T_2400 ? _T_2374 : _T_2188; // @[NV_NVDLA_CSC_dl.scala 988:24:@21016.4]
  assign _GEN_144 = _T_2406 ? _T_2385 : _T_2191; // @[NV_NVDLA_CSC_dl.scala 989:24:@21019.4]
  assign _GEN_145 = _T_2411 ? _T_2352 : _T_2194; // @[NV_NVDLA_CSC_dl.scala 990:28:@21022.4]
  assign _GEN_146 = _T_2419 ? _T_2363 : _T_2197; // @[NV_NVDLA_CSC_dl.scala 991:28:@21025.4]
  assign _GEN_147 = _T_2427 ? _T_2374 : _T_2200; // @[NV_NVDLA_CSC_dl.scala 992:28:@21028.4]
  assign _GEN_148 = _T_2435 ? _T_2385 : _T_2203; // @[NV_NVDLA_CSC_dl.scala 993:28:@21031.4]
  assign _T_2436 = _T_988[7:0]; // @[NV_NVDLA_CSC_dl.scala 1002:55:@21034.4]
  assign _T_2439 = {_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436}; // @[Cat.scala 30:58:@21037.4]
  assign _T_2440 = {_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2439}; // @[Cat.scala 30:58:@21038.4]
  assign _T_2441 = {_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2439,_T_2440}; // @[Cat.scala 30:58:@21039.4]
  assign _T_2442 = {_T_2441,_T_2441}; // @[Cat.scala 30:58:@21040.4]
  assign _T_2443 = _T_2051 ? _T_2442 : _T_2074; // @[NV_NVDLA_CSC_dl.scala 1004:23:@21041.4]
  assign _T_2447 = _T_2063 ? _T_2442 : _T_2082; // @[NV_NVDLA_CSC_dl.scala 1009:23:@21045.4]
  assign _T_2453 = _T_831[26]; // @[NV_NVDLA_CSC_dl.scala 1022:37:@21050.4]
  assign _T_2456 = _T_2285 <= 8'h20; // @[NV_NVDLA_CSC_dl.scala 1023:43:@21051.4]
  assign _T_2457 = _T_2281[0]; // @[NV_NVDLA_CSC_dl.scala 1023:87:@21052.4]
  assign _T_2459 = _T_2457 == 1'h0; // @[NV_NVDLA_CSC_dl.scala 1023:91:@21053.4]
  assign _T_2460 = _T_2456 & _T_2459; // @[NV_NVDLA_CSC_dl.scala 1023:72:@21054.4]
  assign _T_2462 = _T_2443[255:0]; // @[NV_NVDLA_CSC_dl.scala 1023:171:@21055.4]
  assign _T_2463 = {256'h0,_T_2462}; // @[Cat.scala 30:58:@21056.4]
  assign _T_2469 = _T_2456 & _T_2457; // @[NV_NVDLA_CSC_dl.scala 1024:72:@21060.4]
  assign _T_2471 = _T_2443[511:256]; // @[NV_NVDLA_CSC_dl.scala 1024:171:@21061.4]
  assign _T_2472 = {256'h0,_T_2471}; // @[Cat.scala 30:58:@21062.4]
  assign _T_2473 = _T_2469 ? _T_2472 : _T_2443; // @[NV_NVDLA_CSC_dl.scala 1024:27:@21063.4]
  assign _T_2474 = _T_2460 ? _T_2463 : _T_2473; // @[NV_NVDLA_CSC_dl.scala 1023:27:@21064.4]
  assign _T_2475 = _T_2453 ? 512'h0 : _T_2474; // @[NV_NVDLA_CSC_dl.scala 1022:27:@21065.4]
  assign _T_2546 = _T_2475[7:0]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21068.4]
  assign _T_2547 = _T_2475[15:8]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21070.4]
  assign _T_2548 = _T_2475[23:16]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21072.4]
  assign _T_2549 = _T_2475[31:24]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21074.4]
  assign _T_2550 = _T_2475[39:32]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21076.4]
  assign _T_2551 = _T_2475[47:40]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21078.4]
  assign _T_2552 = _T_2475[55:48]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21080.4]
  assign _T_2553 = _T_2475[63:56]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21082.4]
  assign _T_2554 = _T_2475[71:64]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21084.4]
  assign _T_2555 = _T_2475[79:72]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21086.4]
  assign _T_2556 = _T_2475[87:80]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21088.4]
  assign _T_2557 = _T_2475[95:88]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21090.4]
  assign _T_2558 = _T_2475[103:96]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21092.4]
  assign _T_2559 = _T_2475[111:104]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21094.4]
  assign _T_2560 = _T_2475[119:112]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21096.4]
  assign _T_2561 = _T_2475[127:120]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21098.4]
  assign _T_2562 = _T_2475[135:128]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21100.4]
  assign _T_2563 = _T_2475[143:136]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21102.4]
  assign _T_2564 = _T_2475[151:144]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21104.4]
  assign _T_2565 = _T_2475[159:152]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21106.4]
  assign _T_2566 = _T_2475[167:160]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21108.4]
  assign _T_2567 = _T_2475[175:168]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21110.4]
  assign _T_2568 = _T_2475[183:176]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21112.4]
  assign _T_2569 = _T_2475[191:184]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21114.4]
  assign _T_2570 = _T_2475[199:192]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21116.4]
  assign _T_2571 = _T_2475[207:200]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21118.4]
  assign _T_2572 = _T_2475[215:208]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21120.4]
  assign _T_2573 = _T_2475[223:216]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21122.4]
  assign _T_2574 = _T_2475[231:224]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21124.4]
  assign _T_2575 = _T_2475[239:232]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21126.4]
  assign _T_2576 = _T_2475[247:240]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21128.4]
  assign _T_2577 = _T_2475[255:248]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21130.4]
  assign _T_2578 = _T_2475[263:256]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21132.4]
  assign _T_2579 = _T_2475[271:264]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21134.4]
  assign _T_2580 = _T_2475[279:272]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21136.4]
  assign _T_2581 = _T_2475[287:280]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21138.4]
  assign _T_2582 = _T_2475[295:288]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21140.4]
  assign _T_2583 = _T_2475[303:296]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21142.4]
  assign _T_2584 = _T_2475[311:304]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21144.4]
  assign _T_2585 = _T_2475[319:312]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21146.4]
  assign _T_2586 = _T_2475[327:320]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21148.4]
  assign _T_2587 = _T_2475[335:328]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21150.4]
  assign _T_2588 = _T_2475[343:336]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21152.4]
  assign _T_2589 = _T_2475[351:344]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21154.4]
  assign _T_2590 = _T_2475[359:352]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21156.4]
  assign _T_2591 = _T_2475[367:360]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21158.4]
  assign _T_2592 = _T_2475[375:368]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21160.4]
  assign _T_2593 = _T_2475[383:376]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21162.4]
  assign _T_2594 = _T_2475[391:384]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21164.4]
  assign _T_2595 = _T_2475[399:392]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21166.4]
  assign _T_2596 = _T_2475[407:400]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21168.4]
  assign _T_2597 = _T_2475[415:408]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21170.4]
  assign _T_2598 = _T_2475[423:416]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21172.4]
  assign _T_2599 = _T_2475[431:424]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21174.4]
  assign _T_2600 = _T_2475[439:432]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21176.4]
  assign _T_2601 = _T_2475[447:440]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21178.4]
  assign _T_2602 = _T_2475[455:448]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21180.4]
  assign _T_2603 = _T_2475[463:456]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21182.4]
  assign _T_2604 = _T_2475[471:464]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21184.4]
  assign _T_2605 = _T_2475[479:472]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21186.4]
  assign _T_2606 = _T_2475[487:480]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21188.4]
  assign _T_2607 = _T_2475[495:488]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21190.4]
  assign _T_2608 = _T_2475[503:496]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21192.4]
  assign _T_2609 = _T_2475[511:504]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@21194.4]
  assign _T_2622 = _T_831[27]; // @[NV_NVDLA_CSC_dl.scala 1053:39:@21202.4]
  assign _T_2623 = ~ _T_2622; // @[NV_NVDLA_CSC_dl.scala 1053:29:@21203.4]
  assign _T_2625 = {_T_2443,_T_2447}; // @[Cat.scala 30:58:@21204.4]
  assign _T_2626 = _T_2623 ? 1024'h0 : _T_2625; // @[NV_NVDLA_CSC_dl.scala 1053:28:@21205.4]
  assign _T_2627 = _T_831[28]; // @[NV_NVDLA_CSC_dl.scala 1054:39:@21206.4]
  assign _T_2628 = ~ _T_2627; // @[NV_NVDLA_CSC_dl.scala 1054:29:@21207.4]
  assign _T_2630 = {_T_2441,_T_2441,_T_2441,_T_2441}; // @[Cat.scala 30:58:@21208.4]
  assign _T_2631 = _T_2628 ? 1024'h0 : _T_2630; // @[NV_NVDLA_CSC_dl.scala 1054:28:@21209.4]
  assign _T_2632 = _T_831[29]; // @[NV_NVDLA_CSC_dl.scala 1055:39:@21210.4]
  assign _T_2633 = ~ _T_2632; // @[NV_NVDLA_CSC_dl.scala 1055:29:@21211.4]
  assign _T_2636 = _T_2633 ? 1024'h0 : _T_2630; // @[NV_NVDLA_CSC_dl.scala 1055:28:@21213.4]
  assign _T_2637 = _T_831[30]; // @[NV_NVDLA_CSC_dl.scala 1056:39:@21214.4]
  assign _T_2638 = ~ _T_2637; // @[NV_NVDLA_CSC_dl.scala 1056:29:@21215.4]
  assign _T_2641 = _T_2638 ? 1024'h0 : _T_2630; // @[NV_NVDLA_CSC_dl.scala 1056:28:@21217.4]
  assign _T_2643 = {_T_2182,3'h0}; // @[Cat.scala 30:58:@21218.4]
  assign _T_2644 = _T_2626 >> _T_2643; // @[NV_NVDLA_CSC_dl.scala 1058:41:@21219.4]
  assign _T_2645 = _T_2644[511:0]; // @[NV_NVDLA_CSC_dl.scala 1058:82:@21220.4]
  assign _T_2647 = {_T_2185,3'h0}; // @[Cat.scala 30:58:@21221.4]
  assign _T_2648 = _T_2631 >> _T_2647; // @[NV_NVDLA_CSC_dl.scala 1059:41:@21222.4]
  assign _T_2649 = _T_2648[511:0]; // @[NV_NVDLA_CSC_dl.scala 1059:82:@21223.4]
  assign _T_2651 = {_T_2188,3'h0}; // @[Cat.scala 30:58:@21224.4]
  assign _T_2652 = _T_2636 >> _T_2651; // @[NV_NVDLA_CSC_dl.scala 1060:41:@21225.4]
  assign _T_2653 = _T_2652[511:0]; // @[NV_NVDLA_CSC_dl.scala 1060:82:@21226.4]
  assign _T_2655 = {_T_2191,3'h0}; // @[Cat.scala 30:58:@21227.4]
  assign _T_2656 = _T_2641 >> _T_2655; // @[NV_NVDLA_CSC_dl.scala 1061:41:@21228.4]
  assign _T_2657 = _T_2656[511:0]; // @[NV_NVDLA_CSC_dl.scala 1061:82:@21229.4]
  assign _T_2658 = _T_831[32]; // @[NV_NVDLA_CSC_dl.scala 1063:36:@21230.4]
  assign _T_2659 = ~ _T_2658; // @[NV_NVDLA_CSC_dl.scala 1063:26:@21231.4]
  assign _T_2662 = _T_893 == 3'h4; // @[NV_NVDLA_CSC_dl.scala 1064:41:@21232.4]
  assign _T_2663 = _T_2657[127:0]; // @[NV_NVDLA_CSC_dl.scala 1064:81:@21233.4]
  assign _T_2669 = {_T_2663,_T_2621,_T_2619,_T_2615}; // @[Cat.scala 30:58:@21239.4]
  assign _T_2671 = _T_893 == 3'h2; // @[NV_NVDLA_CSC_dl.scala 1065:41:@21240.4]
  assign _T_2672 = _T_2649[255:0]; // @[NV_NVDLA_CSC_dl.scala 1065:81:@21241.4]
  assign _T_2674 = {_T_2672,_T_2611}; // @[Cat.scala 30:58:@21243.4]
  assign _T_2676 = _T_2671 ? _T_2674 : _T_2645; // @[NV_NVDLA_CSC_dl.scala 1065:25:@21245.4]
  assign _T_2677 = _T_2662 ? _T_2669 : _T_2676; // @[NV_NVDLA_CSC_dl.scala 1064:25:@21246.4]
  assign _T_2678 = _T_2659 ? 512'h0 : _T_2677; // @[NV_NVDLA_CSC_dl.scala 1063:25:@21247.4]
  assign _T_2749 = _T_2678[7:0]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21249.4]
  assign _T_2750 = _T_2678[15:8]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21251.4]
  assign _T_2751 = _T_2678[23:16]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21253.4]
  assign _T_2752 = _T_2678[31:24]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21255.4]
  assign _T_2753 = _T_2678[39:32]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21257.4]
  assign _T_2754 = _T_2678[47:40]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21259.4]
  assign _T_2755 = _T_2678[55:48]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21261.4]
  assign _T_2756 = _T_2678[63:56]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21263.4]
  assign _T_2757 = _T_2678[71:64]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21265.4]
  assign _T_2758 = _T_2678[79:72]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21267.4]
  assign _T_2759 = _T_2678[87:80]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21269.4]
  assign _T_2760 = _T_2678[95:88]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21271.4]
  assign _T_2761 = _T_2678[103:96]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21273.4]
  assign _T_2762 = _T_2678[111:104]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21275.4]
  assign _T_2763 = _T_2678[119:112]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21277.4]
  assign _T_2764 = _T_2678[127:120]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21279.4]
  assign _T_2765 = _T_2678[135:128]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21281.4]
  assign _T_2766 = _T_2678[143:136]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21283.4]
  assign _T_2767 = _T_2678[151:144]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21285.4]
  assign _T_2768 = _T_2678[159:152]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21287.4]
  assign _T_2769 = _T_2678[167:160]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21289.4]
  assign _T_2770 = _T_2678[175:168]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21291.4]
  assign _T_2771 = _T_2678[183:176]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21293.4]
  assign _T_2772 = _T_2678[191:184]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21295.4]
  assign _T_2773 = _T_2678[199:192]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21297.4]
  assign _T_2774 = _T_2678[207:200]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21299.4]
  assign _T_2775 = _T_2678[215:208]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21301.4]
  assign _T_2776 = _T_2678[223:216]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21303.4]
  assign _T_2777 = _T_2678[231:224]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21305.4]
  assign _T_2778 = _T_2678[239:232]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21307.4]
  assign _T_2779 = _T_2678[247:240]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21309.4]
  assign _T_2780 = _T_2678[255:248]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21311.4]
  assign _T_2781 = _T_2678[263:256]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21313.4]
  assign _T_2782 = _T_2678[271:264]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21315.4]
  assign _T_2783 = _T_2678[279:272]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21317.4]
  assign _T_2784 = _T_2678[287:280]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21319.4]
  assign _T_2785 = _T_2678[295:288]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21321.4]
  assign _T_2786 = _T_2678[303:296]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21323.4]
  assign _T_2787 = _T_2678[311:304]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21325.4]
  assign _T_2788 = _T_2678[319:312]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21327.4]
  assign _T_2789 = _T_2678[327:320]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21329.4]
  assign _T_2790 = _T_2678[335:328]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21331.4]
  assign _T_2791 = _T_2678[343:336]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21333.4]
  assign _T_2792 = _T_2678[351:344]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21335.4]
  assign _T_2793 = _T_2678[359:352]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21337.4]
  assign _T_2794 = _T_2678[367:360]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21339.4]
  assign _T_2795 = _T_2678[375:368]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21341.4]
  assign _T_2796 = _T_2678[383:376]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21343.4]
  assign _T_2797 = _T_2678[391:384]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21345.4]
  assign _T_2798 = _T_2678[399:392]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21347.4]
  assign _T_2799 = _T_2678[407:400]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21349.4]
  assign _T_2800 = _T_2678[415:408]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21351.4]
  assign _T_2801 = _T_2678[423:416]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21353.4]
  assign _T_2802 = _T_2678[431:424]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21355.4]
  assign _T_2803 = _T_2678[439:432]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21357.4]
  assign _T_2804 = _T_2678[447:440]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21359.4]
  assign _T_2805 = _T_2678[455:448]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21361.4]
  assign _T_2806 = _T_2678[463:456]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21363.4]
  assign _T_2807 = _T_2678[471:464]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21365.4]
  assign _T_2808 = _T_2678[479:472]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21367.4]
  assign _T_2809 = _T_2678[487:480]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21369.4]
  assign _T_2810 = _T_2678[495:488]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21371.4]
  assign _T_2811 = _T_2678[503:496]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21373.4]
  assign _T_2812 = _T_2678[511:504]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@21375.4]
  assign _T_2814 = _T_896 != 3'h1; // @[NV_NVDLA_CSC_dl.scala 1074:59:@21377.4]
  assign _T_2815 = _T_2208 & _T_2814; // @[NV_NVDLA_CSC_dl.scala 1074:41:@21378.4]
  assign _T_2817 = _T_896 == 3'h4; // @[NV_NVDLA_CSC_dl.scala 1075:59:@21379.4]
  assign _T_2818 = _T_2211 & _T_2817; // @[NV_NVDLA_CSC_dl.scala 1075:41:@21380.4]
  assign _T_2821 = _T_2214 & _T_2817; // @[NV_NVDLA_CSC_dl.scala 1076:41:@21382.4]
  assign _GEN_149 = _T_2815 ? _T_2645 : {{256'd0}, _T_2611}; // @[NV_NVDLA_CSC_dl.scala 1078:24:@21383.4]
  assign _GEN_150 = _T_2818 ? _T_2611 : {{128'd0}, _T_2613}; // @[NV_NVDLA_CSC_dl.scala 1081:24:@21386.4]
  assign _GEN_151 = _T_2818 ? _T_2649 : {{384'd0}, _T_2617}; // @[NV_NVDLA_CSC_dl.scala 1081:24:@21386.4]
  assign _GEN_154 = _T_2821 ? _T_2653 : {{384'd0}, _T_2621}; // @[NV_NVDLA_CSC_dl.scala 1085:24:@21390.4]
  assign _T_2827 = 319'hffffffffffffffff << _T_2285; // @[NV_NVDLA_CSC_dl.scala 1094:56:@21396.4]
  assign _T_2828 = _T_2827[63:0]; // @[NV_NVDLA_CSC_dl.scala 1094:73:@21397.4]
  assign _T_2829 = ~ _T_2828; // @[NV_NVDLA_CSC_dl.scala 1094:24:@21398.4]
  assign _T_2831 = _T_2286 >= 2'h1; // @[NV_NVDLA_CSC_dl.scala 1096:51:@21399.4]
  assign _T_2838 = _T_2831 ? 64'hffffffffffffffff : 64'h0; // @[NV_NVDLA_CSC_dl.scala 1096:32:@21401.4]
  assign _T_2840 = _T_2286 >= 2'h2; // @[NV_NVDLA_CSC_dl.scala 1097:51:@21402.4]
  assign _T_2847 = _T_2840 ? 32'hffffffff : 32'h0; // @[NV_NVDLA_CSC_dl.scala 1097:32:@21404.4]
  assign _T_2849 = _T_2286 == 2'h3; // @[NV_NVDLA_CSC_dl.scala 1098:51:@21405.4]
  assign _T_2856 = _T_2849 ? 32'hffffffff : 32'h0; // @[NV_NVDLA_CSC_dl.scala 1098:32:@21407.4]
  assign _T_2857 = _T_2838[31:0]; // @[NV_NVDLA_CSC_dl.scala 1100:57:@21408.4]
  assign _T_2863 = {_T_2857,32'hffffffff}; // @[Cat.scala 30:58:@21410.4]
  assign _T_2864 = _T_2856[15:0]; // @[NV_NVDLA_CSC_dl.scala 1101:57:@21411.4]
  assign _T_2865 = _T_2847[15:0]; // @[NV_NVDLA_CSC_dl.scala 1101:106:@21412.4]
  assign _T_2866 = _T_2838[15:0]; // @[NV_NVDLA_CSC_dl.scala 1101:155:@21413.4]
  assign _T_2874 = {_T_2864,_T_2865,_T_2866,16'hffff}; // @[Cat.scala 30:58:@21417.4]
  assign _T_2876 = _T_902 == 3'h4; // @[NV_NVDLA_CSC_dl.scala 1103:43:@21418.4]
  assign _T_2877 = _T_2829[15:0]; // @[NV_NVDLA_CSC_dl.scala 1103:89:@21419.4]
  assign _T_2879 = {_T_2877,_T_2877,_T_2877,_T_2877}; // @[Cat.scala 30:58:@21421.4]
  assign _T_2880 = _T_2879 & _T_2874; // @[NV_NVDLA_CSC_dl.scala 1103:116:@21422.4]
  assign _T_2882 = _T_902 == 3'h2; // @[NV_NVDLA_CSC_dl.scala 1104:43:@21423.4]
  assign _T_2883 = _T_2829[31:0]; // @[NV_NVDLA_CSC_dl.scala 1104:89:@21424.4]
  assign _T_2884 = {_T_2883,_T_2883}; // @[Cat.scala 30:58:@21425.4]
  assign _T_2885 = _T_2884 & _T_2863; // @[NV_NVDLA_CSC_dl.scala 1104:116:@21426.4]
  assign _T_2886 = _T_2882 ? _T_2885 : _T_2829; // @[NV_NVDLA_CSC_dl.scala 1104:26:@21427.4]
  assign _T_2887 = _T_2876 ? _T_2880 : _T_2886; // @[NV_NVDLA_CSC_dl.scala 1103:26:@21428.4]
  assign _T_2888 = _T_831[33]; // @[NV_NVDLA_CSC_dl.scala 1108:35:@21429.4]
  assign _T_2889_0 = _T_2888 ? _T_2749 : _T_2546; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_1 = _T_2888 ? _T_2750 : _T_2547; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_2 = _T_2888 ? _T_2751 : _T_2548; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_3 = _T_2888 ? _T_2752 : _T_2549; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_4 = _T_2888 ? _T_2753 : _T_2550; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_5 = _T_2888 ? _T_2754 : _T_2551; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_6 = _T_2888 ? _T_2755 : _T_2552; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_7 = _T_2888 ? _T_2756 : _T_2553; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_8 = _T_2888 ? _T_2757 : _T_2554; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_9 = _T_2888 ? _T_2758 : _T_2555; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_10 = _T_2888 ? _T_2759 : _T_2556; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_11 = _T_2888 ? _T_2760 : _T_2557; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_12 = _T_2888 ? _T_2761 : _T_2558; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_13 = _T_2888 ? _T_2762 : _T_2559; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_14 = _T_2888 ? _T_2763 : _T_2560; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_15 = _T_2888 ? _T_2764 : _T_2561; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_16 = _T_2888 ? _T_2765 : _T_2562; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_17 = _T_2888 ? _T_2766 : _T_2563; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_18 = _T_2888 ? _T_2767 : _T_2564; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_19 = _T_2888 ? _T_2768 : _T_2565; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_20 = _T_2888 ? _T_2769 : _T_2566; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_21 = _T_2888 ? _T_2770 : _T_2567; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_22 = _T_2888 ? _T_2771 : _T_2568; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_23 = _T_2888 ? _T_2772 : _T_2569; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_24 = _T_2888 ? _T_2773 : _T_2570; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_25 = _T_2888 ? _T_2774 : _T_2571; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_26 = _T_2888 ? _T_2775 : _T_2572; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_27 = _T_2888 ? _T_2776 : _T_2573; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_28 = _T_2888 ? _T_2777 : _T_2574; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_29 = _T_2888 ? _T_2778 : _T_2575; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_30 = _T_2888 ? _T_2779 : _T_2576; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_31 = _T_2888 ? _T_2780 : _T_2577; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_32 = _T_2888 ? _T_2781 : _T_2578; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_33 = _T_2888 ? _T_2782 : _T_2579; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_34 = _T_2888 ? _T_2783 : _T_2580; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_35 = _T_2888 ? _T_2784 : _T_2581; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_36 = _T_2888 ? _T_2785 : _T_2582; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_37 = _T_2888 ? _T_2786 : _T_2583; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_38 = _T_2888 ? _T_2787 : _T_2584; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_39 = _T_2888 ? _T_2788 : _T_2585; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_40 = _T_2888 ? _T_2789 : _T_2586; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_41 = _T_2888 ? _T_2790 : _T_2587; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_42 = _T_2888 ? _T_2791 : _T_2588; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_43 = _T_2888 ? _T_2792 : _T_2589; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_44 = _T_2888 ? _T_2793 : _T_2590; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_45 = _T_2888 ? _T_2794 : _T_2591; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_46 = _T_2888 ? _T_2795 : _T_2592; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_47 = _T_2888 ? _T_2796 : _T_2593; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_48 = _T_2888 ? _T_2797 : _T_2594; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_49 = _T_2888 ? _T_2798 : _T_2595; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_50 = _T_2888 ? _T_2799 : _T_2596; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_51 = _T_2888 ? _T_2800 : _T_2597; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_52 = _T_2888 ? _T_2801 : _T_2598; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_53 = _T_2888 ? _T_2802 : _T_2599; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_54 = _T_2888 ? _T_2803 : _T_2600; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_55 = _T_2888 ? _T_2804 : _T_2601; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_56 = _T_2888 ? _T_2805 : _T_2602; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_57 = _T_2888 ? _T_2806 : _T_2603; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_58 = _T_2888 ? _T_2807 : _T_2604; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_59 = _T_2888 ? _T_2808 : _T_2605; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_60 = _T_2888 ? _T_2809 : _T_2606; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_61 = _T_2888 ? _T_2810 : _T_2607; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_62 = _T_2888 ? _T_2811 : _T_2608; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_2889_63 = _T_2888 ? _T_2812 : _T_2609; // @[NV_NVDLA_CSC_dl.scala 1108:25:@21430.4]
  assign _T_3022 = _T_2889_0 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21431.4]
  assign _T_3024 = _T_2889_1 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21432.4]
  assign _T_3026 = _T_2889_2 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21433.4]
  assign _T_3028 = _T_2889_3 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21434.4]
  assign _T_3030 = _T_2889_4 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21435.4]
  assign _T_3032 = _T_2889_5 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21436.4]
  assign _T_3034 = _T_2889_6 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21437.4]
  assign _T_3036 = _T_2889_7 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21438.4]
  assign _T_3038 = _T_2889_8 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21439.4]
  assign _T_3040 = _T_2889_9 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21440.4]
  assign _T_3042 = _T_2889_10 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21441.4]
  assign _T_3044 = _T_2889_11 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21442.4]
  assign _T_3046 = _T_2889_12 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21443.4]
  assign _T_3048 = _T_2889_13 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21444.4]
  assign _T_3050 = _T_2889_14 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21445.4]
  assign _T_3052 = _T_2889_15 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21446.4]
  assign _T_3054 = _T_2889_16 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21447.4]
  assign _T_3056 = _T_2889_17 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21448.4]
  assign _T_3058 = _T_2889_18 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21449.4]
  assign _T_3060 = _T_2889_19 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21450.4]
  assign _T_3062 = _T_2889_20 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21451.4]
  assign _T_3064 = _T_2889_21 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21452.4]
  assign _T_3066 = _T_2889_22 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21453.4]
  assign _T_3068 = _T_2889_23 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21454.4]
  assign _T_3070 = _T_2889_24 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21455.4]
  assign _T_3072 = _T_2889_25 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21456.4]
  assign _T_3074 = _T_2889_26 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21457.4]
  assign _T_3076 = _T_2889_27 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21458.4]
  assign _T_3078 = _T_2889_28 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21459.4]
  assign _T_3080 = _T_2889_29 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21460.4]
  assign _T_3082 = _T_2889_30 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21461.4]
  assign _T_3084 = _T_2889_31 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21462.4]
  assign _T_3086 = _T_2889_32 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21463.4]
  assign _T_3088 = _T_2889_33 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21464.4]
  assign _T_3090 = _T_2889_34 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21465.4]
  assign _T_3092 = _T_2889_35 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21466.4]
  assign _T_3094 = _T_2889_36 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21467.4]
  assign _T_3096 = _T_2889_37 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21468.4]
  assign _T_3098 = _T_2889_38 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21469.4]
  assign _T_3100 = _T_2889_39 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21470.4]
  assign _T_3102 = _T_2889_40 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21471.4]
  assign _T_3104 = _T_2889_41 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21472.4]
  assign _T_3106 = _T_2889_42 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21473.4]
  assign _T_3108 = _T_2889_43 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21474.4]
  assign _T_3110 = _T_2889_44 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21475.4]
  assign _T_3112 = _T_2889_45 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21476.4]
  assign _T_3114 = _T_2889_46 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21477.4]
  assign _T_3116 = _T_2889_47 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21478.4]
  assign _T_3118 = _T_2889_48 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21479.4]
  assign _T_3120 = _T_2889_49 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21480.4]
  assign _T_3122 = _T_2889_50 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21481.4]
  assign _T_3124 = _T_2889_51 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21482.4]
  assign _T_3126 = _T_2889_52 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21483.4]
  assign _T_3128 = _T_2889_53 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21484.4]
  assign _T_3130 = _T_2889_54 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21485.4]
  assign _T_3132 = _T_2889_55 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21486.4]
  assign _T_3134 = _T_2889_56 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21487.4]
  assign _T_3136 = _T_2889_57 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21488.4]
  assign _T_3138 = _T_2889_58 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21489.4]
  assign _T_3140 = _T_2889_59 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21490.4]
  assign _T_3142 = _T_2889_60 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21491.4]
  assign _T_3144 = _T_2889_61 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21492.4]
  assign _T_3146 = _T_2889_62 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21493.4]
  assign _T_3148 = _T_2889_63 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@21494.4]
  assign _T_3219 = _T_2887[0]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21560.4]
  assign _T_3220 = _T_3219 & _T_3022; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21561.4]
  assign _T_3221 = _T_2887[1]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21562.4]
  assign _T_3222 = _T_3221 & _T_3024; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21563.4]
  assign _T_3223 = _T_2887[2]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21564.4]
  assign _T_3224 = _T_3223 & _T_3026; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21565.4]
  assign _T_3225 = _T_2887[3]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21566.4]
  assign _T_3226 = _T_3225 & _T_3028; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21567.4]
  assign _T_3227 = _T_2887[4]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21568.4]
  assign _T_3228 = _T_3227 & _T_3030; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21569.4]
  assign _T_3229 = _T_2887[5]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21570.4]
  assign _T_3230 = _T_3229 & _T_3032; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21571.4]
  assign _T_3231 = _T_2887[6]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21572.4]
  assign _T_3232 = _T_3231 & _T_3034; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21573.4]
  assign _T_3233 = _T_2887[7]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21574.4]
  assign _T_3234 = _T_3233 & _T_3036; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21575.4]
  assign _T_3235 = _T_2887[8]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21576.4]
  assign _T_3236 = _T_3235 & _T_3038; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21577.4]
  assign _T_3237 = _T_2887[9]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21578.4]
  assign _T_3238 = _T_3237 & _T_3040; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21579.4]
  assign _T_3239 = _T_2887[10]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21580.4]
  assign _T_3240 = _T_3239 & _T_3042; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21581.4]
  assign _T_3241 = _T_2887[11]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21582.4]
  assign _T_3242 = _T_3241 & _T_3044; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21583.4]
  assign _T_3243 = _T_2887[12]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21584.4]
  assign _T_3244 = _T_3243 & _T_3046; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21585.4]
  assign _T_3245 = _T_2887[13]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21586.4]
  assign _T_3246 = _T_3245 & _T_3048; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21587.4]
  assign _T_3247 = _T_2887[14]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21588.4]
  assign _T_3248 = _T_3247 & _T_3050; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21589.4]
  assign _T_3249 = _T_2887[15]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21590.4]
  assign _T_3250 = _T_3249 & _T_3052; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21591.4]
  assign _T_3251 = _T_2887[16]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21592.4]
  assign _T_3252 = _T_3251 & _T_3054; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21593.4]
  assign _T_3253 = _T_2887[17]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21594.4]
  assign _T_3254 = _T_3253 & _T_3056; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21595.4]
  assign _T_3255 = _T_2887[18]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21596.4]
  assign _T_3256 = _T_3255 & _T_3058; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21597.4]
  assign _T_3257 = _T_2887[19]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21598.4]
  assign _T_3258 = _T_3257 & _T_3060; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21599.4]
  assign _T_3259 = _T_2887[20]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21600.4]
  assign _T_3260 = _T_3259 & _T_3062; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21601.4]
  assign _T_3261 = _T_2887[21]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21602.4]
  assign _T_3262 = _T_3261 & _T_3064; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21603.4]
  assign _T_3263 = _T_2887[22]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21604.4]
  assign _T_3264 = _T_3263 & _T_3066; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21605.4]
  assign _T_3265 = _T_2887[23]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21606.4]
  assign _T_3266 = _T_3265 & _T_3068; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21607.4]
  assign _T_3267 = _T_2887[24]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21608.4]
  assign _T_3268 = _T_3267 & _T_3070; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21609.4]
  assign _T_3269 = _T_2887[25]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21610.4]
  assign _T_3270 = _T_3269 & _T_3072; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21611.4]
  assign _T_3271 = _T_2887[26]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21612.4]
  assign _T_3272 = _T_3271 & _T_3074; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21613.4]
  assign _T_3273 = _T_2887[27]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21614.4]
  assign _T_3274 = _T_3273 & _T_3076; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21615.4]
  assign _T_3275 = _T_2887[28]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21616.4]
  assign _T_3276 = _T_3275 & _T_3078; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21617.4]
  assign _T_3277 = _T_2887[29]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21618.4]
  assign _T_3278 = _T_3277 & _T_3080; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21619.4]
  assign _T_3279 = _T_2887[30]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21620.4]
  assign _T_3280 = _T_3279 & _T_3082; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21621.4]
  assign _T_3281 = _T_2887[31]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21622.4]
  assign _T_3282 = _T_3281 & _T_3084; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21623.4]
  assign _T_3283 = _T_2887[32]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21624.4]
  assign _T_3284 = _T_3283 & _T_3086; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21625.4]
  assign _T_3285 = _T_2887[33]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21626.4]
  assign _T_3286 = _T_3285 & _T_3088; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21627.4]
  assign _T_3287 = _T_2887[34]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21628.4]
  assign _T_3288 = _T_3287 & _T_3090; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21629.4]
  assign _T_3289 = _T_2887[35]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21630.4]
  assign _T_3290 = _T_3289 & _T_3092; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21631.4]
  assign _T_3291 = _T_2887[36]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21632.4]
  assign _T_3292 = _T_3291 & _T_3094; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21633.4]
  assign _T_3293 = _T_2887[37]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21634.4]
  assign _T_3294 = _T_3293 & _T_3096; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21635.4]
  assign _T_3295 = _T_2887[38]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21636.4]
  assign _T_3296 = _T_3295 & _T_3098; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21637.4]
  assign _T_3297 = _T_2887[39]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21638.4]
  assign _T_3298 = _T_3297 & _T_3100; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21639.4]
  assign _T_3299 = _T_2887[40]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21640.4]
  assign _T_3300 = _T_3299 & _T_3102; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21641.4]
  assign _T_3301 = _T_2887[41]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21642.4]
  assign _T_3302 = _T_3301 & _T_3104; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21643.4]
  assign _T_3303 = _T_2887[42]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21644.4]
  assign _T_3304 = _T_3303 & _T_3106; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21645.4]
  assign _T_3305 = _T_2887[43]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21646.4]
  assign _T_3306 = _T_3305 & _T_3108; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21647.4]
  assign _T_3307 = _T_2887[44]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21648.4]
  assign _T_3308 = _T_3307 & _T_3110; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21649.4]
  assign _T_3309 = _T_2887[45]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21650.4]
  assign _T_3310 = _T_3309 & _T_3112; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21651.4]
  assign _T_3311 = _T_2887[46]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21652.4]
  assign _T_3312 = _T_3311 & _T_3114; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21653.4]
  assign _T_3313 = _T_2887[47]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21654.4]
  assign _T_3314 = _T_3313 & _T_3116; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21655.4]
  assign _T_3315 = _T_2887[48]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21656.4]
  assign _T_3316 = _T_3315 & _T_3118; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21657.4]
  assign _T_3317 = _T_2887[49]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21658.4]
  assign _T_3318 = _T_3317 & _T_3120; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21659.4]
  assign _T_3319 = _T_2887[50]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21660.4]
  assign _T_3320 = _T_3319 & _T_3122; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21661.4]
  assign _T_3321 = _T_2887[51]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21662.4]
  assign _T_3322 = _T_3321 & _T_3124; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21663.4]
  assign _T_3323 = _T_2887[52]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21664.4]
  assign _T_3324 = _T_3323 & _T_3126; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21665.4]
  assign _T_3325 = _T_2887[53]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21666.4]
  assign _T_3326 = _T_3325 & _T_3128; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21667.4]
  assign _T_3327 = _T_2887[54]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21668.4]
  assign _T_3328 = _T_3327 & _T_3130; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21669.4]
  assign _T_3329 = _T_2887[55]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21670.4]
  assign _T_3330 = _T_3329 & _T_3132; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21671.4]
  assign _T_3331 = _T_2887[56]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21672.4]
  assign _T_3332 = _T_3331 & _T_3134; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21673.4]
  assign _T_3333 = _T_2887[57]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21674.4]
  assign _T_3334 = _T_3333 & _T_3136; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21675.4]
  assign _T_3335 = _T_2887[58]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21676.4]
  assign _T_3336 = _T_3335 & _T_3138; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21677.4]
  assign _T_3337 = _T_2887[59]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21678.4]
  assign _T_3338 = _T_3337 & _T_3140; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21679.4]
  assign _T_3339 = _T_2887[60]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21680.4]
  assign _T_3340 = _T_3339 & _T_3142; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21681.4]
  assign _T_3341 = _T_2887[61]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21682.4]
  assign _T_3342 = _T_3341 & _T_3144; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21683.4]
  assign _T_3343 = _T_2887[62]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21684.4]
  assign _T_3344 = _T_3343 & _T_3146; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21685.4]
  assign _T_3345 = _T_2887[63]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@21686.4]
  assign _T_3346 = _T_3345 & _T_3148; // @[NV_NVDLA_CSC_dl.scala 1110:83:@21687.4]
  assign _GEN_156 = _T_2248 ? _T_3220 : _T_3689_0; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_157 = _T_2248 ? _T_3222 : _T_3689_1; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_158 = _T_2248 ? _T_3224 : _T_3689_2; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_159 = _T_2248 ? _T_3226 : _T_3689_3; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_160 = _T_2248 ? _T_3228 : _T_3689_4; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_161 = _T_2248 ? _T_3230 : _T_3689_5; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_162 = _T_2248 ? _T_3232 : _T_3689_6; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_163 = _T_2248 ? _T_3234 : _T_3689_7; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_164 = _T_2248 ? _T_3236 : _T_3689_8; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_165 = _T_2248 ? _T_3238 : _T_3689_9; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_166 = _T_2248 ? _T_3240 : _T_3689_10; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_167 = _T_2248 ? _T_3242 : _T_3689_11; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_168 = _T_2248 ? _T_3244 : _T_3689_12; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_169 = _T_2248 ? _T_3246 : _T_3689_13; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_170 = _T_2248 ? _T_3248 : _T_3689_14; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_171 = _T_2248 ? _T_3250 : _T_3689_15; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_172 = _T_2248 ? _T_3252 : _T_3689_16; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_173 = _T_2248 ? _T_3254 : _T_3689_17; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_174 = _T_2248 ? _T_3256 : _T_3689_18; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_175 = _T_2248 ? _T_3258 : _T_3689_19; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_176 = _T_2248 ? _T_3260 : _T_3689_20; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_177 = _T_2248 ? _T_3262 : _T_3689_21; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_178 = _T_2248 ? _T_3264 : _T_3689_22; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_179 = _T_2248 ? _T_3266 : _T_3689_23; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_180 = _T_2248 ? _T_3268 : _T_3689_24; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_181 = _T_2248 ? _T_3270 : _T_3689_25; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_182 = _T_2248 ? _T_3272 : _T_3689_26; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_183 = _T_2248 ? _T_3274 : _T_3689_27; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_184 = _T_2248 ? _T_3276 : _T_3689_28; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_185 = _T_2248 ? _T_3278 : _T_3689_29; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_186 = _T_2248 ? _T_3280 : _T_3689_30; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_187 = _T_2248 ? _T_3282 : _T_3689_31; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_188 = _T_2248 ? _T_3284 : _T_3689_32; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_189 = _T_2248 ? _T_3286 : _T_3689_33; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_190 = _T_2248 ? _T_3288 : _T_3689_34; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_191 = _T_2248 ? _T_3290 : _T_3689_35; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_192 = _T_2248 ? _T_3292 : _T_3689_36; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_193 = _T_2248 ? _T_3294 : _T_3689_37; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_194 = _T_2248 ? _T_3296 : _T_3689_38; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_195 = _T_2248 ? _T_3298 : _T_3689_39; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_196 = _T_2248 ? _T_3300 : _T_3689_40; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_197 = _T_2248 ? _T_3302 : _T_3689_41; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_198 = _T_2248 ? _T_3304 : _T_3689_42; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_199 = _T_2248 ? _T_3306 : _T_3689_43; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_200 = _T_2248 ? _T_3308 : _T_3689_44; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_201 = _T_2248 ? _T_3310 : _T_3689_45; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_202 = _T_2248 ? _T_3312 : _T_3689_46; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_203 = _T_2248 ? _T_3314 : _T_3689_47; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_204 = _T_2248 ? _T_3316 : _T_3689_48; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_205 = _T_2248 ? _T_3318 : _T_3689_49; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_206 = _T_2248 ? _T_3320 : _T_3689_50; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_207 = _T_2248 ? _T_3322 : _T_3689_51; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_208 = _T_2248 ? _T_3324 : _T_3689_52; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_209 = _T_2248 ? _T_3326 : _T_3689_53; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_210 = _T_2248 ? _T_3328 : _T_3689_54; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_211 = _T_2248 ? _T_3330 : _T_3689_55; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_212 = _T_2248 ? _T_3332 : _T_3689_56; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_213 = _T_2248 ? _T_3334 : _T_3689_57; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_214 = _T_2248 ? _T_3336 : _T_3689_58; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_215 = _T_2248 ? _T_3338 : _T_3689_59; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_216 = _T_2248 ? _T_3340 : _T_3689_60; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_217 = _T_2248 ? _T_3342 : _T_3689_61; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_218 = _T_2248 ? _T_3344 : _T_3689_62; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _GEN_219 = _T_2248 ? _T_3346 : _T_3689_63; // @[NV_NVDLA_CSC_dl.scala 1133:30:@21826.4]
  assign _T_3956 = _T_2248 & _T_3220; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21892.4]
  assign _T_3957 = _T_2248 & _T_3222; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21896.4]
  assign _T_3958 = _T_2248 & _T_3224; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21900.4]
  assign _T_3959 = _T_2248 & _T_3226; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21904.4]
  assign _T_3960 = _T_2248 & _T_3228; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21908.4]
  assign _T_3961 = _T_2248 & _T_3230; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21912.4]
  assign _T_3962 = _T_2248 & _T_3232; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21916.4]
  assign _T_3963 = _T_2248 & _T_3234; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21920.4]
  assign _T_3964 = _T_2248 & _T_3236; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21924.4]
  assign _T_3965 = _T_2248 & _T_3238; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21928.4]
  assign _T_3966 = _T_2248 & _T_3240; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21932.4]
  assign _T_3967 = _T_2248 & _T_3242; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21936.4]
  assign _T_3968 = _T_2248 & _T_3244; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21940.4]
  assign _T_3969 = _T_2248 & _T_3246; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21944.4]
  assign _T_3970 = _T_2248 & _T_3248; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21948.4]
  assign _T_3971 = _T_2248 & _T_3250; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21952.4]
  assign _T_3972 = _T_2248 & _T_3252; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21956.4]
  assign _T_3973 = _T_2248 & _T_3254; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21960.4]
  assign _T_3974 = _T_2248 & _T_3256; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21964.4]
  assign _T_3975 = _T_2248 & _T_3258; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21968.4]
  assign _T_3976 = _T_2248 & _T_3260; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21972.4]
  assign _T_3977 = _T_2248 & _T_3262; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21976.4]
  assign _T_3978 = _T_2248 & _T_3264; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21980.4]
  assign _T_3979 = _T_2248 & _T_3266; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21984.4]
  assign _T_3980 = _T_2248 & _T_3268; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21988.4]
  assign _T_3981 = _T_2248 & _T_3270; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21992.4]
  assign _T_3982 = _T_2248 & _T_3272; // @[NV_NVDLA_CSC_dl.scala 1137:34:@21996.4]
  assign _T_3983 = _T_2248 & _T_3274; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22000.4]
  assign _T_3984 = _T_2248 & _T_3276; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22004.4]
  assign _T_3985 = _T_2248 & _T_3278; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22008.4]
  assign _T_3986 = _T_2248 & _T_3280; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22012.4]
  assign _T_3987 = _T_2248 & _T_3282; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22016.4]
  assign _T_3988 = _T_2248 & _T_3284; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22020.4]
  assign _T_3989 = _T_2248 & _T_3286; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22024.4]
  assign _T_3990 = _T_2248 & _T_3288; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22028.4]
  assign _T_3991 = _T_2248 & _T_3290; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22032.4]
  assign _T_3992 = _T_2248 & _T_3292; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22036.4]
  assign _T_3993 = _T_2248 & _T_3294; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22040.4]
  assign _T_3994 = _T_2248 & _T_3296; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22044.4]
  assign _T_3995 = _T_2248 & _T_3298; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22048.4]
  assign _T_3996 = _T_2248 & _T_3300; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22052.4]
  assign _T_3997 = _T_2248 & _T_3302; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22056.4]
  assign _T_3998 = _T_2248 & _T_3304; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22060.4]
  assign _T_3999 = _T_2248 & _T_3306; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22064.4]
  assign _T_4000 = _T_2248 & _T_3308; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22068.4]
  assign _T_4001 = _T_2248 & _T_3310; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22072.4]
  assign _T_4002 = _T_2248 & _T_3312; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22076.4]
  assign _T_4003 = _T_2248 & _T_3314; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22080.4]
  assign _T_4004 = _T_2248 & _T_3316; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22084.4]
  assign _T_4005 = _T_2248 & _T_3318; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22088.4]
  assign _T_4006 = _T_2248 & _T_3320; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22092.4]
  assign _T_4007 = _T_2248 & _T_3322; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22096.4]
  assign _T_4008 = _T_2248 & _T_3324; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22100.4]
  assign _T_4009 = _T_2248 & _T_3326; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22104.4]
  assign _T_4010 = _T_2248 & _T_3328; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22108.4]
  assign _T_4011 = _T_2248 & _T_3330; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22112.4]
  assign _T_4012 = _T_2248 & _T_3332; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22116.4]
  assign _T_4013 = _T_2248 & _T_3334; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22120.4]
  assign _T_4014 = _T_2248 & _T_3336; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22124.4]
  assign _T_4015 = _T_2248 & _T_3338; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22128.4]
  assign _T_4016 = _T_2248 & _T_3340; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22132.4]
  assign _T_4017 = _T_2248 & _T_3342; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22136.4]
  assign _T_4018 = _T_2248 & _T_3344; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22140.4]
  assign _T_4019 = _T_2248 & _T_3346; // @[NV_NVDLA_CSC_dl.scala 1137:34:@22144.4]
  assign _T_4559 = ~ _T_3419; // @[NV_NVDLA_CSC_dl.scala 1151:24:@22217.4]
  assign _T_4694_0 = _T_4559 ? 1'h0 : _T_3689_0; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_1 = _T_4559 ? 1'h0 : _T_3689_1; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_2 = _T_4559 ? 1'h0 : _T_3689_2; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_3 = _T_4559 ? 1'h0 : _T_3689_3; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_4 = _T_4559 ? 1'h0 : _T_3689_4; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_5 = _T_4559 ? 1'h0 : _T_3689_5; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_6 = _T_4559 ? 1'h0 : _T_3689_6; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_7 = _T_4559 ? 1'h0 : _T_3689_7; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_8 = _T_4559 ? 1'h0 : _T_3689_8; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_9 = _T_4559 ? 1'h0 : _T_3689_9; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_10 = _T_4559 ? 1'h0 : _T_3689_10; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_11 = _T_4559 ? 1'h0 : _T_3689_11; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_12 = _T_4559 ? 1'h0 : _T_3689_12; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_13 = _T_4559 ? 1'h0 : _T_3689_13; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_14 = _T_4559 ? 1'h0 : _T_3689_14; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_15 = _T_4559 ? 1'h0 : _T_3689_15; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_16 = _T_4559 ? 1'h0 : _T_3689_16; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_17 = _T_4559 ? 1'h0 : _T_3689_17; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_18 = _T_4559 ? 1'h0 : _T_3689_18; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_19 = _T_4559 ? 1'h0 : _T_3689_19; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_20 = _T_4559 ? 1'h0 : _T_3689_20; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_21 = _T_4559 ? 1'h0 : _T_3689_21; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_22 = _T_4559 ? 1'h0 : _T_3689_22; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_23 = _T_4559 ? 1'h0 : _T_3689_23; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_24 = _T_4559 ? 1'h0 : _T_3689_24; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_25 = _T_4559 ? 1'h0 : _T_3689_25; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_26 = _T_4559 ? 1'h0 : _T_3689_26; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_27 = _T_4559 ? 1'h0 : _T_3689_27; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_28 = _T_4559 ? 1'h0 : _T_3689_28; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_29 = _T_4559 ? 1'h0 : _T_3689_29; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_30 = _T_4559 ? 1'h0 : _T_3689_30; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_31 = _T_4559 ? 1'h0 : _T_3689_31; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_32 = _T_4559 ? 1'h0 : _T_3689_32; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_33 = _T_4559 ? 1'h0 : _T_3689_33; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_34 = _T_4559 ? 1'h0 : _T_3689_34; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_35 = _T_4559 ? 1'h0 : _T_3689_35; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_36 = _T_4559 ? 1'h0 : _T_3689_36; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_37 = _T_4559 ? 1'h0 : _T_3689_37; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_38 = _T_4559 ? 1'h0 : _T_3689_38; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_39 = _T_4559 ? 1'h0 : _T_3689_39; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_40 = _T_4559 ? 1'h0 : _T_3689_40; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_41 = _T_4559 ? 1'h0 : _T_3689_41; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_42 = _T_4559 ? 1'h0 : _T_3689_42; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_43 = _T_4559 ? 1'h0 : _T_3689_43; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_44 = _T_4559 ? 1'h0 : _T_3689_44; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_45 = _T_4559 ? 1'h0 : _T_3689_45; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_46 = _T_4559 ? 1'h0 : _T_3689_46; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_47 = _T_4559 ? 1'h0 : _T_3689_47; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_48 = _T_4559 ? 1'h0 : _T_3689_48; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_49 = _T_4559 ? 1'h0 : _T_3689_49; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_50 = _T_4559 ? 1'h0 : _T_3689_50; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_51 = _T_4559 ? 1'h0 : _T_3689_51; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_52 = _T_4559 ? 1'h0 : _T_3689_52; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_53 = _T_4559 ? 1'h0 : _T_3689_53; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_54 = _T_4559 ? 1'h0 : _T_3689_54; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_55 = _T_4559 ? 1'h0 : _T_3689_55; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_56 = _T_4559 ? 1'h0 : _T_3689_56; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_57 = _T_4559 ? 1'h0 : _T_3689_57; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_58 = _T_4559 ? 1'h0 : _T_3689_58; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_59 = _T_4559 ? 1'h0 : _T_3689_59; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_60 = _T_4559 ? 1'h0 : _T_3689_60; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_61 = _T_4559 ? 1'h0 : _T_3689_61; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_62 = _T_4559 ? 1'h0 : _T_3689_62; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4694_63 = _T_4559 ? 1'h0 : _T_3689_63; // @[NV_NVDLA_CSC_dl.scala 1151:23:@22283.4]
  assign _T_4826 = _T_3419 | _T_4022; // @[NV_NVDLA_CSC_dl.scala 1155:19:@22285.4]
  assign _GEN_284 = _T_4826 ? _T_4694_0 : _T_4289_0; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_285 = _T_4826 ? _T_4694_1 : _T_4289_1; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_286 = _T_4826 ? _T_4694_2 : _T_4289_2; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_287 = _T_4826 ? _T_4694_3 : _T_4289_3; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_288 = _T_4826 ? _T_4694_4 : _T_4289_4; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_289 = _T_4826 ? _T_4694_5 : _T_4289_5; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_290 = _T_4826 ? _T_4694_6 : _T_4289_6; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_291 = _T_4826 ? _T_4694_7 : _T_4289_7; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_292 = _T_4826 ? _T_4694_8 : _T_4289_8; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_293 = _T_4826 ? _T_4694_9 : _T_4289_9; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_294 = _T_4826 ? _T_4694_10 : _T_4289_10; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_295 = _T_4826 ? _T_4694_11 : _T_4289_11; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_296 = _T_4826 ? _T_4694_12 : _T_4289_12; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_297 = _T_4826 ? _T_4694_13 : _T_4289_13; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_298 = _T_4826 ? _T_4694_14 : _T_4289_14; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_299 = _T_4826 ? _T_4694_15 : _T_4289_15; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_300 = _T_4826 ? _T_4694_16 : _T_4289_16; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_301 = _T_4826 ? _T_4694_17 : _T_4289_17; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_302 = _T_4826 ? _T_4694_18 : _T_4289_18; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_303 = _T_4826 ? _T_4694_19 : _T_4289_19; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_304 = _T_4826 ? _T_4694_20 : _T_4289_20; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_305 = _T_4826 ? _T_4694_21 : _T_4289_21; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_306 = _T_4826 ? _T_4694_22 : _T_4289_22; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_307 = _T_4826 ? _T_4694_23 : _T_4289_23; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_308 = _T_4826 ? _T_4694_24 : _T_4289_24; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_309 = _T_4826 ? _T_4694_25 : _T_4289_25; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_310 = _T_4826 ? _T_4694_26 : _T_4289_26; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_311 = _T_4826 ? _T_4694_27 : _T_4289_27; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_312 = _T_4826 ? _T_4694_28 : _T_4289_28; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_313 = _T_4826 ? _T_4694_29 : _T_4289_29; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_314 = _T_4826 ? _T_4694_30 : _T_4289_30; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_315 = _T_4826 ? _T_4694_31 : _T_4289_31; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_316 = _T_4826 ? _T_4694_32 : _T_4289_32; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_317 = _T_4826 ? _T_4694_33 : _T_4289_33; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_318 = _T_4826 ? _T_4694_34 : _T_4289_34; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_319 = _T_4826 ? _T_4694_35 : _T_4289_35; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_320 = _T_4826 ? _T_4694_36 : _T_4289_36; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_321 = _T_4826 ? _T_4694_37 : _T_4289_37; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_322 = _T_4826 ? _T_4694_38 : _T_4289_38; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_323 = _T_4826 ? _T_4694_39 : _T_4289_39; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_324 = _T_4826 ? _T_4694_40 : _T_4289_40; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_325 = _T_4826 ? _T_4694_41 : _T_4289_41; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_326 = _T_4826 ? _T_4694_42 : _T_4289_42; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_327 = _T_4826 ? _T_4694_43 : _T_4289_43; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_328 = _T_4826 ? _T_4694_44 : _T_4289_44; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_329 = _T_4826 ? _T_4694_45 : _T_4289_45; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_330 = _T_4826 ? _T_4694_46 : _T_4289_46; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_331 = _T_4826 ? _T_4694_47 : _T_4289_47; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_332 = _T_4826 ? _T_4694_48 : _T_4289_48; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_333 = _T_4826 ? _T_4694_49 : _T_4289_49; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_334 = _T_4826 ? _T_4694_50 : _T_4289_50; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_335 = _T_4826 ? _T_4694_51 : _T_4289_51; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_336 = _T_4826 ? _T_4694_52 : _T_4289_52; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_337 = _T_4826 ? _T_4694_53 : _T_4289_53; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_338 = _T_4826 ? _T_4694_54 : _T_4289_54; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_339 = _T_4826 ? _T_4694_55 : _T_4289_55; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_340 = _T_4826 ? _T_4694_56 : _T_4289_56; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_341 = _T_4826 ? _T_4694_57 : _T_4289_57; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_342 = _T_4826 ? _T_4694_58 : _T_4289_58; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_343 = _T_4826 ? _T_4694_59 : _T_4289_59; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_344 = _T_4826 ? _T_4694_60 : _T_4289_60; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_345 = _T_4826 ? _T_4694_61 : _T_4289_61; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_346 = _T_4826 ? _T_4694_62 : _T_4289_62; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_347 = _T_4826 ? _T_4694_63 : _T_4289_63; // @[NV_NVDLA_CSC_dl.scala 1155:33:@22286.4]
  assign _GEN_348 = _T_3419 ? {{8'd0}, _T_3419} : _T_4488; // @[NV_NVDLA_CSC_dl.scala 1158:19:@22352.4]
  assign _T_4830 = ~ _T_4022; // @[NV_NVDLA_CSC_dl.scala 1172:27:@22549.4]
  assign _T_4832 = _T_4830 ? 9'h0 : _T_4488; // @[NV_NVDLA_CSC_dl.scala 1172:26:@22550.4]
  assign _T_4840 = _T_4022 | _T_4829; // @[NV_NVDLA_CSC_dl.scala 1176:85:@22557.4]
  assign _GEN_413 = _T_4840 ? _T_4832 : _T_4842; // @[Reg.scala 20:19:@22559.4]
  assign _GEN_414 = _T_4840 ? _T_4832 : _T_4846; // @[Reg.scala 20:19:@22565.4]
  assign _GEN_415 = _T_4840 ? _T_4289_0 : _T_5114_0; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_416 = _T_4840 ? _T_4289_1 : _T_5114_1; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_417 = _T_4840 ? _T_4289_2 : _T_5114_2; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_418 = _T_4840 ? _T_4289_3 : _T_5114_3; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_419 = _T_4840 ? _T_4289_4 : _T_5114_4; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_420 = _T_4840 ? _T_4289_5 : _T_5114_5; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_421 = _T_4840 ? _T_4289_6 : _T_5114_6; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_422 = _T_4840 ? _T_4289_7 : _T_5114_7; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_423 = _T_4840 ? _T_4289_8 : _T_5114_8; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_424 = _T_4840 ? _T_4289_9 : _T_5114_9; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_425 = _T_4840 ? _T_4289_10 : _T_5114_10; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_426 = _T_4840 ? _T_4289_11 : _T_5114_11; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_427 = _T_4840 ? _T_4289_12 : _T_5114_12; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_428 = _T_4840 ? _T_4289_13 : _T_5114_13; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_429 = _T_4840 ? _T_4289_14 : _T_5114_14; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_430 = _T_4840 ? _T_4289_15 : _T_5114_15; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_431 = _T_4840 ? _T_4289_16 : _T_5114_16; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_432 = _T_4840 ? _T_4289_17 : _T_5114_17; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_433 = _T_4840 ? _T_4289_18 : _T_5114_18; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_434 = _T_4840 ? _T_4289_19 : _T_5114_19; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_435 = _T_4840 ? _T_4289_20 : _T_5114_20; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_436 = _T_4840 ? _T_4289_21 : _T_5114_21; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_437 = _T_4840 ? _T_4289_22 : _T_5114_22; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_438 = _T_4840 ? _T_4289_23 : _T_5114_23; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_439 = _T_4840 ? _T_4289_24 : _T_5114_24; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_440 = _T_4840 ? _T_4289_25 : _T_5114_25; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_441 = _T_4840 ? _T_4289_26 : _T_5114_26; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_442 = _T_4840 ? _T_4289_27 : _T_5114_27; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_443 = _T_4840 ? _T_4289_28 : _T_5114_28; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_444 = _T_4840 ? _T_4289_29 : _T_5114_29; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_445 = _T_4840 ? _T_4289_30 : _T_5114_30; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_446 = _T_4840 ? _T_4289_31 : _T_5114_31; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_447 = _T_4840 ? _T_4289_32 : _T_5114_32; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_448 = _T_4840 ? _T_4289_33 : _T_5114_33; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_449 = _T_4840 ? _T_4289_34 : _T_5114_34; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_450 = _T_4840 ? _T_4289_35 : _T_5114_35; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_451 = _T_4840 ? _T_4289_36 : _T_5114_36; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_452 = _T_4840 ? _T_4289_37 : _T_5114_37; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_453 = _T_4840 ? _T_4289_38 : _T_5114_38; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_454 = _T_4840 ? _T_4289_39 : _T_5114_39; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_455 = _T_4840 ? _T_4289_40 : _T_5114_40; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_456 = _T_4840 ? _T_4289_41 : _T_5114_41; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_457 = _T_4840 ? _T_4289_42 : _T_5114_42; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_458 = _T_4840 ? _T_4289_43 : _T_5114_43; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_459 = _T_4840 ? _T_4289_44 : _T_5114_44; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_460 = _T_4840 ? _T_4289_45 : _T_5114_45; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_461 = _T_4840 ? _T_4289_46 : _T_5114_46; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_462 = _T_4840 ? _T_4289_47 : _T_5114_47; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_463 = _T_4840 ? _T_4289_48 : _T_5114_48; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_464 = _T_4840 ? _T_4289_49 : _T_5114_49; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_465 = _T_4840 ? _T_4289_50 : _T_5114_50; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_466 = _T_4840 ? _T_4289_51 : _T_5114_51; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_467 = _T_4840 ? _T_4289_52 : _T_5114_52; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_468 = _T_4840 ? _T_4289_53 : _T_5114_53; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_469 = _T_4840 ? _T_4289_54 : _T_5114_54; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_470 = _T_4840 ? _T_4289_55 : _T_5114_55; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_471 = _T_4840 ? _T_4289_56 : _T_5114_56; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_472 = _T_4840 ? _T_4289_57 : _T_5114_57; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_473 = _T_4840 ? _T_4289_58 : _T_5114_58; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_474 = _T_4840 ? _T_4289_59 : _T_5114_59; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_475 = _T_4840 ? _T_4289_60 : _T_5114_60; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_476 = _T_4840 ? _T_4289_61 : _T_5114_61; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_477 = _T_4840 ? _T_4289_62 : _T_5114_62; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_478 = _T_4840 ? _T_4289_63 : _T_5114_63; // @[Reg.scala 20:19:@22636.4]
  assign _GEN_479 = _T_4840 ? _T_4289_0 : _T_5578_0; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_480 = _T_4840 ? _T_4289_1 : _T_5578_1; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_481 = _T_4840 ? _T_4289_2 : _T_5578_2; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_482 = _T_4840 ? _T_4289_3 : _T_5578_3; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_483 = _T_4840 ? _T_4289_4 : _T_5578_4; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_484 = _T_4840 ? _T_4289_5 : _T_5578_5; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_485 = _T_4840 ? _T_4289_6 : _T_5578_6; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_486 = _T_4840 ? _T_4289_7 : _T_5578_7; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_487 = _T_4840 ? _T_4289_8 : _T_5578_8; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_488 = _T_4840 ? _T_4289_9 : _T_5578_9; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_489 = _T_4840 ? _T_4289_10 : _T_5578_10; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_490 = _T_4840 ? _T_4289_11 : _T_5578_11; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_491 = _T_4840 ? _T_4289_12 : _T_5578_12; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_492 = _T_4840 ? _T_4289_13 : _T_5578_13; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_493 = _T_4840 ? _T_4289_14 : _T_5578_14; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_494 = _T_4840 ? _T_4289_15 : _T_5578_15; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_495 = _T_4840 ? _T_4289_16 : _T_5578_16; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_496 = _T_4840 ? _T_4289_17 : _T_5578_17; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_497 = _T_4840 ? _T_4289_18 : _T_5578_18; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_498 = _T_4840 ? _T_4289_19 : _T_5578_19; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_499 = _T_4840 ? _T_4289_20 : _T_5578_20; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_500 = _T_4840 ? _T_4289_21 : _T_5578_21; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_501 = _T_4840 ? _T_4289_22 : _T_5578_22; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_502 = _T_4840 ? _T_4289_23 : _T_5578_23; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_503 = _T_4840 ? _T_4289_24 : _T_5578_24; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_504 = _T_4840 ? _T_4289_25 : _T_5578_25; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_505 = _T_4840 ? _T_4289_26 : _T_5578_26; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_506 = _T_4840 ? _T_4289_27 : _T_5578_27; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_507 = _T_4840 ? _T_4289_28 : _T_5578_28; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_508 = _T_4840 ? _T_4289_29 : _T_5578_29; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_509 = _T_4840 ? _T_4289_30 : _T_5578_30; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_510 = _T_4840 ? _T_4289_31 : _T_5578_31; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_511 = _T_4840 ? _T_4289_32 : _T_5578_32; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_512 = _T_4840 ? _T_4289_33 : _T_5578_33; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_513 = _T_4840 ? _T_4289_34 : _T_5578_34; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_514 = _T_4840 ? _T_4289_35 : _T_5578_35; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_515 = _T_4840 ? _T_4289_36 : _T_5578_36; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_516 = _T_4840 ? _T_4289_37 : _T_5578_37; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_517 = _T_4840 ? _T_4289_38 : _T_5578_38; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_518 = _T_4840 ? _T_4289_39 : _T_5578_39; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_519 = _T_4840 ? _T_4289_40 : _T_5578_40; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_520 = _T_4840 ? _T_4289_41 : _T_5578_41; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_521 = _T_4840 ? _T_4289_42 : _T_5578_42; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_522 = _T_4840 ? _T_4289_43 : _T_5578_43; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_523 = _T_4840 ? _T_4289_44 : _T_5578_44; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_524 = _T_4840 ? _T_4289_45 : _T_5578_45; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_525 = _T_4840 ? _T_4289_46 : _T_5578_46; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_526 = _T_4840 ? _T_4289_47 : _T_5578_47; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_527 = _T_4840 ? _T_4289_48 : _T_5578_48; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_528 = _T_4840 ? _T_4289_49 : _T_5578_49; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_529 = _T_4840 ? _T_4289_50 : _T_5578_50; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_530 = _T_4840 ? _T_4289_51 : _T_5578_51; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_531 = _T_4840 ? _T_4289_52 : _T_5578_52; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_532 = _T_4840 ? _T_4289_53 : _T_5578_53; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_533 = _T_4840 ? _T_4289_54 : _T_5578_54; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_534 = _T_4840 ? _T_4289_55 : _T_5578_55; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_535 = _T_4840 ? _T_4289_56 : _T_5578_56; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_536 = _T_4840 ? _T_4289_57 : _T_5578_57; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_537 = _T_4840 ? _T_4289_58 : _T_5578_58; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_538 = _T_4840 ? _T_4289_59 : _T_5578_59; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_539 = _T_4840 ? _T_4289_60 : _T_5578_60; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_540 = _T_4840 ? _T_4289_61 : _T_5578_61; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_541 = _T_4840 ? _T_4289_62 : _T_5578_62; // @[Reg.scala 20:19:@22833.4]
  assign _GEN_542 = _T_4840 ? _T_4289_63 : _T_5578_63; // @[Reg.scala 20:19:@22833.4]
  assign io_sc2cdma_dat_updt_valid = _T_1166; // @[NV_NVDLA_CSC_dl.scala 308:27:@19950.4]
  assign io_sc2cdma_dat_updt_bits_entries = _T_1172; // @[NV_NVDLA_CSC_dl.scala 310:34:@19960.4]
  assign io_sc2cdma_dat_updt_bits_slices = _T_1169; // @[NV_NVDLA_CSC_dl.scala 309:33:@19955.4]
  assign io_sc2buf_dat_rd_addr_valid = _T_1778; // @[NV_NVDLA_CSC_dl.scala 725:29:@20557.4]
  assign io_sc2buf_dat_rd_addr_bits = _T_1785[12:0]; // @[NV_NVDLA_CSC_dl.scala 726:28:@20558.4]
  assign io_sc2mac_dat_a_valid = _T_4835; // @[NV_NVDLA_CSC_dl.scala 1174:23:@22553.4]
  assign io_sc2mac_dat_a_bits_mask_0 = _T_5114_0; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22702.4]
  assign io_sc2mac_dat_a_bits_mask_1 = _T_5114_1; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22703.4]
  assign io_sc2mac_dat_a_bits_mask_2 = _T_5114_2; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22704.4]
  assign io_sc2mac_dat_a_bits_mask_3 = _T_5114_3; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22705.4]
  assign io_sc2mac_dat_a_bits_mask_4 = _T_5114_4; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22706.4]
  assign io_sc2mac_dat_a_bits_mask_5 = _T_5114_5; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22707.4]
  assign io_sc2mac_dat_a_bits_mask_6 = _T_5114_6; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22708.4]
  assign io_sc2mac_dat_a_bits_mask_7 = _T_5114_7; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22709.4]
  assign io_sc2mac_dat_a_bits_mask_8 = _T_5114_8; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22710.4]
  assign io_sc2mac_dat_a_bits_mask_9 = _T_5114_9; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22711.4]
  assign io_sc2mac_dat_a_bits_mask_10 = _T_5114_10; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22712.4]
  assign io_sc2mac_dat_a_bits_mask_11 = _T_5114_11; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22713.4]
  assign io_sc2mac_dat_a_bits_mask_12 = _T_5114_12; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22714.4]
  assign io_sc2mac_dat_a_bits_mask_13 = _T_5114_13; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22715.4]
  assign io_sc2mac_dat_a_bits_mask_14 = _T_5114_14; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22716.4]
  assign io_sc2mac_dat_a_bits_mask_15 = _T_5114_15; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22717.4]
  assign io_sc2mac_dat_a_bits_mask_16 = _T_5114_16; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22718.4]
  assign io_sc2mac_dat_a_bits_mask_17 = _T_5114_17; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22719.4]
  assign io_sc2mac_dat_a_bits_mask_18 = _T_5114_18; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22720.4]
  assign io_sc2mac_dat_a_bits_mask_19 = _T_5114_19; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22721.4]
  assign io_sc2mac_dat_a_bits_mask_20 = _T_5114_20; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22722.4]
  assign io_sc2mac_dat_a_bits_mask_21 = _T_5114_21; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22723.4]
  assign io_sc2mac_dat_a_bits_mask_22 = _T_5114_22; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22724.4]
  assign io_sc2mac_dat_a_bits_mask_23 = _T_5114_23; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22725.4]
  assign io_sc2mac_dat_a_bits_mask_24 = _T_5114_24; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22726.4]
  assign io_sc2mac_dat_a_bits_mask_25 = _T_5114_25; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22727.4]
  assign io_sc2mac_dat_a_bits_mask_26 = _T_5114_26; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22728.4]
  assign io_sc2mac_dat_a_bits_mask_27 = _T_5114_27; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22729.4]
  assign io_sc2mac_dat_a_bits_mask_28 = _T_5114_28; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22730.4]
  assign io_sc2mac_dat_a_bits_mask_29 = _T_5114_29; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22731.4]
  assign io_sc2mac_dat_a_bits_mask_30 = _T_5114_30; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22732.4]
  assign io_sc2mac_dat_a_bits_mask_31 = _T_5114_31; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22733.4]
  assign io_sc2mac_dat_a_bits_mask_32 = _T_5114_32; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22734.4]
  assign io_sc2mac_dat_a_bits_mask_33 = _T_5114_33; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22735.4]
  assign io_sc2mac_dat_a_bits_mask_34 = _T_5114_34; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22736.4]
  assign io_sc2mac_dat_a_bits_mask_35 = _T_5114_35; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22737.4]
  assign io_sc2mac_dat_a_bits_mask_36 = _T_5114_36; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22738.4]
  assign io_sc2mac_dat_a_bits_mask_37 = _T_5114_37; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22739.4]
  assign io_sc2mac_dat_a_bits_mask_38 = _T_5114_38; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22740.4]
  assign io_sc2mac_dat_a_bits_mask_39 = _T_5114_39; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22741.4]
  assign io_sc2mac_dat_a_bits_mask_40 = _T_5114_40; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22742.4]
  assign io_sc2mac_dat_a_bits_mask_41 = _T_5114_41; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22743.4]
  assign io_sc2mac_dat_a_bits_mask_42 = _T_5114_42; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22744.4]
  assign io_sc2mac_dat_a_bits_mask_43 = _T_5114_43; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22745.4]
  assign io_sc2mac_dat_a_bits_mask_44 = _T_5114_44; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22746.4]
  assign io_sc2mac_dat_a_bits_mask_45 = _T_5114_45; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22747.4]
  assign io_sc2mac_dat_a_bits_mask_46 = _T_5114_46; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22748.4]
  assign io_sc2mac_dat_a_bits_mask_47 = _T_5114_47; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22749.4]
  assign io_sc2mac_dat_a_bits_mask_48 = _T_5114_48; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22750.4]
  assign io_sc2mac_dat_a_bits_mask_49 = _T_5114_49; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22751.4]
  assign io_sc2mac_dat_a_bits_mask_50 = _T_5114_50; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22752.4]
  assign io_sc2mac_dat_a_bits_mask_51 = _T_5114_51; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22753.4]
  assign io_sc2mac_dat_a_bits_mask_52 = _T_5114_52; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22754.4]
  assign io_sc2mac_dat_a_bits_mask_53 = _T_5114_53; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22755.4]
  assign io_sc2mac_dat_a_bits_mask_54 = _T_5114_54; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22756.4]
  assign io_sc2mac_dat_a_bits_mask_55 = _T_5114_55; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22757.4]
  assign io_sc2mac_dat_a_bits_mask_56 = _T_5114_56; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22758.4]
  assign io_sc2mac_dat_a_bits_mask_57 = _T_5114_57; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22759.4]
  assign io_sc2mac_dat_a_bits_mask_58 = _T_5114_58; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22760.4]
  assign io_sc2mac_dat_a_bits_mask_59 = _T_5114_59; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22761.4]
  assign io_sc2mac_dat_a_bits_mask_60 = _T_5114_60; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22762.4]
  assign io_sc2mac_dat_a_bits_mask_61 = _T_5114_61; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22763.4]
  assign io_sc2mac_dat_a_bits_mask_62 = _T_5114_62; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22764.4]
  assign io_sc2mac_dat_a_bits_mask_63 = _T_5114_63; // @[NV_NVDLA_CSC_dl.scala 1178:27:@22765.4]
  assign io_sc2mac_dat_a_bits_data_0 = _T_5776; // @[NV_NVDLA_CSC_dl.scala 1181:34:@22967.4]
  assign io_sc2mac_dat_a_bits_data_1 = _T_5780; // @[NV_NVDLA_CSC_dl.scala 1181:34:@22977.4]
  assign io_sc2mac_dat_a_bits_data_2 = _T_5784; // @[NV_NVDLA_CSC_dl.scala 1181:34:@22987.4]
  assign io_sc2mac_dat_a_bits_data_3 = _T_5788; // @[NV_NVDLA_CSC_dl.scala 1181:34:@22997.4]
  assign io_sc2mac_dat_a_bits_data_4 = _T_5792; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23007.4]
  assign io_sc2mac_dat_a_bits_data_5 = _T_5796; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23017.4]
  assign io_sc2mac_dat_a_bits_data_6 = _T_5800; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23027.4]
  assign io_sc2mac_dat_a_bits_data_7 = _T_5804; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23037.4]
  assign io_sc2mac_dat_a_bits_data_8 = _T_5808; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23047.4]
  assign io_sc2mac_dat_a_bits_data_9 = _T_5812; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23057.4]
  assign io_sc2mac_dat_a_bits_data_10 = _T_5816; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23067.4]
  assign io_sc2mac_dat_a_bits_data_11 = _T_5820; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23077.4]
  assign io_sc2mac_dat_a_bits_data_12 = _T_5824; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23087.4]
  assign io_sc2mac_dat_a_bits_data_13 = _T_5828; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23097.4]
  assign io_sc2mac_dat_a_bits_data_14 = _T_5832; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23107.4]
  assign io_sc2mac_dat_a_bits_data_15 = _T_5836; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23117.4]
  assign io_sc2mac_dat_a_bits_data_16 = _T_5840; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23127.4]
  assign io_sc2mac_dat_a_bits_data_17 = _T_5844; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23137.4]
  assign io_sc2mac_dat_a_bits_data_18 = _T_5848; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23147.4]
  assign io_sc2mac_dat_a_bits_data_19 = _T_5852; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23157.4]
  assign io_sc2mac_dat_a_bits_data_20 = _T_5856; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23167.4]
  assign io_sc2mac_dat_a_bits_data_21 = _T_5860; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23177.4]
  assign io_sc2mac_dat_a_bits_data_22 = _T_5864; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23187.4]
  assign io_sc2mac_dat_a_bits_data_23 = _T_5868; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23197.4]
  assign io_sc2mac_dat_a_bits_data_24 = _T_5872; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23207.4]
  assign io_sc2mac_dat_a_bits_data_25 = _T_5876; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23217.4]
  assign io_sc2mac_dat_a_bits_data_26 = _T_5880; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23227.4]
  assign io_sc2mac_dat_a_bits_data_27 = _T_5884; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23237.4]
  assign io_sc2mac_dat_a_bits_data_28 = _T_5888; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23247.4]
  assign io_sc2mac_dat_a_bits_data_29 = _T_5892; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23257.4]
  assign io_sc2mac_dat_a_bits_data_30 = _T_5896; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23267.4]
  assign io_sc2mac_dat_a_bits_data_31 = _T_5900; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23277.4]
  assign io_sc2mac_dat_a_bits_data_32 = _T_5904; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23287.4]
  assign io_sc2mac_dat_a_bits_data_33 = _T_5908; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23297.4]
  assign io_sc2mac_dat_a_bits_data_34 = _T_5912; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23307.4]
  assign io_sc2mac_dat_a_bits_data_35 = _T_5916; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23317.4]
  assign io_sc2mac_dat_a_bits_data_36 = _T_5920; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23327.4]
  assign io_sc2mac_dat_a_bits_data_37 = _T_5924; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23337.4]
  assign io_sc2mac_dat_a_bits_data_38 = _T_5928; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23347.4]
  assign io_sc2mac_dat_a_bits_data_39 = _T_5932; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23357.4]
  assign io_sc2mac_dat_a_bits_data_40 = _T_5936; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23367.4]
  assign io_sc2mac_dat_a_bits_data_41 = _T_5940; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23377.4]
  assign io_sc2mac_dat_a_bits_data_42 = _T_5944; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23387.4]
  assign io_sc2mac_dat_a_bits_data_43 = _T_5948; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23397.4]
  assign io_sc2mac_dat_a_bits_data_44 = _T_5952; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23407.4]
  assign io_sc2mac_dat_a_bits_data_45 = _T_5956; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23417.4]
  assign io_sc2mac_dat_a_bits_data_46 = _T_5960; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23427.4]
  assign io_sc2mac_dat_a_bits_data_47 = _T_5964; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23437.4]
  assign io_sc2mac_dat_a_bits_data_48 = _T_5968; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23447.4]
  assign io_sc2mac_dat_a_bits_data_49 = _T_5972; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23457.4]
  assign io_sc2mac_dat_a_bits_data_50 = _T_5976; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23467.4]
  assign io_sc2mac_dat_a_bits_data_51 = _T_5980; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23477.4]
  assign io_sc2mac_dat_a_bits_data_52 = _T_5984; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23487.4]
  assign io_sc2mac_dat_a_bits_data_53 = _T_5988; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23497.4]
  assign io_sc2mac_dat_a_bits_data_54 = _T_5992; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23507.4]
  assign io_sc2mac_dat_a_bits_data_55 = _T_5996; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23517.4]
  assign io_sc2mac_dat_a_bits_data_56 = _T_6000; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23527.4]
  assign io_sc2mac_dat_a_bits_data_57 = _T_6004; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23537.4]
  assign io_sc2mac_dat_a_bits_data_58 = _T_6008; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23547.4]
  assign io_sc2mac_dat_a_bits_data_59 = _T_6012; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23557.4]
  assign io_sc2mac_dat_a_bits_data_60 = _T_6016; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23567.4]
  assign io_sc2mac_dat_a_bits_data_61 = _T_6020; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23577.4]
  assign io_sc2mac_dat_a_bits_data_62 = _T_6024; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23587.4]
  assign io_sc2mac_dat_a_bits_data_63 = _T_6028; // @[NV_NVDLA_CSC_dl.scala 1181:34:@23597.4]
  assign io_sc2mac_dat_a_bits_pd = _T_4842; // @[NV_NVDLA_CSC_dl.scala 1176:25:@22562.4]
  assign io_sc2mac_dat_b_valid = _T_4838; // @[NV_NVDLA_CSC_dl.scala 1175:23:@22556.4]
  assign io_sc2mac_dat_b_bits_mask_0 = _T_5578_0; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22899.4]
  assign io_sc2mac_dat_b_bits_mask_1 = _T_5578_1; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22900.4]
  assign io_sc2mac_dat_b_bits_mask_2 = _T_5578_2; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22901.4]
  assign io_sc2mac_dat_b_bits_mask_3 = _T_5578_3; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22902.4]
  assign io_sc2mac_dat_b_bits_mask_4 = _T_5578_4; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22903.4]
  assign io_sc2mac_dat_b_bits_mask_5 = _T_5578_5; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22904.4]
  assign io_sc2mac_dat_b_bits_mask_6 = _T_5578_6; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22905.4]
  assign io_sc2mac_dat_b_bits_mask_7 = _T_5578_7; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22906.4]
  assign io_sc2mac_dat_b_bits_mask_8 = _T_5578_8; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22907.4]
  assign io_sc2mac_dat_b_bits_mask_9 = _T_5578_9; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22908.4]
  assign io_sc2mac_dat_b_bits_mask_10 = _T_5578_10; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22909.4]
  assign io_sc2mac_dat_b_bits_mask_11 = _T_5578_11; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22910.4]
  assign io_sc2mac_dat_b_bits_mask_12 = _T_5578_12; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22911.4]
  assign io_sc2mac_dat_b_bits_mask_13 = _T_5578_13; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22912.4]
  assign io_sc2mac_dat_b_bits_mask_14 = _T_5578_14; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22913.4]
  assign io_sc2mac_dat_b_bits_mask_15 = _T_5578_15; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22914.4]
  assign io_sc2mac_dat_b_bits_mask_16 = _T_5578_16; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22915.4]
  assign io_sc2mac_dat_b_bits_mask_17 = _T_5578_17; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22916.4]
  assign io_sc2mac_dat_b_bits_mask_18 = _T_5578_18; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22917.4]
  assign io_sc2mac_dat_b_bits_mask_19 = _T_5578_19; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22918.4]
  assign io_sc2mac_dat_b_bits_mask_20 = _T_5578_20; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22919.4]
  assign io_sc2mac_dat_b_bits_mask_21 = _T_5578_21; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22920.4]
  assign io_sc2mac_dat_b_bits_mask_22 = _T_5578_22; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22921.4]
  assign io_sc2mac_dat_b_bits_mask_23 = _T_5578_23; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22922.4]
  assign io_sc2mac_dat_b_bits_mask_24 = _T_5578_24; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22923.4]
  assign io_sc2mac_dat_b_bits_mask_25 = _T_5578_25; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22924.4]
  assign io_sc2mac_dat_b_bits_mask_26 = _T_5578_26; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22925.4]
  assign io_sc2mac_dat_b_bits_mask_27 = _T_5578_27; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22926.4]
  assign io_sc2mac_dat_b_bits_mask_28 = _T_5578_28; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22927.4]
  assign io_sc2mac_dat_b_bits_mask_29 = _T_5578_29; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22928.4]
  assign io_sc2mac_dat_b_bits_mask_30 = _T_5578_30; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22929.4]
  assign io_sc2mac_dat_b_bits_mask_31 = _T_5578_31; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22930.4]
  assign io_sc2mac_dat_b_bits_mask_32 = _T_5578_32; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22931.4]
  assign io_sc2mac_dat_b_bits_mask_33 = _T_5578_33; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22932.4]
  assign io_sc2mac_dat_b_bits_mask_34 = _T_5578_34; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22933.4]
  assign io_sc2mac_dat_b_bits_mask_35 = _T_5578_35; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22934.4]
  assign io_sc2mac_dat_b_bits_mask_36 = _T_5578_36; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22935.4]
  assign io_sc2mac_dat_b_bits_mask_37 = _T_5578_37; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22936.4]
  assign io_sc2mac_dat_b_bits_mask_38 = _T_5578_38; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22937.4]
  assign io_sc2mac_dat_b_bits_mask_39 = _T_5578_39; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22938.4]
  assign io_sc2mac_dat_b_bits_mask_40 = _T_5578_40; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22939.4]
  assign io_sc2mac_dat_b_bits_mask_41 = _T_5578_41; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22940.4]
  assign io_sc2mac_dat_b_bits_mask_42 = _T_5578_42; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22941.4]
  assign io_sc2mac_dat_b_bits_mask_43 = _T_5578_43; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22942.4]
  assign io_sc2mac_dat_b_bits_mask_44 = _T_5578_44; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22943.4]
  assign io_sc2mac_dat_b_bits_mask_45 = _T_5578_45; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22944.4]
  assign io_sc2mac_dat_b_bits_mask_46 = _T_5578_46; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22945.4]
  assign io_sc2mac_dat_b_bits_mask_47 = _T_5578_47; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22946.4]
  assign io_sc2mac_dat_b_bits_mask_48 = _T_5578_48; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22947.4]
  assign io_sc2mac_dat_b_bits_mask_49 = _T_5578_49; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22948.4]
  assign io_sc2mac_dat_b_bits_mask_50 = _T_5578_50; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22949.4]
  assign io_sc2mac_dat_b_bits_mask_51 = _T_5578_51; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22950.4]
  assign io_sc2mac_dat_b_bits_mask_52 = _T_5578_52; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22951.4]
  assign io_sc2mac_dat_b_bits_mask_53 = _T_5578_53; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22952.4]
  assign io_sc2mac_dat_b_bits_mask_54 = _T_5578_54; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22953.4]
  assign io_sc2mac_dat_b_bits_mask_55 = _T_5578_55; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22954.4]
  assign io_sc2mac_dat_b_bits_mask_56 = _T_5578_56; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22955.4]
  assign io_sc2mac_dat_b_bits_mask_57 = _T_5578_57; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22956.4]
  assign io_sc2mac_dat_b_bits_mask_58 = _T_5578_58; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22957.4]
  assign io_sc2mac_dat_b_bits_mask_59 = _T_5578_59; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22958.4]
  assign io_sc2mac_dat_b_bits_mask_60 = _T_5578_60; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22959.4]
  assign io_sc2mac_dat_b_bits_mask_61 = _T_5578_61; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22960.4]
  assign io_sc2mac_dat_b_bits_mask_62 = _T_5578_62; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22961.4]
  assign io_sc2mac_dat_b_bits_mask_63 = _T_5578_63; // @[NV_NVDLA_CSC_dl.scala 1179:27:@22962.4]
  assign io_sc2mac_dat_b_bits_data_0 = _T_5778; // @[NV_NVDLA_CSC_dl.scala 1182:34:@22972.4]
  assign io_sc2mac_dat_b_bits_data_1 = _T_5782; // @[NV_NVDLA_CSC_dl.scala 1182:34:@22982.4]
  assign io_sc2mac_dat_b_bits_data_2 = _T_5786; // @[NV_NVDLA_CSC_dl.scala 1182:34:@22992.4]
  assign io_sc2mac_dat_b_bits_data_3 = _T_5790; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23002.4]
  assign io_sc2mac_dat_b_bits_data_4 = _T_5794; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23012.4]
  assign io_sc2mac_dat_b_bits_data_5 = _T_5798; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23022.4]
  assign io_sc2mac_dat_b_bits_data_6 = _T_5802; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23032.4]
  assign io_sc2mac_dat_b_bits_data_7 = _T_5806; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23042.4]
  assign io_sc2mac_dat_b_bits_data_8 = _T_5810; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23052.4]
  assign io_sc2mac_dat_b_bits_data_9 = _T_5814; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23062.4]
  assign io_sc2mac_dat_b_bits_data_10 = _T_5818; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23072.4]
  assign io_sc2mac_dat_b_bits_data_11 = _T_5822; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23082.4]
  assign io_sc2mac_dat_b_bits_data_12 = _T_5826; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23092.4]
  assign io_sc2mac_dat_b_bits_data_13 = _T_5830; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23102.4]
  assign io_sc2mac_dat_b_bits_data_14 = _T_5834; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23112.4]
  assign io_sc2mac_dat_b_bits_data_15 = _T_5838; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23122.4]
  assign io_sc2mac_dat_b_bits_data_16 = _T_5842; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23132.4]
  assign io_sc2mac_dat_b_bits_data_17 = _T_5846; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23142.4]
  assign io_sc2mac_dat_b_bits_data_18 = _T_5850; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23152.4]
  assign io_sc2mac_dat_b_bits_data_19 = _T_5854; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23162.4]
  assign io_sc2mac_dat_b_bits_data_20 = _T_5858; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23172.4]
  assign io_sc2mac_dat_b_bits_data_21 = _T_5862; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23182.4]
  assign io_sc2mac_dat_b_bits_data_22 = _T_5866; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23192.4]
  assign io_sc2mac_dat_b_bits_data_23 = _T_5870; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23202.4]
  assign io_sc2mac_dat_b_bits_data_24 = _T_5874; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23212.4]
  assign io_sc2mac_dat_b_bits_data_25 = _T_5878; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23222.4]
  assign io_sc2mac_dat_b_bits_data_26 = _T_5882; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23232.4]
  assign io_sc2mac_dat_b_bits_data_27 = _T_5886; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23242.4]
  assign io_sc2mac_dat_b_bits_data_28 = _T_5890; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23252.4]
  assign io_sc2mac_dat_b_bits_data_29 = _T_5894; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23262.4]
  assign io_sc2mac_dat_b_bits_data_30 = _T_5898; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23272.4]
  assign io_sc2mac_dat_b_bits_data_31 = _T_5902; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23282.4]
  assign io_sc2mac_dat_b_bits_data_32 = _T_5906; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23292.4]
  assign io_sc2mac_dat_b_bits_data_33 = _T_5910; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23302.4]
  assign io_sc2mac_dat_b_bits_data_34 = _T_5914; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23312.4]
  assign io_sc2mac_dat_b_bits_data_35 = _T_5918; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23322.4]
  assign io_sc2mac_dat_b_bits_data_36 = _T_5922; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23332.4]
  assign io_sc2mac_dat_b_bits_data_37 = _T_5926; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23342.4]
  assign io_sc2mac_dat_b_bits_data_38 = _T_5930; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23352.4]
  assign io_sc2mac_dat_b_bits_data_39 = _T_5934; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23362.4]
  assign io_sc2mac_dat_b_bits_data_40 = _T_5938; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23372.4]
  assign io_sc2mac_dat_b_bits_data_41 = _T_5942; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23382.4]
  assign io_sc2mac_dat_b_bits_data_42 = _T_5946; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23392.4]
  assign io_sc2mac_dat_b_bits_data_43 = _T_5950; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23402.4]
  assign io_sc2mac_dat_b_bits_data_44 = _T_5954; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23412.4]
  assign io_sc2mac_dat_b_bits_data_45 = _T_5958; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23422.4]
  assign io_sc2mac_dat_b_bits_data_46 = _T_5962; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23432.4]
  assign io_sc2mac_dat_b_bits_data_47 = _T_5966; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23442.4]
  assign io_sc2mac_dat_b_bits_data_48 = _T_5970; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23452.4]
  assign io_sc2mac_dat_b_bits_data_49 = _T_5974; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23462.4]
  assign io_sc2mac_dat_b_bits_data_50 = _T_5978; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23472.4]
  assign io_sc2mac_dat_b_bits_data_51 = _T_5982; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23482.4]
  assign io_sc2mac_dat_b_bits_data_52 = _T_5986; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23492.4]
  assign io_sc2mac_dat_b_bits_data_53 = _T_5990; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23502.4]
  assign io_sc2mac_dat_b_bits_data_54 = _T_5994; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23512.4]
  assign io_sc2mac_dat_b_bits_data_55 = _T_5998; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23522.4]
  assign io_sc2mac_dat_b_bits_data_56 = _T_6002; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23532.4]
  assign io_sc2mac_dat_b_bits_data_57 = _T_6006; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23542.4]
  assign io_sc2mac_dat_b_bits_data_58 = _T_6010; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23552.4]
  assign io_sc2mac_dat_b_bits_data_59 = _T_6014; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23562.4]
  assign io_sc2mac_dat_b_bits_data_60 = _T_6018; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23572.4]
  assign io_sc2mac_dat_b_bits_data_61 = _T_6022; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23582.4]
  assign io_sc2mac_dat_b_bits_data_62 = _T_6026; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23592.4]
  assign io_sc2mac_dat_b_bits_data_63 = _T_6030; // @[NV_NVDLA_CSC_dl.scala 1182:34:@23602.4]
  assign io_sc2mac_dat_b_bits_pd = _T_4846; // @[NV_NVDLA_CSC_dl.scala 1177:25:@22568.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_715 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_722 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_729 = _RAND_2[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_736 = _RAND_3[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_743 = _RAND_4[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_750 = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_757 = _RAND_6[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_771 = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_778 = _RAND_8[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_785 = _RAND_9[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_792 = _RAND_10[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  _T_831 = _RAND_11[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_838 = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_845 = _RAND_13[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_852 = _RAND_14[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_859 = _RAND_15[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_866 = _RAND_16[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_869 = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_872 = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_878 = _RAND_19[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_881 = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_884 = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_887 = _RAND_22[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_893 = _RAND_23[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_896 = _RAND_24[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_902 = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_905 = _RAND_26[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_908 = _RAND_27[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_915 = _RAND_28[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_922 = _RAND_29[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_932 = _RAND_30[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_939 = _RAND_31[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_946 = _RAND_32[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_953 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_960 = _RAND_34[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_967 = _RAND_35[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_974 = _RAND_36[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_981 = _RAND_37[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_988 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_995 = _RAND_39[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_1002 = _RAND_40[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_1009 = _RAND_41[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_1016 = _RAND_42[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_1023 = _RAND_43[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_1076 = _RAND_44[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_2217 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_2211 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_2208 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_2231 = _RAND_48[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_2225 = _RAND_49[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_2222 = _RAND_50[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_1166 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_1169 = _RAND_52[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_1172 = _RAND_53[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_1177 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_1180 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_1183 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_1186 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_1189 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_1211 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_1214 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_1217 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_1220 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_1225 = _RAND_63[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_1228 = _RAND_64[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_1231 = _RAND_65[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_1234 = _RAND_66[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_1279 = _RAND_67[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_1290 = _RAND_68[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_1306 = _RAND_69[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_1335 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_1329 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_1332 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_1361 = _RAND_73[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_1366 = _RAND_74[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_1369 = _RAND_75[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_1390 = _RAND_76[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_1404 = _RAND_77[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_1407 = _RAND_78[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_1410 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_1413 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_1416 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_1419 = _RAND_82[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_1424 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_1427 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_1539 = _RAND_85[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_1542 = _RAND_86[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_1616 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_1619 = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_1622 = _RAND_89[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_1625 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_1628 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_1631 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_1634 = _RAND_93[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_1637 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_1640 = _RAND_95[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_1643 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_1648 = _RAND_97[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_1651 = _RAND_98[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_1654 = _RAND_99[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_1657 = _RAND_100[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_1660 = _RAND_101[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_1663 = _RAND_102[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_1666 = _RAND_103[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_1759_0 = _RAND_104[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_1759_1 = _RAND_105[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_1759_2 = _RAND_106[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_1759_3 = _RAND_107[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_1778 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_1785 = _RAND_109[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_1788 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_1794 = _RAND_111[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_1797 = _RAND_112[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_1800 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_1803 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_1806 = _RAND_115[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_1809 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_1812 = _RAND_117[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_1815 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_1818 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_1821 = _RAND_120[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_1943 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_1946 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_1949 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_1952 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_1955 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_1958 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_1963 = _RAND_127[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_1966 = _RAND_128[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_1969 = _RAND_129[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_1972 = _RAND_130[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_1975 = _RAND_131[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_1978 = _RAND_132[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_2051 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_2063 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {16{`RANDOM}};
  _T_2074 = _RAND_135[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {16{`RANDOM}};
  _T_2082 = _RAND_136[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_2182 = _RAND_137[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_2185 = _RAND_138[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_2188 = _RAND_139[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_2191 = _RAND_140[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_2194 = _RAND_141[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_2197 = _RAND_142[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_2200 = _RAND_143[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_2203 = _RAND_144[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_2214 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_2228 = _RAND_146[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {8{`RANDOM}};
  _T_2611 = _RAND_147[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {4{`RANDOM}};
  _T_2613 = _RAND_148[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {4{`RANDOM}};
  _T_2615 = _RAND_149[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {4{`RANDOM}};
  _T_2617 = _RAND_150[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {4{`RANDOM}};
  _T_2619 = _RAND_151[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {4{`RANDOM}};
  _T_2621 = _RAND_152[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_3419 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_3689_0 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_3689_1 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_3689_2 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_3689_3 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_3689_4 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_3689_5 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_3689_6 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_3689_7 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_3689_8 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_3689_9 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_3689_10 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_3689_11 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_3689_12 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_3689_13 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_3689_14 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_3689_15 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_3689_16 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_3689_17 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_3689_18 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_3689_19 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_3689_20 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_3689_21 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_3689_22 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_3689_23 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_3689_24 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_3689_25 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_3689_26 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_3689_27 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_3689_28 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_3689_29 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_3689_30 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_3689_31 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_3689_32 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_3689_33 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_3689_34 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_3689_35 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_3689_36 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_3689_37 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_3689_38 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_3689_39 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_3689_40 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_3689_41 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_3689_42 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_3689_43 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_3689_44 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_3689_45 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_3689_46 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_3689_47 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_3689_48 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_3689_49 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_3689_50 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_3689_51 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_3689_52 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_3689_53 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_3689_54 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_3689_55 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_3689_56 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_3689_57 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_3689_58 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_3689_59 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_3689_60 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_3689_61 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_3689_62 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_3689_63 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_3889_0 = _RAND_218[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_3889_1 = _RAND_219[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_3889_2 = _RAND_220[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_3889_3 = _RAND_221[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_3889_4 = _RAND_222[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_3889_5 = _RAND_223[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_3889_6 = _RAND_224[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_3889_7 = _RAND_225[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_3889_8 = _RAND_226[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_3889_9 = _RAND_227[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_3889_10 = _RAND_228[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_3889_11 = _RAND_229[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_3889_12 = _RAND_230[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_3889_13 = _RAND_231[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_3889_14 = _RAND_232[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_3889_15 = _RAND_233[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_3889_16 = _RAND_234[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_3889_17 = _RAND_235[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_3889_18 = _RAND_236[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_3889_19 = _RAND_237[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_3889_20 = _RAND_238[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_3889_21 = _RAND_239[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_3889_22 = _RAND_240[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_3889_23 = _RAND_241[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_3889_24 = _RAND_242[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_3889_25 = _RAND_243[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_3889_26 = _RAND_244[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_3889_27 = _RAND_245[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_3889_28 = _RAND_246[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_3889_29 = _RAND_247[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_3889_30 = _RAND_248[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_3889_31 = _RAND_249[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_3889_32 = _RAND_250[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_3889_33 = _RAND_251[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_3889_34 = _RAND_252[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_3889_35 = _RAND_253[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_3889_36 = _RAND_254[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_3889_37 = _RAND_255[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_3889_38 = _RAND_256[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_3889_39 = _RAND_257[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_3889_40 = _RAND_258[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_3889_41 = _RAND_259[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_3889_42 = _RAND_260[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_3889_43 = _RAND_261[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_3889_44 = _RAND_262[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_3889_45 = _RAND_263[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_3889_46 = _RAND_264[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_3889_47 = _RAND_265[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_3889_48 = _RAND_266[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_3889_49 = _RAND_267[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_3889_50 = _RAND_268[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_3889_51 = _RAND_269[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_3889_52 = _RAND_270[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_3889_53 = _RAND_271[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_3889_54 = _RAND_272[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_3889_55 = _RAND_273[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_3889_56 = _RAND_274[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_3889_57 = _RAND_275[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_3889_58 = _RAND_276[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_3889_59 = _RAND_277[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_3889_60 = _RAND_278[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_3889_61 = _RAND_279[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_3889_62 = _RAND_280[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_3889_63 = _RAND_281[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_4022 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_4289_0 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_4289_1 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_4289_2 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_4289_3 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_4289_4 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_4289_5 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_4289_6 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_4289_7 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_4289_8 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_4289_9 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_4289_10 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_4289_11 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_4289_12 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_4289_13 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_4289_14 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_4289_15 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_4289_16 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_4289_17 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_4289_18 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_4289_19 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_4289_20 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_4289_21 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_4289_22 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_4289_23 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_4289_24 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_4289_25 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_4289_26 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_4289_27 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_4289_28 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_4289_29 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_4289_30 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_4289_31 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_4289_32 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_4289_33 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_4289_34 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_4289_35 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_4289_36 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_4289_37 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_4289_38 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_4289_39 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_4289_40 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_4289_41 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_4289_42 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_4289_43 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_4289_44 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_4289_45 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_4289_46 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_4289_47 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_4289_48 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_4289_49 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_4289_50 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_4289_51 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_4289_52 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_4289_53 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_4289_54 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_4289_55 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_4289_56 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_4289_57 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_4289_58 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_4289_59 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_4289_60 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_4289_61 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_4289_62 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_4289_63 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_4488 = _RAND_347[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_4492_0 = _RAND_348[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_4492_1 = _RAND_349[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_4492_2 = _RAND_350[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_4492_3 = _RAND_351[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_4492_4 = _RAND_352[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_4492_5 = _RAND_353[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_4492_6 = _RAND_354[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_4492_7 = _RAND_355[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_4492_8 = _RAND_356[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_4492_9 = _RAND_357[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_4492_10 = _RAND_358[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_4492_11 = _RAND_359[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_4492_12 = _RAND_360[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_4492_13 = _RAND_361[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_4492_14 = _RAND_362[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_4492_15 = _RAND_363[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_4492_16 = _RAND_364[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_4492_17 = _RAND_365[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_4492_18 = _RAND_366[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_4492_19 = _RAND_367[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_4492_20 = _RAND_368[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_4492_21 = _RAND_369[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_4492_22 = _RAND_370[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_4492_23 = _RAND_371[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_4492_24 = _RAND_372[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_4492_25 = _RAND_373[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_4492_26 = _RAND_374[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_4492_27 = _RAND_375[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_4492_28 = _RAND_376[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_4492_29 = _RAND_377[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_4492_30 = _RAND_378[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_4492_31 = _RAND_379[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_4492_32 = _RAND_380[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_4492_33 = _RAND_381[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_4492_34 = _RAND_382[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_4492_35 = _RAND_383[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_4492_36 = _RAND_384[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_4492_37 = _RAND_385[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_4492_38 = _RAND_386[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_4492_39 = _RAND_387[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_4492_40 = _RAND_388[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_4492_41 = _RAND_389[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_4492_42 = _RAND_390[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_4492_43 = _RAND_391[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_4492_44 = _RAND_392[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_4492_45 = _RAND_393[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_4492_46 = _RAND_394[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_4492_47 = _RAND_395[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_4492_48 = _RAND_396[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_4492_49 = _RAND_397[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_4492_50 = _RAND_398[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_4492_51 = _RAND_399[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_4492_52 = _RAND_400[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_4492_53 = _RAND_401[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_4492_54 = _RAND_402[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_4492_55 = _RAND_403[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_4492_56 = _RAND_404[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_4492_57 = _RAND_405[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_4492_58 = _RAND_406[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_4492_59 = _RAND_407[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_4492_60 = _RAND_408[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_4492_61 = _RAND_409[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_4492_62 = _RAND_410[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_4492_63 = _RAND_411[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_4829 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_4835 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_4838 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_4842 = _RAND_415[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_4846 = _RAND_416[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_5114_0 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_5114_1 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_5114_2 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_5114_3 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_5114_4 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_5114_5 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_5114_6 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_5114_7 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_5114_8 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_5114_9 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_5114_10 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_5114_11 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_5114_12 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_5114_13 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_5114_14 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_5114_15 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_5114_16 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_5114_17 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_5114_18 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_5114_19 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_5114_20 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_5114_21 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_5114_22 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_5114_23 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_5114_24 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_5114_25 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_5114_26 = _RAND_443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_5114_27 = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_5114_28 = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_5114_29 = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_5114_30 = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_5114_31 = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_5114_32 = _RAND_449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_5114_33 = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_5114_34 = _RAND_451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_5114_35 = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_5114_36 = _RAND_453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_5114_37 = _RAND_454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_5114_38 = _RAND_455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_5114_39 = _RAND_456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_5114_40 = _RAND_457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_5114_41 = _RAND_458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_5114_42 = _RAND_459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_5114_43 = _RAND_460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_5114_44 = _RAND_461[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_5114_45 = _RAND_462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_5114_46 = _RAND_463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_5114_47 = _RAND_464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_5114_48 = _RAND_465[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_5114_49 = _RAND_466[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_5114_50 = _RAND_467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_5114_51 = _RAND_468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_5114_52 = _RAND_469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_5114_53 = _RAND_470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_5114_54 = _RAND_471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_5114_55 = _RAND_472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_5114_56 = _RAND_473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_5114_57 = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_5114_58 = _RAND_475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_5114_59 = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_5114_60 = _RAND_477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_5114_61 = _RAND_478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_5114_62 = _RAND_479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_5114_63 = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_5578_0 = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_5578_1 = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_5578_2 = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_5578_3 = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_5578_4 = _RAND_485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_5578_5 = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_5578_6 = _RAND_487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_5578_7 = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_5578_8 = _RAND_489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_5578_9 = _RAND_490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_5578_10 = _RAND_491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_5578_11 = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_5578_12 = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_5578_13 = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_5578_14 = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_5578_15 = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_5578_16 = _RAND_497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_5578_17 = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_5578_18 = _RAND_499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_5578_19 = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_5578_20 = _RAND_501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_5578_21 = _RAND_502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_5578_22 = _RAND_503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_5578_23 = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_5578_24 = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_5578_25 = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_5578_26 = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_5578_27 = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_5578_28 = _RAND_509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_5578_29 = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_5578_30 = _RAND_511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_5578_31 = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_5578_32 = _RAND_513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_5578_33 = _RAND_514[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_5578_34 = _RAND_515[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_5578_35 = _RAND_516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_5578_36 = _RAND_517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_5578_37 = _RAND_518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  _T_5578_38 = _RAND_519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  _T_5578_39 = _RAND_520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  _T_5578_40 = _RAND_521[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  _T_5578_41 = _RAND_522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  _T_5578_42 = _RAND_523[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  _T_5578_43 = _RAND_524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  _T_5578_44 = _RAND_525[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  _T_5578_45 = _RAND_526[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  _T_5578_46 = _RAND_527[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  _T_5578_47 = _RAND_528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  _T_5578_48 = _RAND_529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  _T_5578_49 = _RAND_530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  _T_5578_50 = _RAND_531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  _T_5578_51 = _RAND_532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  _T_5578_52 = _RAND_533[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  _T_5578_53 = _RAND_534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  _T_5578_54 = _RAND_535[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  _T_5578_55 = _RAND_536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  _T_5578_56 = _RAND_537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  _T_5578_57 = _RAND_538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  _T_5578_58 = _RAND_539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  _T_5578_59 = _RAND_540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  _T_5578_60 = _RAND_541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  _T_5578_61 = _RAND_542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  _T_5578_62 = _RAND_543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  _T_5578_63 = _RAND_544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  _T_5776 = _RAND_545[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  _T_5778 = _RAND_546[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  _T_5780 = _RAND_547[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  _T_5782 = _RAND_548[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  _T_5784 = _RAND_549[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  _T_5786 = _RAND_550[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  _T_5788 = _RAND_551[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  _T_5790 = _RAND_552[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  _T_5792 = _RAND_553[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  _T_5794 = _RAND_554[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  _T_5796 = _RAND_555[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  _T_5798 = _RAND_556[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  _T_5800 = _RAND_557[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  _T_5802 = _RAND_558[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  _T_5804 = _RAND_559[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  _T_5806 = _RAND_560[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  _T_5808 = _RAND_561[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  _T_5810 = _RAND_562[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  _T_5812 = _RAND_563[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  _T_5814 = _RAND_564[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  _T_5816 = _RAND_565[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  _T_5818 = _RAND_566[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  _T_5820 = _RAND_567[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  _T_5822 = _RAND_568[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  _T_5824 = _RAND_569[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  _T_5826 = _RAND_570[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  _T_5828 = _RAND_571[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  _T_5830 = _RAND_572[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  _T_5832 = _RAND_573[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  _T_5834 = _RAND_574[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  _T_5836 = _RAND_575[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  _T_5838 = _RAND_576[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  _T_5840 = _RAND_577[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  _T_5842 = _RAND_578[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  _T_5844 = _RAND_579[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  _T_5846 = _RAND_580[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  _T_5848 = _RAND_581[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  _T_5850 = _RAND_582[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  _T_5852 = _RAND_583[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  _T_5854 = _RAND_584[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  _T_5856 = _RAND_585[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  _T_5858 = _RAND_586[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  _T_5860 = _RAND_587[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  _T_5862 = _RAND_588[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  _T_5864 = _RAND_589[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  _T_5866 = _RAND_590[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  _T_5868 = _RAND_591[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  _T_5870 = _RAND_592[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  _T_5872 = _RAND_593[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  _T_5874 = _RAND_594[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  _T_5876 = _RAND_595[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  _T_5878 = _RAND_596[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  _T_5880 = _RAND_597[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  _T_5882 = _RAND_598[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  _T_5884 = _RAND_599[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  _T_5886 = _RAND_600[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  _T_5888 = _RAND_601[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  _T_5890 = _RAND_602[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  _T_5892 = _RAND_603[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  _T_5894 = _RAND_604[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  _T_5896 = _RAND_605[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  _T_5898 = _RAND_606[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  _T_5900 = _RAND_607[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  _T_5902 = _RAND_608[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  _T_5904 = _RAND_609[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  _T_5906 = _RAND_610[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  _T_5908 = _RAND_611[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  _T_5910 = _RAND_612[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  _T_5912 = _RAND_613[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  _T_5914 = _RAND_614[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  _T_5916 = _RAND_615[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  _T_5918 = _RAND_616[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  _T_5920 = _RAND_617[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  _T_5922 = _RAND_618[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  _T_5924 = _RAND_619[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  _T_5926 = _RAND_620[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  _T_5928 = _RAND_621[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  _T_5930 = _RAND_622[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  _T_5932 = _RAND_623[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  _T_5934 = _RAND_624[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  _T_5936 = _RAND_625[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  _T_5938 = _RAND_626[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  _T_5940 = _RAND_627[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  _T_5942 = _RAND_628[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  _T_5944 = _RAND_629[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  _T_5946 = _RAND_630[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  _T_5948 = _RAND_631[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  _T_5950 = _RAND_632[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  _T_5952 = _RAND_633[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  _T_5954 = _RAND_634[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  _T_5956 = _RAND_635[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  _T_5958 = _RAND_636[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  _T_5960 = _RAND_637[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  _T_5962 = _RAND_638[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  _T_5964 = _RAND_639[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  _T_5966 = _RAND_640[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  _T_5968 = _RAND_641[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  _T_5970 = _RAND_642[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  _T_5972 = _RAND_643[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  _T_5974 = _RAND_644[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  _T_5976 = _RAND_645[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  _T_5978 = _RAND_646[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  _T_5980 = _RAND_647[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  _T_5982 = _RAND_648[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  _T_5984 = _RAND_649[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  _T_5986 = _RAND_650[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  _T_5988 = _RAND_651[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  _T_5990 = _RAND_652[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  _T_5992 = _RAND_653[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  _T_5994 = _RAND_654[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  _T_5996 = _RAND_655[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  _T_5998 = _RAND_656[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  _T_6000 = _RAND_657[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  _T_6002 = _RAND_658[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  _T_6004 = _RAND_659[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  _T_6006 = _RAND_660[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  _T_6008 = _RAND_661[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  _T_6010 = _RAND_662[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  _T_6012 = _RAND_663[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  _T_6014 = _RAND_664[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  _T_6016 = _RAND_665[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  _T_6018 = _RAND_666[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  _T_6020 = _RAND_667[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  _T_6022 = _RAND_668[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  _T_6024 = _RAND_669[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  _T_6026 = _RAND_670[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  _T_6028 = _RAND_671[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  _T_6030 = _RAND_672[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_715 <= 1'h0;
    end else begin
      _T_715 <= _T_630;
    end
    if (reset) begin
      _T_722 <= 6'h0;
    end else begin
      if (_T_630) begin
        _T_722 <= 6'h1;
      end
    end
    if (reset) begin
      _T_729 <= 14'h0;
    end else begin
      if (_T_630) begin
        _T_729 <= {{2'd0}, _T_805};
      end
    end
    if (reset) begin
      _T_736 <= 14'h0;
    end else begin
      if (_T_630) begin
        _T_736 <= {{2'd0}, _T_798};
      end
    end
    if (reset) begin
      _T_743 <= 15'h0;
    end else begin
      if (_T_630) begin
        _T_743 <= _T_794;
      end
    end
    if (reset) begin
      _T_750 <= 15'h0;
    end else begin
      if (_T_630) begin
        _T_750 <= _T_797;
      end
    end
    if (reset) begin
      _T_757 <= 13'h0;
    end else begin
      if (_T_630) begin
        _T_757 <= io_reg2dp_dataout_width;
      end
    end
    if (reset) begin
      _T_771 <= 15'h0;
    end else begin
      if (_T_715) begin
        _T_771 <= _T_813;
      end
    end
    if (reset) begin
      _T_778 <= 12'h0;
    end else begin
      if (_T_715) begin
        _T_778 <= _T_800;
      end
    end
    if (reset) begin
      _T_785 <= 12'h0;
    end else begin
      if (_T_715) begin
        _T_785 <= _T_802;
      end
    end
    if (reset) begin
      _T_792 <= 14'h0;
    end else begin
      if (_T_630) begin
        if (io_reg2dp_skip_data_rls) begin
          _T_792 <= _T_807;
        end else begin
          _T_792 <= _T_809;
        end
      end
    end
    if (reset) begin
      _T_831 <= 34'h0;
    end else begin
      if (_T_630) begin
        if (_T_635) begin
          _T_831 <= 34'h3ffffffff;
        end else begin
          _T_831 <= 34'h0;
        end
      end
    end
    if (reset) begin
      _T_838 <= 5'h0;
    end else begin
      if (_T_630) begin
        _T_838 <= _T_1041;
      end
    end
    if (reset) begin
      _T_845 <= 14'h0;
    end else begin
      if (_T_630) begin
        _T_845 <= _T_1043;
      end
    end
    if (reset) begin
      _T_852 <= 13'h0;
    end else begin
      if (_T_630) begin
        _T_852 <= io_reg2dp_datain_width_ext;
      end
    end
    if (reset) begin
      _T_859 <= 13'h0;
    end else begin
      if (_T_630) begin
        _T_859 <= io_reg2dp_datain_height_ext;
      end
    end
    if (reset) begin
      _T_866 <= 11'h0;
    end else begin
      if (_T_630) begin
        _T_866 <= _T_1050;
      end
    end
    if (reset) begin
      _T_869 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_869 <= _T_643;
      end
    end
    if (reset) begin
      _T_872 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_872 <= _T_643;
      end
    end
    if (reset) begin
      _T_878 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_878 <= _T_643;
      end
    end
    if (reset) begin
      _T_881 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_881 <= _T_643;
      end
    end
    if (reset) begin
      _T_884 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_884 <= _T_643;
      end
    end
    if (reset) begin
      _T_887 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_887 <= _T_643;
      end
    end
    if (reset) begin
      _T_893 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_893 <= _T_643;
      end
    end
    if (reset) begin
      _T_896 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_896 <= _T_643;
      end
    end
    if (reset) begin
      _T_902 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_902 <= _T_643;
      end
    end
    if (reset) begin
      _T_905 <= 3'h1;
    end else begin
      if (_T_630) begin
        if (_T_635) begin
          _T_905 <= _T_643;
        end else begin
          _T_905 <= 3'h1;
        end
      end
    end
    if (reset) begin
      _T_908 <= 3'h1;
    end else begin
      if (_T_630) begin
        if (_T_635) begin
          _T_908 <= _T_643;
        end else begin
          _T_908 <= 3'h1;
        end
      end
    end
    if (reset) begin
      _T_915 <= 4'h0;
    end else begin
      if (_T_630) begin
        _T_915 <= _T_650;
      end
    end
    if (reset) begin
      _T_922 <= 4'h0;
    end else begin
      if (_T_630) begin
        _T_922 <= _T_704;
      end
    end
    if (reset) begin
      _T_932 <= 5'h0;
    end else begin
      if (_T_630) begin
        _T_932 <= 5'h0;
      end
    end
    if (reset) begin
      _T_939 <= 7'h0;
    end else begin
      if (_T_630) begin
        if (_T_686) begin
          _T_939 <= _T_679;
        end else begin
          _T_939 <= {{1'd0}, _T_685};
        end
      end
    end
    if (reset) begin
      _T_946 <= 7'h0;
    end else begin
      if (_T_630) begin
        _T_946 <= _T_690;
      end
    end
    if (reset) begin
      _T_953 <= 8'h0;
    end else begin
      if (_T_630) begin
        if (_T_686) begin
          _T_953 <= _T_693;
        end else begin
          _T_953 <= {{1'd0}, _T_698};
        end
      end
    end
    if (reset) begin
      _T_960 <= 7'h0;
    end else begin
      if (_T_630) begin
        _T_960 <= {{1'd0}, _T_662};
      end
    end
    if (reset) begin
      _T_967 <= 12'h0;
    end else begin
      if (_T_630) begin
        _T_967 <= _T_702;
      end
    end
    if (reset) begin
      _T_974 <= 6'h0;
    end else begin
      if (_T_630) begin
        if (_T_635) begin
          _T_974 <= 6'h1;
        end else begin
          _T_974 <= _T_707;
        end
      end
    end
    if (reset) begin
      _T_981 <= 6'h0;
    end else begin
      if (_T_630) begin
        if (_T_635) begin
          _T_981 <= 6'h1;
        end else begin
          _T_981 <= _T_711;
        end
      end
    end
    if (reset) begin
      _T_988 <= 16'h0;
    end else begin
      if (_T_630) begin
        _T_988 <= io_reg2dp_pad_value;
      end
    end
    if (reset) begin
      _T_995 <= 15'h0;
    end else begin
      if (_T_630) begin
        _T_995 <= _T_1054;
      end
    end
    if (reset) begin
      _T_1002 <= 15'h0;
    end else begin
      if (_T_715) begin
        _T_1002 <= _T_743;
      end
    end
    if (reset) begin
      _T_1009 <= 15'h0;
    end else begin
      if (_T_715) begin
        _T_1009 <= _T_743;
      end
    end
    if (reset) begin
      _T_1016 <= 14'h0;
    end else begin
      if (_T_626) begin
        _T_1016 <= _T_792;
      end
    end
    if (reset) begin
      _T_1023 <= 15'h0;
    end else begin
      if (_T_626) begin
        _T_1023 <= _T_813;
      end
    end
    if (reset) begin
      _T_2217 <= 1'h0;
    end else begin
      _T_2217 <= _T_2214;
    end
    if (reset) begin
      _T_2211 <= 1'h0;
    end else begin
      _T_2211 <= _T_2208;
    end
    if (reset) begin
      _T_2208 <= 1'h0;
    end else begin
      _T_2208 <= _T_1958;
    end
    if (reset) begin
      _T_2231 <= 27'h0;
    end else begin
      if (_T_2214) begin
        _T_2231 <= _T_2228;
      end
    end
    if (reset) begin
      _T_2225 <= 27'h0;
    end else begin
      if (_T_2208) begin
        _T_2225 <= _T_2222;
      end
    end
    if (reset) begin
      _T_2222 <= 27'h0;
    end else begin
      if (_T_1958) begin
        _T_2222 <= _T_2240;
      end
    end
    if (reset) begin
      _T_1166 <= 1'h0;
    end else begin
      _T_1166 <= _T_1161;
    end
    if (reset) begin
      _T_1169 <= 14'h0;
    end else begin
      if (_T_1161) begin
        if (_T_1154) begin
          _T_1169 <= _T_729;
        end else begin
          _T_1169 <= _T_1016;
        end
      end
    end
    if (reset) begin
      _T_1172 <= 15'h0;
    end else begin
      if (_T_1161) begin
        if (_T_1154) begin
          _T_1172 <= _T_771;
        end else begin
          _T_1172 <= _T_1023;
        end
      end
    end
    if (reset) begin
      _T_1177 <= 1'h0;
    end else begin
      _T_1177 <= io_sg2dl_pd_valid;
    end
    if (reset) begin
      _T_1180 <= 1'h0;
    end else begin
      _T_1180 <= _T_1177;
    end
    if (reset) begin
      _T_1183 <= 1'h0;
    end else begin
      _T_1183 <= _T_1180;
    end
    if (reset) begin
      _T_1186 <= 1'h0;
    end else begin
      _T_1186 <= _T_1183;
    end
    if (reset) begin
      _T_1189 <= 1'h0;
    end else begin
      _T_1189 <= _T_1186;
    end
    if (reset) begin
      _T_1211 <= 1'h0;
    end else begin
      _T_1211 <= _T_1189;
    end
    if (reset) begin
      _T_1214 <= 1'h0;
    end else begin
      _T_1214 <= _T_1211;
    end
    if (reset) begin
      _T_1217 <= 1'h0;
    end else begin
      _T_1217 <= _T_1214;
    end
    if (reset) begin
      _T_1220 <= 1'h0;
    end else begin
      _T_1220 <= _T_1217;
    end
    if (reset) begin
      _T_1225 <= 31'h0;
    end else begin
      if (_T_1189) begin
        _T_1225 <= _T_1222;
      end
    end
    if (reset) begin
      _T_1228 <= 31'h0;
    end else begin
      if (_T_1211) begin
        _T_1228 <= _T_1225;
      end
    end
    if (reset) begin
      _T_1231 <= 31'h0;
    end else begin
      if (_T_1214) begin
        _T_1231 <= _T_1228;
      end
    end
    if (reset) begin
      _T_1234 <= 31'h0;
    end else begin
      if (_T_1217) begin
        _T_1234 <= _T_1231;
      end
    end
    if (reset) begin
      _T_1279 <= 5'h0;
    end else begin
      if (_T_630) begin
        _T_1279 <= 5'h0;
      end else begin
        if (_T_1287) begin
          _T_1279 <= 5'h0;
        end else begin
          _T_1279 <= _T_1284;
        end
      end
    end
    if (reset) begin
      _T_1290 <= 2'h0;
    end else begin
      if (_T_1300) begin
        if (_T_1301) begin
          _T_1290 <= 2'h0;
        end else begin
          _T_1290 <= _T_1295;
        end
      end
    end
    if (reset) begin
      _T_1306 <= 7'h0;
    end else begin
      if (_T_1318) begin
        if (_T_630) begin
          _T_1306 <= 7'h0;
        end else begin
          if (_T_1321) begin
            _T_1306 <= 7'h0;
          end else begin
            if (_T_1316) begin
              _T_1306 <= 7'h0;
            end else begin
              _T_1306 <= _T_1313;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1335 <= 1'h0;
    end else begin
      if (_T_1242) begin
        _T_1335 <= 1'h1;
      end else begin
        if (_T_1355) begin
          _T_1335 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_1329 <= 1'h0;
    end else begin
      if (_T_1338) begin
        _T_1329 <= 1'h0;
      end else begin
        if (_T_1242) begin
          _T_1329 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_1332 <= 1'h0;
    end else begin
      _T_1332 <= _T_1343;
    end
    if (reset) begin
      _T_1361 <= 8'h0;
    end else begin
      if (_T_1358) begin
        _T_1361 <= _T_1363;
      end
    end
    if (reset) begin
      _T_1366 <= 13'h0;
    end else begin
      if (_T_1384) begin
        if (_T_630) begin
          _T_1366 <= {{9'd0}, _T_648};
        end else begin
          if (_T_1378) begin
            _T_1366 <= _T_1369;
          end else begin
            if (_T_1374) begin
              _T_1366 <= {{9'd0}, _T_648};
            end else begin
              _T_1366 <= _T_1371;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1369 <= 13'h0;
    end else begin
      if (_T_1387) begin
        if (_T_630) begin
          _T_1369 <= {{9'd0}, _T_648};
        end else begin
          if (!(_T_1378)) begin
            if (_T_1374) begin
              _T_1369 <= {{9'd0}, _T_648};
            end else begin
              _T_1369 <= _T_1371;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1390 <= 11'h0;
    end else begin
      if (_T_1394) begin
        if (_T_630) begin
          _T_1390 <= 11'h0;
        end else begin
          if (_T_1269) begin
            _T_1390 <= 11'h0;
          end else begin
            _T_1390 <= _T_1399;
          end
        end
      end
    end
    if (reset) begin
      _T_1404 <= 14'h0;
    end else begin
      if (_T_1448) begin
        if (_T_630) begin
          if (_T_635) begin
            _T_1404 <= 14'h0;
          end else begin
            _T_1404 <= _T_1431;
          end
        end else begin
          if (_T_1378) begin
            _T_1404 <= _T_1407;
          end else begin
            if (_T_1374) begin
              if (_T_635) begin
                _T_1404 <= 14'h0;
              end else begin
                _T_1404 <= _T_1431;
              end
            end else begin
              _T_1404 <= _T_1434;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1407 <= 14'h0;
    end else begin
      if (_T_1454) begin
        if (_T_630) begin
          if (_T_635) begin
            _T_1407 <= 14'h0;
          end else begin
            _T_1407 <= _T_1431;
          end
        end else begin
          if (!(_T_1378)) begin
            if (_T_1374) begin
              if (_T_635) begin
                _T_1407 <= 14'h0;
              end else begin
                _T_1407 <= _T_1431;
              end
            end else begin
              _T_1407 <= _T_1434;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1410 <= 16'h0;
    end else begin
      if (_T_1448) begin
        if (_T_715) begin
          _T_1410 <= {{9'd0}, _T_939};
        end else begin
          if (_T_1477) begin
            _T_1410 <= {{9'd0}, _T_939};
          end else begin
            if (_T_1481) begin
              _T_1410 <= _T_1483;
            end else begin
              if (_T_1485) begin
                _T_1410 <= _T_1487;
              end else begin
                if (_T_1490) begin
                  _T_1410 <= _T_1493;
                end else begin
                  if (_T_1495) begin
                    _T_1410 <= _T_1413;
                  end else begin
                    _T_1410 <= _T_1497;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1413 <= 16'h0;
    end else begin
      if (_T_1454) begin
        if (_T_715) begin
          _T_1413 <= {{9'd0}, _T_939};
        end else begin
          if (_T_1477) begin
            _T_1413 <= {{9'd0}, _T_939};
          end else begin
            if (_T_1481) begin
              _T_1413 <= _T_1483;
            end else begin
              if (_T_1485) begin
                _T_1413 <= _T_1487;
              end else begin
                if (_T_1490) begin
                  _T_1413 <= _T_1493;
                end else begin
                  if (!(_T_1495)) begin
                    _T_1413 <= _T_1497;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1416 <= 16'h0;
    end else begin
      if (_T_1526) begin
        if (_T_715) begin
          _T_1416 <= {{9'd0}, _T_939};
        end else begin
          if (_T_1477) begin
            _T_1416 <= {{9'd0}, _T_939};
          end else begin
            if (_T_1481) begin
              _T_1416 <= _T_1483;
            end else begin
              if (_T_1485) begin
                _T_1416 <= _T_1487;
              end else begin
                if (_T_1490) begin
                  _T_1416 <= _T_1493;
                end else begin
                  if (_T_1495) begin
                    _T_1416 <= _T_1413;
                  end else begin
                    _T_1416 <= _T_1497;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1419 <= 13'h2;
    end else begin
      if (_T_1466) begin
        _T_1419 <= 13'h2;
      end else begin
        if (_T_1468) begin
          _T_1419 <= _T_1471;
        end
      end
    end
    if (reset) begin
      _T_1424 <= 1'h0;
    end else begin
      if (_T_1358) begin
        _T_1424 <= _T_1536;
      end
    end
    if (reset) begin
      _T_1427 <= 1'h0;
    end else begin
      if (_T_1358) begin
        if (_T_1528) begin
          _T_1427 <= 1'h1;
        end else begin
          if (_T_1424) begin
            _T_1427 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_1539 <= 14'h0;
    end else begin
      if (_T_1560) begin
        if (_T_1550) begin
          _T_1539 <= _T_1546;
        end else begin
          if (_T_1378) begin
            _T_1539 <= _T_1542;
          end else begin
            if (_T_1374) begin
              _T_1539 <= _T_1548;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1542 <= 14'h0;
    end else begin
      if (_T_1387) begin
        if (_T_1550) begin
          _T_1542 <= _T_1546;
        end else begin
          if (!(_T_1378)) begin
            if (_T_1374) begin
              _T_1542 <= _T_1548;
            end else begin
              _T_1542 <= _T_1539;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1616 <= 1'h0;
    end else begin
      _T_1616 <= _T_1600;
    end
    if (reset) begin
      _T_1619 <= 2'h0;
    end else begin
      if (_T_1358) begin
        _T_1619 <= _T_1605;
      end
    end
    if (reset) begin
      _T_1622 <= 2'h0;
    end else begin
      if (_T_1358) begin
        _T_1622 <= _T_1290;
      end
    end
    if (reset) begin
      _T_1625 <= 1'h0;
    end else begin
      if (_T_1358) begin
        if (_T_1602) begin
          _T_1625 <= _T_1603;
        end else begin
          _T_1625 <= _T_1268;
        end
      end
    end
    if (reset) begin
      _T_1628 <= 1'h0;
    end else begin
      if (_T_1358) begin
        _T_1628 <= _T_1391;
      end
    end
    if (reset) begin
      _T_1631 <= 1'h0;
    end else begin
      if (_T_1358) begin
        if (_T_1242) begin
          _T_1631 <= 1'h1;
        end else begin
          if (_T_1355) begin
            _T_1631 <= 1'h0;
          end else begin
            _T_1631 <= _T_1335;
          end
        end
      end
    end
    if (reset) begin
      _T_1634 <= 2'h0;
    end else begin
      if (_T_1358) begin
        _T_1634 <= _T_1267;
      end
    end
    if (reset) begin
      _T_1637 <= 1'h0;
    end else begin
      if (_T_1608) begin
        _T_1637 <= _T_1242;
      end
    end
    if (reset) begin
      _T_1640 <= 9'h0;
    end else begin
      if (_T_1358) begin
        _T_1640 <= _T_1613;
      end
    end
    if (reset) begin
      _T_1643 <= 1'h0;
    end else begin
      if (_T_1358) begin
        _T_1643 <= _T_1645;
      end
    end
    if (reset) begin
      _T_1648 <= 13'h0;
    end else begin
      if (_T_1394) begin
        if (_T_630) begin
          _T_1648 <= 13'h0;
        end else begin
          if (_T_1673) begin
            _T_1648 <= 13'h0;
          end else begin
            _T_1648 <= _T_1676;
          end
        end
      end
    end
    if (reset) begin
      _T_1651 <= 13'h0;
    end else begin
      if (_T_1682) begin
        _T_1651 <= _T_1648;
      end
    end
    if (reset) begin
      _T_1654 <= 13'h0;
    end else begin
      if (_T_1715) begin
        _T_1654 <= _T_1684;
      end
    end
    if (reset) begin
      _T_1657 <= 13'h0;
    end else begin
      if (_T_1715) begin
        _T_1657 <= _T_1686;
      end
    end
    if (reset) begin
      _T_1660 <= 13'h0;
    end else begin
      if (_T_1715) begin
        _T_1660 <= _T_1688;
      end
    end
    if (reset) begin
      _T_1663 <= 13'h0;
    end else begin
      if (_T_1716) begin
        _T_1663 <= _T_1692;
      end
    end
    if (reset) begin
      _T_1666 <= 13'h0;
    end else begin
      _T_1666 <= _GEN_95[12:0];
    end
    if (reset) begin
      _T_1759_0 <= 13'h1fff;
    end else begin
      _T_1759_0 <= _GEN_96[12:0];
    end
    if (reset) begin
      _T_1759_1 <= 13'h1fff;
    end else begin
      _T_1759_1 <= _GEN_97[12:0];
    end
    if (reset) begin
      _T_1759_2 <= 13'h1fff;
    end else begin
      _T_1759_2 <= _GEN_98[12:0];
    end
    if (reset) begin
      _T_1759_3 <= 13'h1fff;
    end else begin
      _T_1759_3 <= _GEN_99[12:0];
    end
    if (reset) begin
      _T_1778 <= 1'h0;
    end else begin
      _T_1778 <= _T_1891;
    end
    if (reset) begin
      _T_1785 <= 15'h1fff;
    end else begin
      if (_T_1922) begin
        if (_T_1850) begin
          _T_1785 <= 15'h1fff;
        end else begin
          if (_T_1840) begin
            _T_1785 <= _T_1849;
          end else begin
            _T_1785 <= _T_1833;
          end
        end
      end
    end
    if (reset) begin
      _T_1788 <= 1'h0;
    end else begin
      _T_1788 <= _T_1332;
    end
    if (reset) begin
      _T_1794 <= 2'h0;
    end else begin
      if (_T_1335) begin
        _T_1794 <= _T_1619;
      end
    end
    if (reset) begin
      _T_1797 <= 2'h0;
    end else begin
      if (_T_1335) begin
        _T_1797 <= _T_1622;
      end
    end
    if (reset) begin
      _T_1800 <= 1'h0;
    end else begin
      if (_T_1335) begin
        _T_1800 <= _T_1625;
      end
    end
    if (reset) begin
      _T_1803 <= 1'h0;
    end else begin
      if (_T_1335) begin
        _T_1803 <= _T_1628;
      end
    end
    if (reset) begin
      _T_1806 <= 8'h0;
    end else begin
      if (_T_1335) begin
        _T_1806 <= _T_1361;
      end
    end
    if (reset) begin
      _T_1809 <= 1'h0;
    end else begin
      if (_T_1335) begin
        _T_1809 <= _T_1631;
      end
    end
    if (reset) begin
      _T_1812 <= 2'h0;
    end else begin
      if (_T_1335) begin
        _T_1812 <= _T_1634;
      end
    end
    if (reset) begin
      _T_1815 <= 1'h0;
    end else begin
      if (_T_1335) begin
        _T_1815 <= _T_1637;
      end
    end
    if (reset) begin
      _T_1818 <= 1'h0;
    end else begin
      if (_T_1335) begin
        _T_1818 <= _T_1643;
      end
    end
    if (reset) begin
      _T_1821 <= 9'h0;
    end else begin
      if (_T_1335) begin
        _T_1821 <= _T_1640;
      end else begin
        _T_1821 <= {{8'd0}, _T_1335};
      end
    end
    if (reset) begin
      _T_1943 <= 1'h0;
    end else begin
      _T_1943 <= _T_1788;
    end
    if (reset) begin
      _T_1946 <= 1'h0;
    end else begin
      _T_1946 <= _T_1943;
    end
    if (reset) begin
      _T_1949 <= 1'h0;
    end else begin
      _T_1949 <= _T_1946;
    end
    if (reset) begin
      _T_1952 <= 1'h0;
    end else begin
      _T_1952 <= _T_1949;
    end
    if (reset) begin
      _T_1955 <= 1'h0;
    end else begin
      _T_1955 <= _T_1952;
    end
    if (reset) begin
      _T_1958 <= 1'h0;
    end else begin
      _T_1958 <= _T_1955;
    end
    if (reset) begin
      _T_1963 <= 29'h0;
    end else begin
      if (_T_1788) begin
        _T_1963 <= _T_1938;
      end
    end
    if (reset) begin
      _T_1966 <= 29'h0;
    end else begin
      if (_T_1943) begin
        _T_1966 <= _T_1963;
      end
    end
    if (reset) begin
      _T_1969 <= 29'h0;
    end else begin
      if (_T_1946) begin
        _T_1969 <= _T_1966;
      end
    end
    if (reset) begin
      _T_1972 <= 29'h0;
    end else begin
      if (_T_1949) begin
        _T_1972 <= _T_1969;
      end
    end
    if (reset) begin
      _T_1975 <= 29'h0;
    end else begin
      if (_T_1952) begin
        _T_1975 <= _T_1972;
      end
    end
    if (reset) begin
      _T_1978 <= 29'h0;
    end else begin
      if (_T_1955) begin
        _T_1978 <= _T_1975;
      end
    end
    if (reset) begin
      _T_2051 <= 1'h1;
    end else begin
      if (io_sc2buf_dat_rd_data_valid) begin
        _T_2051 <= 1'h0;
      end
    end
    if (reset) begin
      _T_2063 <= 1'h1;
    end else begin
      if (_T_2108) begin
        _T_2063 <= 1'h0;
      end else begin
        if (io_sc2buf_dat_rd_data_valid) begin
          _T_2063 <= _T_2051;
        end
      end
    end
    if (io_sc2buf_dat_rd_data_valid) begin
      _T_2074 <= io_sc2buf_dat_rd_data_bits;
    end
    if (_T_2108) begin
      _T_2082 <= _T_2074;
    end
    if (reset) begin
      _T_2182 <= 8'h0;
    end else begin
      if (_T_2388) begin
        if (_T_630) begin
          _T_2182 <= 8'h40;
        end else begin
          if (_T_2344) begin
            _T_2182 <= _T_2194;
          end else begin
            if (_T_2345) begin
              _T_2182 <= 8'h40;
            end else begin
              if (_T_2307) begin
                _T_2182 <= 8'h40;
              end else begin
                _T_2182 <= _T_2313;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2185 <= 8'h0;
    end else begin
      if (_T_2394) begin
        if (_T_630) begin
          _T_2185 <= 8'h40;
        end else begin
          if (_T_2355) begin
            _T_2185 <= _T_2197;
          end else begin
            if (_T_2356) begin
              _T_2185 <= 8'h40;
            end else begin
              if (_T_2307) begin
                _T_2185 <= 8'h40;
              end else begin
                _T_2185 <= _T_2322;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2188 <= 8'h0;
    end else begin
      if (_T_2400) begin
        if (_T_630) begin
          _T_2188 <= 8'h40;
        end else begin
          if (_T_2366) begin
            _T_2188 <= _T_2200;
          end else begin
            if (_T_2367) begin
              _T_2188 <= 8'h40;
            end else begin
              if (_T_2307) begin
                _T_2188 <= 8'h40;
              end else begin
                _T_2188 <= _T_2331;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2191 <= 8'h0;
    end else begin
      if (_T_2406) begin
        if (_T_630) begin
          _T_2191 <= 8'h40;
        end else begin
          if (_T_2377) begin
            _T_2191 <= _T_2203;
          end else begin
            if (_T_2378) begin
              _T_2191 <= 8'h40;
            end else begin
              if (_T_2307) begin
                _T_2191 <= 8'h40;
              end else begin
                _T_2191 <= _T_2340;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2194 <= 8'h0;
    end else begin
      if (_T_2411) begin
        if (_T_630) begin
          _T_2194 <= 8'h40;
        end else begin
          if (!(_T_2344)) begin
            if (_T_2345) begin
              _T_2194 <= 8'h40;
            end else begin
              if (_T_2307) begin
                _T_2194 <= 8'h40;
              end else begin
                _T_2194 <= _T_2313;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2197 <= 8'h0;
    end else begin
      if (_T_2419) begin
        if (_T_630) begin
          _T_2197 <= 8'h40;
        end else begin
          if (!(_T_2355)) begin
            if (_T_2356) begin
              _T_2197 <= 8'h40;
            end else begin
              if (_T_2307) begin
                _T_2197 <= 8'h40;
              end else begin
                _T_2197 <= _T_2322;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2200 <= 8'h0;
    end else begin
      if (_T_2427) begin
        if (_T_630) begin
          _T_2200 <= 8'h40;
        end else begin
          if (!(_T_2366)) begin
            if (_T_2367) begin
              _T_2200 <= 8'h40;
            end else begin
              if (_T_2307) begin
                _T_2200 <= 8'h40;
              end else begin
                _T_2200 <= _T_2331;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2203 <= 8'h0;
    end else begin
      if (_T_2435) begin
        if (_T_630) begin
          _T_2203 <= 8'h40;
        end else begin
          if (!(_T_2377)) begin
            if (_T_2378) begin
              _T_2203 <= 8'h40;
            end else begin
              if (_T_2307) begin
                _T_2203 <= 8'h40;
              end else begin
                _T_2203 <= _T_2340;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2214 <= 1'h0;
    end else begin
      _T_2214 <= _T_2211;
    end
    if (reset) begin
      _T_2228 <= 27'h0;
    end else begin
      if (_T_2211) begin
        _T_2228 <= _T_2225;
      end
    end
    _T_2611 <= _GEN_149[255:0];
    _T_2613 <= _GEN_150[127:0];
    if (_T_2821) begin
      _T_2615 <= _T_2613;
    end
    _T_2617 <= _GEN_151[127:0];
    if (_T_2821) begin
      _T_2619 <= _T_2617;
    end
    _T_2621 <= _GEN_154[127:0];
    if (reset) begin
      _T_3419 <= 1'h0;
    end else begin
      _T_3419 <= _T_2248;
    end
    if (reset) begin
      _T_3689_0 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_0 <= _T_3220;
      end
    end
    if (reset) begin
      _T_3689_1 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_1 <= _T_3222;
      end
    end
    if (reset) begin
      _T_3689_2 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_2 <= _T_3224;
      end
    end
    if (reset) begin
      _T_3689_3 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_3 <= _T_3226;
      end
    end
    if (reset) begin
      _T_3689_4 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_4 <= _T_3228;
      end
    end
    if (reset) begin
      _T_3689_5 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_5 <= _T_3230;
      end
    end
    if (reset) begin
      _T_3689_6 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_6 <= _T_3232;
      end
    end
    if (reset) begin
      _T_3689_7 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_7 <= _T_3234;
      end
    end
    if (reset) begin
      _T_3689_8 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_8 <= _T_3236;
      end
    end
    if (reset) begin
      _T_3689_9 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_9 <= _T_3238;
      end
    end
    if (reset) begin
      _T_3689_10 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_10 <= _T_3240;
      end
    end
    if (reset) begin
      _T_3689_11 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_11 <= _T_3242;
      end
    end
    if (reset) begin
      _T_3689_12 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_12 <= _T_3244;
      end
    end
    if (reset) begin
      _T_3689_13 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_13 <= _T_3246;
      end
    end
    if (reset) begin
      _T_3689_14 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_14 <= _T_3248;
      end
    end
    if (reset) begin
      _T_3689_15 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_15 <= _T_3250;
      end
    end
    if (reset) begin
      _T_3689_16 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_16 <= _T_3252;
      end
    end
    if (reset) begin
      _T_3689_17 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_17 <= _T_3254;
      end
    end
    if (reset) begin
      _T_3689_18 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_18 <= _T_3256;
      end
    end
    if (reset) begin
      _T_3689_19 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_19 <= _T_3258;
      end
    end
    if (reset) begin
      _T_3689_20 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_20 <= _T_3260;
      end
    end
    if (reset) begin
      _T_3689_21 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_21 <= _T_3262;
      end
    end
    if (reset) begin
      _T_3689_22 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_22 <= _T_3264;
      end
    end
    if (reset) begin
      _T_3689_23 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_23 <= _T_3266;
      end
    end
    if (reset) begin
      _T_3689_24 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_24 <= _T_3268;
      end
    end
    if (reset) begin
      _T_3689_25 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_25 <= _T_3270;
      end
    end
    if (reset) begin
      _T_3689_26 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_26 <= _T_3272;
      end
    end
    if (reset) begin
      _T_3689_27 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_27 <= _T_3274;
      end
    end
    if (reset) begin
      _T_3689_28 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_28 <= _T_3276;
      end
    end
    if (reset) begin
      _T_3689_29 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_29 <= _T_3278;
      end
    end
    if (reset) begin
      _T_3689_30 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_30 <= _T_3280;
      end
    end
    if (reset) begin
      _T_3689_31 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_31 <= _T_3282;
      end
    end
    if (reset) begin
      _T_3689_32 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_32 <= _T_3284;
      end
    end
    if (reset) begin
      _T_3689_33 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_33 <= _T_3286;
      end
    end
    if (reset) begin
      _T_3689_34 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_34 <= _T_3288;
      end
    end
    if (reset) begin
      _T_3689_35 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_35 <= _T_3290;
      end
    end
    if (reset) begin
      _T_3689_36 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_36 <= _T_3292;
      end
    end
    if (reset) begin
      _T_3689_37 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_37 <= _T_3294;
      end
    end
    if (reset) begin
      _T_3689_38 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_38 <= _T_3296;
      end
    end
    if (reset) begin
      _T_3689_39 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_39 <= _T_3298;
      end
    end
    if (reset) begin
      _T_3689_40 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_40 <= _T_3300;
      end
    end
    if (reset) begin
      _T_3689_41 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_41 <= _T_3302;
      end
    end
    if (reset) begin
      _T_3689_42 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_42 <= _T_3304;
      end
    end
    if (reset) begin
      _T_3689_43 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_43 <= _T_3306;
      end
    end
    if (reset) begin
      _T_3689_44 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_44 <= _T_3308;
      end
    end
    if (reset) begin
      _T_3689_45 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_45 <= _T_3310;
      end
    end
    if (reset) begin
      _T_3689_46 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_46 <= _T_3312;
      end
    end
    if (reset) begin
      _T_3689_47 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_47 <= _T_3314;
      end
    end
    if (reset) begin
      _T_3689_48 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_48 <= _T_3316;
      end
    end
    if (reset) begin
      _T_3689_49 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_49 <= _T_3318;
      end
    end
    if (reset) begin
      _T_3689_50 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_50 <= _T_3320;
      end
    end
    if (reset) begin
      _T_3689_51 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_51 <= _T_3322;
      end
    end
    if (reset) begin
      _T_3689_52 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_52 <= _T_3324;
      end
    end
    if (reset) begin
      _T_3689_53 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_53 <= _T_3326;
      end
    end
    if (reset) begin
      _T_3689_54 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_54 <= _T_3328;
      end
    end
    if (reset) begin
      _T_3689_55 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_55 <= _T_3330;
      end
    end
    if (reset) begin
      _T_3689_56 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_56 <= _T_3332;
      end
    end
    if (reset) begin
      _T_3689_57 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_57 <= _T_3334;
      end
    end
    if (reset) begin
      _T_3689_58 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_58 <= _T_3336;
      end
    end
    if (reset) begin
      _T_3689_59 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_59 <= _T_3338;
      end
    end
    if (reset) begin
      _T_3689_60 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_60 <= _T_3340;
      end
    end
    if (reset) begin
      _T_3689_61 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_61 <= _T_3342;
      end
    end
    if (reset) begin
      _T_3689_62 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_62 <= _T_3344;
      end
    end
    if (reset) begin
      _T_3689_63 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_63 <= _T_3346;
      end
    end
    if (_T_3956) begin
      if (_T_2888) begin
        _T_3889_0 <= _T_2749;
      end else begin
        _T_3889_0 <= _T_2546;
      end
    end
    if (_T_3957) begin
      if (_T_2888) begin
        _T_3889_1 <= _T_2750;
      end else begin
        _T_3889_1 <= _T_2547;
      end
    end
    if (_T_3958) begin
      if (_T_2888) begin
        _T_3889_2 <= _T_2751;
      end else begin
        _T_3889_2 <= _T_2548;
      end
    end
    if (_T_3959) begin
      if (_T_2888) begin
        _T_3889_3 <= _T_2752;
      end else begin
        _T_3889_3 <= _T_2549;
      end
    end
    if (_T_3960) begin
      if (_T_2888) begin
        _T_3889_4 <= _T_2753;
      end else begin
        _T_3889_4 <= _T_2550;
      end
    end
    if (_T_3961) begin
      if (_T_2888) begin
        _T_3889_5 <= _T_2754;
      end else begin
        _T_3889_5 <= _T_2551;
      end
    end
    if (_T_3962) begin
      if (_T_2888) begin
        _T_3889_6 <= _T_2755;
      end else begin
        _T_3889_6 <= _T_2552;
      end
    end
    if (_T_3963) begin
      if (_T_2888) begin
        _T_3889_7 <= _T_2756;
      end else begin
        _T_3889_7 <= _T_2553;
      end
    end
    if (_T_3964) begin
      if (_T_2888) begin
        _T_3889_8 <= _T_2757;
      end else begin
        _T_3889_8 <= _T_2554;
      end
    end
    if (_T_3965) begin
      if (_T_2888) begin
        _T_3889_9 <= _T_2758;
      end else begin
        _T_3889_9 <= _T_2555;
      end
    end
    if (_T_3966) begin
      if (_T_2888) begin
        _T_3889_10 <= _T_2759;
      end else begin
        _T_3889_10 <= _T_2556;
      end
    end
    if (_T_3967) begin
      if (_T_2888) begin
        _T_3889_11 <= _T_2760;
      end else begin
        _T_3889_11 <= _T_2557;
      end
    end
    if (_T_3968) begin
      if (_T_2888) begin
        _T_3889_12 <= _T_2761;
      end else begin
        _T_3889_12 <= _T_2558;
      end
    end
    if (_T_3969) begin
      if (_T_2888) begin
        _T_3889_13 <= _T_2762;
      end else begin
        _T_3889_13 <= _T_2559;
      end
    end
    if (_T_3970) begin
      if (_T_2888) begin
        _T_3889_14 <= _T_2763;
      end else begin
        _T_3889_14 <= _T_2560;
      end
    end
    if (_T_3971) begin
      if (_T_2888) begin
        _T_3889_15 <= _T_2764;
      end else begin
        _T_3889_15 <= _T_2561;
      end
    end
    if (_T_3972) begin
      if (_T_2888) begin
        _T_3889_16 <= _T_2765;
      end else begin
        _T_3889_16 <= _T_2562;
      end
    end
    if (_T_3973) begin
      if (_T_2888) begin
        _T_3889_17 <= _T_2766;
      end else begin
        _T_3889_17 <= _T_2563;
      end
    end
    if (_T_3974) begin
      if (_T_2888) begin
        _T_3889_18 <= _T_2767;
      end else begin
        _T_3889_18 <= _T_2564;
      end
    end
    if (_T_3975) begin
      if (_T_2888) begin
        _T_3889_19 <= _T_2768;
      end else begin
        _T_3889_19 <= _T_2565;
      end
    end
    if (_T_3976) begin
      if (_T_2888) begin
        _T_3889_20 <= _T_2769;
      end else begin
        _T_3889_20 <= _T_2566;
      end
    end
    if (_T_3977) begin
      if (_T_2888) begin
        _T_3889_21 <= _T_2770;
      end else begin
        _T_3889_21 <= _T_2567;
      end
    end
    if (_T_3978) begin
      if (_T_2888) begin
        _T_3889_22 <= _T_2771;
      end else begin
        _T_3889_22 <= _T_2568;
      end
    end
    if (_T_3979) begin
      if (_T_2888) begin
        _T_3889_23 <= _T_2772;
      end else begin
        _T_3889_23 <= _T_2569;
      end
    end
    if (_T_3980) begin
      if (_T_2888) begin
        _T_3889_24 <= _T_2773;
      end else begin
        _T_3889_24 <= _T_2570;
      end
    end
    if (_T_3981) begin
      if (_T_2888) begin
        _T_3889_25 <= _T_2774;
      end else begin
        _T_3889_25 <= _T_2571;
      end
    end
    if (_T_3982) begin
      if (_T_2888) begin
        _T_3889_26 <= _T_2775;
      end else begin
        _T_3889_26 <= _T_2572;
      end
    end
    if (_T_3983) begin
      if (_T_2888) begin
        _T_3889_27 <= _T_2776;
      end else begin
        _T_3889_27 <= _T_2573;
      end
    end
    if (_T_3984) begin
      if (_T_2888) begin
        _T_3889_28 <= _T_2777;
      end else begin
        _T_3889_28 <= _T_2574;
      end
    end
    if (_T_3985) begin
      if (_T_2888) begin
        _T_3889_29 <= _T_2778;
      end else begin
        _T_3889_29 <= _T_2575;
      end
    end
    if (_T_3986) begin
      if (_T_2888) begin
        _T_3889_30 <= _T_2779;
      end else begin
        _T_3889_30 <= _T_2576;
      end
    end
    if (_T_3987) begin
      if (_T_2888) begin
        _T_3889_31 <= _T_2780;
      end else begin
        _T_3889_31 <= _T_2577;
      end
    end
    if (_T_3988) begin
      if (_T_2888) begin
        _T_3889_32 <= _T_2781;
      end else begin
        _T_3889_32 <= _T_2578;
      end
    end
    if (_T_3989) begin
      if (_T_2888) begin
        _T_3889_33 <= _T_2782;
      end else begin
        _T_3889_33 <= _T_2579;
      end
    end
    if (_T_3990) begin
      if (_T_2888) begin
        _T_3889_34 <= _T_2783;
      end else begin
        _T_3889_34 <= _T_2580;
      end
    end
    if (_T_3991) begin
      if (_T_2888) begin
        _T_3889_35 <= _T_2784;
      end else begin
        _T_3889_35 <= _T_2581;
      end
    end
    if (_T_3992) begin
      if (_T_2888) begin
        _T_3889_36 <= _T_2785;
      end else begin
        _T_3889_36 <= _T_2582;
      end
    end
    if (_T_3993) begin
      if (_T_2888) begin
        _T_3889_37 <= _T_2786;
      end else begin
        _T_3889_37 <= _T_2583;
      end
    end
    if (_T_3994) begin
      if (_T_2888) begin
        _T_3889_38 <= _T_2787;
      end else begin
        _T_3889_38 <= _T_2584;
      end
    end
    if (_T_3995) begin
      if (_T_2888) begin
        _T_3889_39 <= _T_2788;
      end else begin
        _T_3889_39 <= _T_2585;
      end
    end
    if (_T_3996) begin
      if (_T_2888) begin
        _T_3889_40 <= _T_2789;
      end else begin
        _T_3889_40 <= _T_2586;
      end
    end
    if (_T_3997) begin
      if (_T_2888) begin
        _T_3889_41 <= _T_2790;
      end else begin
        _T_3889_41 <= _T_2587;
      end
    end
    if (_T_3998) begin
      if (_T_2888) begin
        _T_3889_42 <= _T_2791;
      end else begin
        _T_3889_42 <= _T_2588;
      end
    end
    if (_T_3999) begin
      if (_T_2888) begin
        _T_3889_43 <= _T_2792;
      end else begin
        _T_3889_43 <= _T_2589;
      end
    end
    if (_T_4000) begin
      if (_T_2888) begin
        _T_3889_44 <= _T_2793;
      end else begin
        _T_3889_44 <= _T_2590;
      end
    end
    if (_T_4001) begin
      if (_T_2888) begin
        _T_3889_45 <= _T_2794;
      end else begin
        _T_3889_45 <= _T_2591;
      end
    end
    if (_T_4002) begin
      if (_T_2888) begin
        _T_3889_46 <= _T_2795;
      end else begin
        _T_3889_46 <= _T_2592;
      end
    end
    if (_T_4003) begin
      if (_T_2888) begin
        _T_3889_47 <= _T_2796;
      end else begin
        _T_3889_47 <= _T_2593;
      end
    end
    if (_T_4004) begin
      if (_T_2888) begin
        _T_3889_48 <= _T_2797;
      end else begin
        _T_3889_48 <= _T_2594;
      end
    end
    if (_T_4005) begin
      if (_T_2888) begin
        _T_3889_49 <= _T_2798;
      end else begin
        _T_3889_49 <= _T_2595;
      end
    end
    if (_T_4006) begin
      if (_T_2888) begin
        _T_3889_50 <= _T_2799;
      end else begin
        _T_3889_50 <= _T_2596;
      end
    end
    if (_T_4007) begin
      if (_T_2888) begin
        _T_3889_51 <= _T_2800;
      end else begin
        _T_3889_51 <= _T_2597;
      end
    end
    if (_T_4008) begin
      if (_T_2888) begin
        _T_3889_52 <= _T_2801;
      end else begin
        _T_3889_52 <= _T_2598;
      end
    end
    if (_T_4009) begin
      if (_T_2888) begin
        _T_3889_53 <= _T_2802;
      end else begin
        _T_3889_53 <= _T_2599;
      end
    end
    if (_T_4010) begin
      if (_T_2888) begin
        _T_3889_54 <= _T_2803;
      end else begin
        _T_3889_54 <= _T_2600;
      end
    end
    if (_T_4011) begin
      if (_T_2888) begin
        _T_3889_55 <= _T_2804;
      end else begin
        _T_3889_55 <= _T_2601;
      end
    end
    if (_T_4012) begin
      if (_T_2888) begin
        _T_3889_56 <= _T_2805;
      end else begin
        _T_3889_56 <= _T_2602;
      end
    end
    if (_T_4013) begin
      if (_T_2888) begin
        _T_3889_57 <= _T_2806;
      end else begin
        _T_3889_57 <= _T_2603;
      end
    end
    if (_T_4014) begin
      if (_T_2888) begin
        _T_3889_58 <= _T_2807;
      end else begin
        _T_3889_58 <= _T_2604;
      end
    end
    if (_T_4015) begin
      if (_T_2888) begin
        _T_3889_59 <= _T_2808;
      end else begin
        _T_3889_59 <= _T_2605;
      end
    end
    if (_T_4016) begin
      if (_T_2888) begin
        _T_3889_60 <= _T_2809;
      end else begin
        _T_3889_60 <= _T_2606;
      end
    end
    if (_T_4017) begin
      if (_T_2888) begin
        _T_3889_61 <= _T_2810;
      end else begin
        _T_3889_61 <= _T_2607;
      end
    end
    if (_T_4018) begin
      if (_T_2888) begin
        _T_3889_62 <= _T_2811;
      end else begin
        _T_3889_62 <= _T_2608;
      end
    end
    if (_T_4019) begin
      if (_T_2888) begin
        _T_3889_63 <= _T_2812;
      end else begin
        _T_3889_63 <= _T_2609;
      end
    end
    if (reset) begin
      _T_4022 <= 1'h0;
    end else begin
      _T_4022 <= _T_3419;
    end
    if (reset) begin
      _T_4289_0 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_0 <= 1'h0;
        end else begin
          _T_4289_0 <= _T_3689_0;
        end
      end
    end
    if (reset) begin
      _T_4289_1 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_1 <= 1'h0;
        end else begin
          _T_4289_1 <= _T_3689_1;
        end
      end
    end
    if (reset) begin
      _T_4289_2 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_2 <= 1'h0;
        end else begin
          _T_4289_2 <= _T_3689_2;
        end
      end
    end
    if (reset) begin
      _T_4289_3 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_3 <= 1'h0;
        end else begin
          _T_4289_3 <= _T_3689_3;
        end
      end
    end
    if (reset) begin
      _T_4289_4 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_4 <= 1'h0;
        end else begin
          _T_4289_4 <= _T_3689_4;
        end
      end
    end
    if (reset) begin
      _T_4289_5 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_5 <= 1'h0;
        end else begin
          _T_4289_5 <= _T_3689_5;
        end
      end
    end
    if (reset) begin
      _T_4289_6 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_6 <= 1'h0;
        end else begin
          _T_4289_6 <= _T_3689_6;
        end
      end
    end
    if (reset) begin
      _T_4289_7 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_7 <= 1'h0;
        end else begin
          _T_4289_7 <= _T_3689_7;
        end
      end
    end
    if (reset) begin
      _T_4289_8 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_8 <= 1'h0;
        end else begin
          _T_4289_8 <= _T_3689_8;
        end
      end
    end
    if (reset) begin
      _T_4289_9 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_9 <= 1'h0;
        end else begin
          _T_4289_9 <= _T_3689_9;
        end
      end
    end
    if (reset) begin
      _T_4289_10 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_10 <= 1'h0;
        end else begin
          _T_4289_10 <= _T_3689_10;
        end
      end
    end
    if (reset) begin
      _T_4289_11 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_11 <= 1'h0;
        end else begin
          _T_4289_11 <= _T_3689_11;
        end
      end
    end
    if (reset) begin
      _T_4289_12 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_12 <= 1'h0;
        end else begin
          _T_4289_12 <= _T_3689_12;
        end
      end
    end
    if (reset) begin
      _T_4289_13 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_13 <= 1'h0;
        end else begin
          _T_4289_13 <= _T_3689_13;
        end
      end
    end
    if (reset) begin
      _T_4289_14 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_14 <= 1'h0;
        end else begin
          _T_4289_14 <= _T_3689_14;
        end
      end
    end
    if (reset) begin
      _T_4289_15 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_15 <= 1'h0;
        end else begin
          _T_4289_15 <= _T_3689_15;
        end
      end
    end
    if (reset) begin
      _T_4289_16 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_16 <= 1'h0;
        end else begin
          _T_4289_16 <= _T_3689_16;
        end
      end
    end
    if (reset) begin
      _T_4289_17 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_17 <= 1'h0;
        end else begin
          _T_4289_17 <= _T_3689_17;
        end
      end
    end
    if (reset) begin
      _T_4289_18 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_18 <= 1'h0;
        end else begin
          _T_4289_18 <= _T_3689_18;
        end
      end
    end
    if (reset) begin
      _T_4289_19 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_19 <= 1'h0;
        end else begin
          _T_4289_19 <= _T_3689_19;
        end
      end
    end
    if (reset) begin
      _T_4289_20 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_20 <= 1'h0;
        end else begin
          _T_4289_20 <= _T_3689_20;
        end
      end
    end
    if (reset) begin
      _T_4289_21 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_21 <= 1'h0;
        end else begin
          _T_4289_21 <= _T_3689_21;
        end
      end
    end
    if (reset) begin
      _T_4289_22 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_22 <= 1'h0;
        end else begin
          _T_4289_22 <= _T_3689_22;
        end
      end
    end
    if (reset) begin
      _T_4289_23 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_23 <= 1'h0;
        end else begin
          _T_4289_23 <= _T_3689_23;
        end
      end
    end
    if (reset) begin
      _T_4289_24 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_24 <= 1'h0;
        end else begin
          _T_4289_24 <= _T_3689_24;
        end
      end
    end
    if (reset) begin
      _T_4289_25 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_25 <= 1'h0;
        end else begin
          _T_4289_25 <= _T_3689_25;
        end
      end
    end
    if (reset) begin
      _T_4289_26 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_26 <= 1'h0;
        end else begin
          _T_4289_26 <= _T_3689_26;
        end
      end
    end
    if (reset) begin
      _T_4289_27 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_27 <= 1'h0;
        end else begin
          _T_4289_27 <= _T_3689_27;
        end
      end
    end
    if (reset) begin
      _T_4289_28 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_28 <= 1'h0;
        end else begin
          _T_4289_28 <= _T_3689_28;
        end
      end
    end
    if (reset) begin
      _T_4289_29 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_29 <= 1'h0;
        end else begin
          _T_4289_29 <= _T_3689_29;
        end
      end
    end
    if (reset) begin
      _T_4289_30 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_30 <= 1'h0;
        end else begin
          _T_4289_30 <= _T_3689_30;
        end
      end
    end
    if (reset) begin
      _T_4289_31 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_31 <= 1'h0;
        end else begin
          _T_4289_31 <= _T_3689_31;
        end
      end
    end
    if (reset) begin
      _T_4289_32 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_32 <= 1'h0;
        end else begin
          _T_4289_32 <= _T_3689_32;
        end
      end
    end
    if (reset) begin
      _T_4289_33 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_33 <= 1'h0;
        end else begin
          _T_4289_33 <= _T_3689_33;
        end
      end
    end
    if (reset) begin
      _T_4289_34 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_34 <= 1'h0;
        end else begin
          _T_4289_34 <= _T_3689_34;
        end
      end
    end
    if (reset) begin
      _T_4289_35 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_35 <= 1'h0;
        end else begin
          _T_4289_35 <= _T_3689_35;
        end
      end
    end
    if (reset) begin
      _T_4289_36 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_36 <= 1'h0;
        end else begin
          _T_4289_36 <= _T_3689_36;
        end
      end
    end
    if (reset) begin
      _T_4289_37 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_37 <= 1'h0;
        end else begin
          _T_4289_37 <= _T_3689_37;
        end
      end
    end
    if (reset) begin
      _T_4289_38 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_38 <= 1'h0;
        end else begin
          _T_4289_38 <= _T_3689_38;
        end
      end
    end
    if (reset) begin
      _T_4289_39 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_39 <= 1'h0;
        end else begin
          _T_4289_39 <= _T_3689_39;
        end
      end
    end
    if (reset) begin
      _T_4289_40 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_40 <= 1'h0;
        end else begin
          _T_4289_40 <= _T_3689_40;
        end
      end
    end
    if (reset) begin
      _T_4289_41 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_41 <= 1'h0;
        end else begin
          _T_4289_41 <= _T_3689_41;
        end
      end
    end
    if (reset) begin
      _T_4289_42 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_42 <= 1'h0;
        end else begin
          _T_4289_42 <= _T_3689_42;
        end
      end
    end
    if (reset) begin
      _T_4289_43 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_43 <= 1'h0;
        end else begin
          _T_4289_43 <= _T_3689_43;
        end
      end
    end
    if (reset) begin
      _T_4289_44 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_44 <= 1'h0;
        end else begin
          _T_4289_44 <= _T_3689_44;
        end
      end
    end
    if (reset) begin
      _T_4289_45 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_45 <= 1'h0;
        end else begin
          _T_4289_45 <= _T_3689_45;
        end
      end
    end
    if (reset) begin
      _T_4289_46 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_46 <= 1'h0;
        end else begin
          _T_4289_46 <= _T_3689_46;
        end
      end
    end
    if (reset) begin
      _T_4289_47 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_47 <= 1'h0;
        end else begin
          _T_4289_47 <= _T_3689_47;
        end
      end
    end
    if (reset) begin
      _T_4289_48 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_48 <= 1'h0;
        end else begin
          _T_4289_48 <= _T_3689_48;
        end
      end
    end
    if (reset) begin
      _T_4289_49 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_49 <= 1'h0;
        end else begin
          _T_4289_49 <= _T_3689_49;
        end
      end
    end
    if (reset) begin
      _T_4289_50 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_50 <= 1'h0;
        end else begin
          _T_4289_50 <= _T_3689_50;
        end
      end
    end
    if (reset) begin
      _T_4289_51 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_51 <= 1'h0;
        end else begin
          _T_4289_51 <= _T_3689_51;
        end
      end
    end
    if (reset) begin
      _T_4289_52 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_52 <= 1'h0;
        end else begin
          _T_4289_52 <= _T_3689_52;
        end
      end
    end
    if (reset) begin
      _T_4289_53 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_53 <= 1'h0;
        end else begin
          _T_4289_53 <= _T_3689_53;
        end
      end
    end
    if (reset) begin
      _T_4289_54 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_54 <= 1'h0;
        end else begin
          _T_4289_54 <= _T_3689_54;
        end
      end
    end
    if (reset) begin
      _T_4289_55 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_55 <= 1'h0;
        end else begin
          _T_4289_55 <= _T_3689_55;
        end
      end
    end
    if (reset) begin
      _T_4289_56 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_56 <= 1'h0;
        end else begin
          _T_4289_56 <= _T_3689_56;
        end
      end
    end
    if (reset) begin
      _T_4289_57 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_57 <= 1'h0;
        end else begin
          _T_4289_57 <= _T_3689_57;
        end
      end
    end
    if (reset) begin
      _T_4289_58 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_58 <= 1'h0;
        end else begin
          _T_4289_58 <= _T_3689_58;
        end
      end
    end
    if (reset) begin
      _T_4289_59 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_59 <= 1'h0;
        end else begin
          _T_4289_59 <= _T_3689_59;
        end
      end
    end
    if (reset) begin
      _T_4289_60 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_60 <= 1'h0;
        end else begin
          _T_4289_60 <= _T_3689_60;
        end
      end
    end
    if (reset) begin
      _T_4289_61 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_61 <= 1'h0;
        end else begin
          _T_4289_61 <= _T_3689_61;
        end
      end
    end
    if (reset) begin
      _T_4289_62 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_62 <= 1'h0;
        end else begin
          _T_4289_62 <= _T_3689_62;
        end
      end
    end
    if (reset) begin
      _T_4289_63 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_63 <= 1'h0;
        end else begin
          _T_4289_63 <= _T_3689_63;
        end
      end
    end
    if (reset) begin
      _T_4488 <= 9'h0;
    end else begin
      if (_T_3419) begin
        _T_4488 <= {{8'd0}, _T_3419};
      end
    end
    if (_T_4694_0) begin
      _T_4492_0 <= _T_3889_0;
    end
    if (_T_4694_1) begin
      _T_4492_1 <= _T_3889_1;
    end
    if (_T_4694_2) begin
      _T_4492_2 <= _T_3889_2;
    end
    if (_T_4694_3) begin
      _T_4492_3 <= _T_3889_3;
    end
    if (_T_4694_4) begin
      _T_4492_4 <= _T_3889_4;
    end
    if (_T_4694_5) begin
      _T_4492_5 <= _T_3889_5;
    end
    if (_T_4694_6) begin
      _T_4492_6 <= _T_3889_6;
    end
    if (_T_4694_7) begin
      _T_4492_7 <= _T_3889_7;
    end
    if (_T_4694_8) begin
      _T_4492_8 <= _T_3889_8;
    end
    if (_T_4694_9) begin
      _T_4492_9 <= _T_3889_9;
    end
    if (_T_4694_10) begin
      _T_4492_10 <= _T_3889_10;
    end
    if (_T_4694_11) begin
      _T_4492_11 <= _T_3889_11;
    end
    if (_T_4694_12) begin
      _T_4492_12 <= _T_3889_12;
    end
    if (_T_4694_13) begin
      _T_4492_13 <= _T_3889_13;
    end
    if (_T_4694_14) begin
      _T_4492_14 <= _T_3889_14;
    end
    if (_T_4694_15) begin
      _T_4492_15 <= _T_3889_15;
    end
    if (_T_4694_16) begin
      _T_4492_16 <= _T_3889_16;
    end
    if (_T_4694_17) begin
      _T_4492_17 <= _T_3889_17;
    end
    if (_T_4694_18) begin
      _T_4492_18 <= _T_3889_18;
    end
    if (_T_4694_19) begin
      _T_4492_19 <= _T_3889_19;
    end
    if (_T_4694_20) begin
      _T_4492_20 <= _T_3889_20;
    end
    if (_T_4694_21) begin
      _T_4492_21 <= _T_3889_21;
    end
    if (_T_4694_22) begin
      _T_4492_22 <= _T_3889_22;
    end
    if (_T_4694_23) begin
      _T_4492_23 <= _T_3889_23;
    end
    if (_T_4694_24) begin
      _T_4492_24 <= _T_3889_24;
    end
    if (_T_4694_25) begin
      _T_4492_25 <= _T_3889_25;
    end
    if (_T_4694_26) begin
      _T_4492_26 <= _T_3889_26;
    end
    if (_T_4694_27) begin
      _T_4492_27 <= _T_3889_27;
    end
    if (_T_4694_28) begin
      _T_4492_28 <= _T_3889_28;
    end
    if (_T_4694_29) begin
      _T_4492_29 <= _T_3889_29;
    end
    if (_T_4694_30) begin
      _T_4492_30 <= _T_3889_30;
    end
    if (_T_4694_31) begin
      _T_4492_31 <= _T_3889_31;
    end
    if (_T_4694_32) begin
      _T_4492_32 <= _T_3889_32;
    end
    if (_T_4694_33) begin
      _T_4492_33 <= _T_3889_33;
    end
    if (_T_4694_34) begin
      _T_4492_34 <= _T_3889_34;
    end
    if (_T_4694_35) begin
      _T_4492_35 <= _T_3889_35;
    end
    if (_T_4694_36) begin
      _T_4492_36 <= _T_3889_36;
    end
    if (_T_4694_37) begin
      _T_4492_37 <= _T_3889_37;
    end
    if (_T_4694_38) begin
      _T_4492_38 <= _T_3889_38;
    end
    if (_T_4694_39) begin
      _T_4492_39 <= _T_3889_39;
    end
    if (_T_4694_40) begin
      _T_4492_40 <= _T_3889_40;
    end
    if (_T_4694_41) begin
      _T_4492_41 <= _T_3889_41;
    end
    if (_T_4694_42) begin
      _T_4492_42 <= _T_3889_42;
    end
    if (_T_4694_43) begin
      _T_4492_43 <= _T_3889_43;
    end
    if (_T_4694_44) begin
      _T_4492_44 <= _T_3889_44;
    end
    if (_T_4694_45) begin
      _T_4492_45 <= _T_3889_45;
    end
    if (_T_4694_46) begin
      _T_4492_46 <= _T_3889_46;
    end
    if (_T_4694_47) begin
      _T_4492_47 <= _T_3889_47;
    end
    if (_T_4694_48) begin
      _T_4492_48 <= _T_3889_48;
    end
    if (_T_4694_49) begin
      _T_4492_49 <= _T_3889_49;
    end
    if (_T_4694_50) begin
      _T_4492_50 <= _T_3889_50;
    end
    if (_T_4694_51) begin
      _T_4492_51 <= _T_3889_51;
    end
    if (_T_4694_52) begin
      _T_4492_52 <= _T_3889_52;
    end
    if (_T_4694_53) begin
      _T_4492_53 <= _T_3889_53;
    end
    if (_T_4694_54) begin
      _T_4492_54 <= _T_3889_54;
    end
    if (_T_4694_55) begin
      _T_4492_55 <= _T_3889_55;
    end
    if (_T_4694_56) begin
      _T_4492_56 <= _T_3889_56;
    end
    if (_T_4694_57) begin
      _T_4492_57 <= _T_3889_57;
    end
    if (_T_4694_58) begin
      _T_4492_58 <= _T_3889_58;
    end
    if (_T_4694_59) begin
      _T_4492_59 <= _T_3889_59;
    end
    if (_T_4694_60) begin
      _T_4492_60 <= _T_3889_60;
    end
    if (_T_4694_61) begin
      _T_4492_61 <= _T_3889_61;
    end
    if (_T_4694_62) begin
      _T_4492_62 <= _T_3889_62;
    end
    if (_T_4694_63) begin
      _T_4492_63 <= _T_3889_63;
    end
    if (reset) begin
      _T_4829 <= 1'h0;
    end else begin
      _T_4829 <= _T_4022;
    end
    if (reset) begin
      _T_4835 <= 1'h0;
    end else begin
      _T_4835 <= _T_4022;
    end
    if (reset) begin
      _T_4838 <= 1'h0;
    end else begin
      _T_4838 <= _T_4022;
    end
    if (reset) begin
      _T_4842 <= 9'h0;
    end else begin
      if (_T_4840) begin
        if (_T_4830) begin
          _T_4842 <= 9'h0;
        end else begin
          _T_4842 <= _T_4488;
        end
      end
    end
    if (reset) begin
      _T_4846 <= 9'h0;
    end else begin
      if (_T_4840) begin
        if (_T_4830) begin
          _T_4846 <= 9'h0;
        end else begin
          _T_4846 <= _T_4488;
        end
      end
    end
    if (reset) begin
      _T_5114_0 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_0 <= _T_4289_0;
      end
    end
    if (reset) begin
      _T_5114_1 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_1 <= _T_4289_1;
      end
    end
    if (reset) begin
      _T_5114_2 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_2 <= _T_4289_2;
      end
    end
    if (reset) begin
      _T_5114_3 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_3 <= _T_4289_3;
      end
    end
    if (reset) begin
      _T_5114_4 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_4 <= _T_4289_4;
      end
    end
    if (reset) begin
      _T_5114_5 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_5 <= _T_4289_5;
      end
    end
    if (reset) begin
      _T_5114_6 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_6 <= _T_4289_6;
      end
    end
    if (reset) begin
      _T_5114_7 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_7 <= _T_4289_7;
      end
    end
    if (reset) begin
      _T_5114_8 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_8 <= _T_4289_8;
      end
    end
    if (reset) begin
      _T_5114_9 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_9 <= _T_4289_9;
      end
    end
    if (reset) begin
      _T_5114_10 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_10 <= _T_4289_10;
      end
    end
    if (reset) begin
      _T_5114_11 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_11 <= _T_4289_11;
      end
    end
    if (reset) begin
      _T_5114_12 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_12 <= _T_4289_12;
      end
    end
    if (reset) begin
      _T_5114_13 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_13 <= _T_4289_13;
      end
    end
    if (reset) begin
      _T_5114_14 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_14 <= _T_4289_14;
      end
    end
    if (reset) begin
      _T_5114_15 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_15 <= _T_4289_15;
      end
    end
    if (reset) begin
      _T_5114_16 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_16 <= _T_4289_16;
      end
    end
    if (reset) begin
      _T_5114_17 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_17 <= _T_4289_17;
      end
    end
    if (reset) begin
      _T_5114_18 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_18 <= _T_4289_18;
      end
    end
    if (reset) begin
      _T_5114_19 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_19 <= _T_4289_19;
      end
    end
    if (reset) begin
      _T_5114_20 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_20 <= _T_4289_20;
      end
    end
    if (reset) begin
      _T_5114_21 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_21 <= _T_4289_21;
      end
    end
    if (reset) begin
      _T_5114_22 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_22 <= _T_4289_22;
      end
    end
    if (reset) begin
      _T_5114_23 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_23 <= _T_4289_23;
      end
    end
    if (reset) begin
      _T_5114_24 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_24 <= _T_4289_24;
      end
    end
    if (reset) begin
      _T_5114_25 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_25 <= _T_4289_25;
      end
    end
    if (reset) begin
      _T_5114_26 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_26 <= _T_4289_26;
      end
    end
    if (reset) begin
      _T_5114_27 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_27 <= _T_4289_27;
      end
    end
    if (reset) begin
      _T_5114_28 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_28 <= _T_4289_28;
      end
    end
    if (reset) begin
      _T_5114_29 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_29 <= _T_4289_29;
      end
    end
    if (reset) begin
      _T_5114_30 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_30 <= _T_4289_30;
      end
    end
    if (reset) begin
      _T_5114_31 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_31 <= _T_4289_31;
      end
    end
    if (reset) begin
      _T_5114_32 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_32 <= _T_4289_32;
      end
    end
    if (reset) begin
      _T_5114_33 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_33 <= _T_4289_33;
      end
    end
    if (reset) begin
      _T_5114_34 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_34 <= _T_4289_34;
      end
    end
    if (reset) begin
      _T_5114_35 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_35 <= _T_4289_35;
      end
    end
    if (reset) begin
      _T_5114_36 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_36 <= _T_4289_36;
      end
    end
    if (reset) begin
      _T_5114_37 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_37 <= _T_4289_37;
      end
    end
    if (reset) begin
      _T_5114_38 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_38 <= _T_4289_38;
      end
    end
    if (reset) begin
      _T_5114_39 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_39 <= _T_4289_39;
      end
    end
    if (reset) begin
      _T_5114_40 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_40 <= _T_4289_40;
      end
    end
    if (reset) begin
      _T_5114_41 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_41 <= _T_4289_41;
      end
    end
    if (reset) begin
      _T_5114_42 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_42 <= _T_4289_42;
      end
    end
    if (reset) begin
      _T_5114_43 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_43 <= _T_4289_43;
      end
    end
    if (reset) begin
      _T_5114_44 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_44 <= _T_4289_44;
      end
    end
    if (reset) begin
      _T_5114_45 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_45 <= _T_4289_45;
      end
    end
    if (reset) begin
      _T_5114_46 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_46 <= _T_4289_46;
      end
    end
    if (reset) begin
      _T_5114_47 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_47 <= _T_4289_47;
      end
    end
    if (reset) begin
      _T_5114_48 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_48 <= _T_4289_48;
      end
    end
    if (reset) begin
      _T_5114_49 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_49 <= _T_4289_49;
      end
    end
    if (reset) begin
      _T_5114_50 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_50 <= _T_4289_50;
      end
    end
    if (reset) begin
      _T_5114_51 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_51 <= _T_4289_51;
      end
    end
    if (reset) begin
      _T_5114_52 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_52 <= _T_4289_52;
      end
    end
    if (reset) begin
      _T_5114_53 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_53 <= _T_4289_53;
      end
    end
    if (reset) begin
      _T_5114_54 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_54 <= _T_4289_54;
      end
    end
    if (reset) begin
      _T_5114_55 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_55 <= _T_4289_55;
      end
    end
    if (reset) begin
      _T_5114_56 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_56 <= _T_4289_56;
      end
    end
    if (reset) begin
      _T_5114_57 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_57 <= _T_4289_57;
      end
    end
    if (reset) begin
      _T_5114_58 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_58 <= _T_4289_58;
      end
    end
    if (reset) begin
      _T_5114_59 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_59 <= _T_4289_59;
      end
    end
    if (reset) begin
      _T_5114_60 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_60 <= _T_4289_60;
      end
    end
    if (reset) begin
      _T_5114_61 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_61 <= _T_4289_61;
      end
    end
    if (reset) begin
      _T_5114_62 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_62 <= _T_4289_62;
      end
    end
    if (reset) begin
      _T_5114_63 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_63 <= _T_4289_63;
      end
    end
    if (reset) begin
      _T_5578_0 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_0 <= _T_4289_0;
      end
    end
    if (reset) begin
      _T_5578_1 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_1 <= _T_4289_1;
      end
    end
    if (reset) begin
      _T_5578_2 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_2 <= _T_4289_2;
      end
    end
    if (reset) begin
      _T_5578_3 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_3 <= _T_4289_3;
      end
    end
    if (reset) begin
      _T_5578_4 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_4 <= _T_4289_4;
      end
    end
    if (reset) begin
      _T_5578_5 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_5 <= _T_4289_5;
      end
    end
    if (reset) begin
      _T_5578_6 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_6 <= _T_4289_6;
      end
    end
    if (reset) begin
      _T_5578_7 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_7 <= _T_4289_7;
      end
    end
    if (reset) begin
      _T_5578_8 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_8 <= _T_4289_8;
      end
    end
    if (reset) begin
      _T_5578_9 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_9 <= _T_4289_9;
      end
    end
    if (reset) begin
      _T_5578_10 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_10 <= _T_4289_10;
      end
    end
    if (reset) begin
      _T_5578_11 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_11 <= _T_4289_11;
      end
    end
    if (reset) begin
      _T_5578_12 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_12 <= _T_4289_12;
      end
    end
    if (reset) begin
      _T_5578_13 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_13 <= _T_4289_13;
      end
    end
    if (reset) begin
      _T_5578_14 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_14 <= _T_4289_14;
      end
    end
    if (reset) begin
      _T_5578_15 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_15 <= _T_4289_15;
      end
    end
    if (reset) begin
      _T_5578_16 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_16 <= _T_4289_16;
      end
    end
    if (reset) begin
      _T_5578_17 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_17 <= _T_4289_17;
      end
    end
    if (reset) begin
      _T_5578_18 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_18 <= _T_4289_18;
      end
    end
    if (reset) begin
      _T_5578_19 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_19 <= _T_4289_19;
      end
    end
    if (reset) begin
      _T_5578_20 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_20 <= _T_4289_20;
      end
    end
    if (reset) begin
      _T_5578_21 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_21 <= _T_4289_21;
      end
    end
    if (reset) begin
      _T_5578_22 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_22 <= _T_4289_22;
      end
    end
    if (reset) begin
      _T_5578_23 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_23 <= _T_4289_23;
      end
    end
    if (reset) begin
      _T_5578_24 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_24 <= _T_4289_24;
      end
    end
    if (reset) begin
      _T_5578_25 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_25 <= _T_4289_25;
      end
    end
    if (reset) begin
      _T_5578_26 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_26 <= _T_4289_26;
      end
    end
    if (reset) begin
      _T_5578_27 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_27 <= _T_4289_27;
      end
    end
    if (reset) begin
      _T_5578_28 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_28 <= _T_4289_28;
      end
    end
    if (reset) begin
      _T_5578_29 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_29 <= _T_4289_29;
      end
    end
    if (reset) begin
      _T_5578_30 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_30 <= _T_4289_30;
      end
    end
    if (reset) begin
      _T_5578_31 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_31 <= _T_4289_31;
      end
    end
    if (reset) begin
      _T_5578_32 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_32 <= _T_4289_32;
      end
    end
    if (reset) begin
      _T_5578_33 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_33 <= _T_4289_33;
      end
    end
    if (reset) begin
      _T_5578_34 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_34 <= _T_4289_34;
      end
    end
    if (reset) begin
      _T_5578_35 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_35 <= _T_4289_35;
      end
    end
    if (reset) begin
      _T_5578_36 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_36 <= _T_4289_36;
      end
    end
    if (reset) begin
      _T_5578_37 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_37 <= _T_4289_37;
      end
    end
    if (reset) begin
      _T_5578_38 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_38 <= _T_4289_38;
      end
    end
    if (reset) begin
      _T_5578_39 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_39 <= _T_4289_39;
      end
    end
    if (reset) begin
      _T_5578_40 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_40 <= _T_4289_40;
      end
    end
    if (reset) begin
      _T_5578_41 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_41 <= _T_4289_41;
      end
    end
    if (reset) begin
      _T_5578_42 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_42 <= _T_4289_42;
      end
    end
    if (reset) begin
      _T_5578_43 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_43 <= _T_4289_43;
      end
    end
    if (reset) begin
      _T_5578_44 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_44 <= _T_4289_44;
      end
    end
    if (reset) begin
      _T_5578_45 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_45 <= _T_4289_45;
      end
    end
    if (reset) begin
      _T_5578_46 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_46 <= _T_4289_46;
      end
    end
    if (reset) begin
      _T_5578_47 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_47 <= _T_4289_47;
      end
    end
    if (reset) begin
      _T_5578_48 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_48 <= _T_4289_48;
      end
    end
    if (reset) begin
      _T_5578_49 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_49 <= _T_4289_49;
      end
    end
    if (reset) begin
      _T_5578_50 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_50 <= _T_4289_50;
      end
    end
    if (reset) begin
      _T_5578_51 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_51 <= _T_4289_51;
      end
    end
    if (reset) begin
      _T_5578_52 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_52 <= _T_4289_52;
      end
    end
    if (reset) begin
      _T_5578_53 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_53 <= _T_4289_53;
      end
    end
    if (reset) begin
      _T_5578_54 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_54 <= _T_4289_54;
      end
    end
    if (reset) begin
      _T_5578_55 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_55 <= _T_4289_55;
      end
    end
    if (reset) begin
      _T_5578_56 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_56 <= _T_4289_56;
      end
    end
    if (reset) begin
      _T_5578_57 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_57 <= _T_4289_57;
      end
    end
    if (reset) begin
      _T_5578_58 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_58 <= _T_4289_58;
      end
    end
    if (reset) begin
      _T_5578_59 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_59 <= _T_4289_59;
      end
    end
    if (reset) begin
      _T_5578_60 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_60 <= _T_4289_60;
      end
    end
    if (reset) begin
      _T_5578_61 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_61 <= _T_4289_61;
      end
    end
    if (reset) begin
      _T_5578_62 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_62 <= _T_4289_62;
      end
    end
    if (reset) begin
      _T_5578_63 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_63 <= _T_4289_63;
      end
    end
    if (_T_4289_0) begin
      _T_5776 <= _T_4492_0;
    end
    if (_T_4289_0) begin
      _T_5778 <= _T_4492_0;
    end
    if (_T_4289_1) begin
      _T_5780 <= _T_4492_1;
    end
    if (_T_4289_1) begin
      _T_5782 <= _T_4492_1;
    end
    if (_T_4289_2) begin
      _T_5784 <= _T_4492_2;
    end
    if (_T_4289_2) begin
      _T_5786 <= _T_4492_2;
    end
    if (_T_4289_3) begin
      _T_5788 <= _T_4492_3;
    end
    if (_T_4289_3) begin
      _T_5790 <= _T_4492_3;
    end
    if (_T_4289_4) begin
      _T_5792 <= _T_4492_4;
    end
    if (_T_4289_4) begin
      _T_5794 <= _T_4492_4;
    end
    if (_T_4289_5) begin
      _T_5796 <= _T_4492_5;
    end
    if (_T_4289_5) begin
      _T_5798 <= _T_4492_5;
    end
    if (_T_4289_6) begin
      _T_5800 <= _T_4492_6;
    end
    if (_T_4289_6) begin
      _T_5802 <= _T_4492_6;
    end
    if (_T_4289_7) begin
      _T_5804 <= _T_4492_7;
    end
    if (_T_4289_7) begin
      _T_5806 <= _T_4492_7;
    end
    if (_T_4289_8) begin
      _T_5808 <= _T_4492_8;
    end
    if (_T_4289_8) begin
      _T_5810 <= _T_4492_8;
    end
    if (_T_4289_9) begin
      _T_5812 <= _T_4492_9;
    end
    if (_T_4289_9) begin
      _T_5814 <= _T_4492_9;
    end
    if (_T_4289_10) begin
      _T_5816 <= _T_4492_10;
    end
    if (_T_4289_10) begin
      _T_5818 <= _T_4492_10;
    end
    if (_T_4289_11) begin
      _T_5820 <= _T_4492_11;
    end
    if (_T_4289_11) begin
      _T_5822 <= _T_4492_11;
    end
    if (_T_4289_12) begin
      _T_5824 <= _T_4492_12;
    end
    if (_T_4289_12) begin
      _T_5826 <= _T_4492_12;
    end
    if (_T_4289_13) begin
      _T_5828 <= _T_4492_13;
    end
    if (_T_4289_13) begin
      _T_5830 <= _T_4492_13;
    end
    if (_T_4289_14) begin
      _T_5832 <= _T_4492_14;
    end
    if (_T_4289_14) begin
      _T_5834 <= _T_4492_14;
    end
    if (_T_4289_15) begin
      _T_5836 <= _T_4492_15;
    end
    if (_T_4289_15) begin
      _T_5838 <= _T_4492_15;
    end
    if (_T_4289_16) begin
      _T_5840 <= _T_4492_16;
    end
    if (_T_4289_16) begin
      _T_5842 <= _T_4492_16;
    end
    if (_T_4289_17) begin
      _T_5844 <= _T_4492_17;
    end
    if (_T_4289_17) begin
      _T_5846 <= _T_4492_17;
    end
    if (_T_4289_18) begin
      _T_5848 <= _T_4492_18;
    end
    if (_T_4289_18) begin
      _T_5850 <= _T_4492_18;
    end
    if (_T_4289_19) begin
      _T_5852 <= _T_4492_19;
    end
    if (_T_4289_19) begin
      _T_5854 <= _T_4492_19;
    end
    if (_T_4289_20) begin
      _T_5856 <= _T_4492_20;
    end
    if (_T_4289_20) begin
      _T_5858 <= _T_4492_20;
    end
    if (_T_4289_21) begin
      _T_5860 <= _T_4492_21;
    end
    if (_T_4289_21) begin
      _T_5862 <= _T_4492_21;
    end
    if (_T_4289_22) begin
      _T_5864 <= _T_4492_22;
    end
    if (_T_4289_22) begin
      _T_5866 <= _T_4492_22;
    end
    if (_T_4289_23) begin
      _T_5868 <= _T_4492_23;
    end
    if (_T_4289_23) begin
      _T_5870 <= _T_4492_23;
    end
    if (_T_4289_24) begin
      _T_5872 <= _T_4492_24;
    end
    if (_T_4289_24) begin
      _T_5874 <= _T_4492_24;
    end
    if (_T_4289_25) begin
      _T_5876 <= _T_4492_25;
    end
    if (_T_4289_25) begin
      _T_5878 <= _T_4492_25;
    end
    if (_T_4289_26) begin
      _T_5880 <= _T_4492_26;
    end
    if (_T_4289_26) begin
      _T_5882 <= _T_4492_26;
    end
    if (_T_4289_27) begin
      _T_5884 <= _T_4492_27;
    end
    if (_T_4289_27) begin
      _T_5886 <= _T_4492_27;
    end
    if (_T_4289_28) begin
      _T_5888 <= _T_4492_28;
    end
    if (_T_4289_28) begin
      _T_5890 <= _T_4492_28;
    end
    if (_T_4289_29) begin
      _T_5892 <= _T_4492_29;
    end
    if (_T_4289_29) begin
      _T_5894 <= _T_4492_29;
    end
    if (_T_4289_30) begin
      _T_5896 <= _T_4492_30;
    end
    if (_T_4289_30) begin
      _T_5898 <= _T_4492_30;
    end
    if (_T_4289_31) begin
      _T_5900 <= _T_4492_31;
    end
    if (_T_4289_31) begin
      _T_5902 <= _T_4492_31;
    end
    if (_T_4289_32) begin
      _T_5904 <= _T_4492_32;
    end
    if (_T_4289_32) begin
      _T_5906 <= _T_4492_32;
    end
    if (_T_4289_33) begin
      _T_5908 <= _T_4492_33;
    end
    if (_T_4289_33) begin
      _T_5910 <= _T_4492_33;
    end
    if (_T_4289_34) begin
      _T_5912 <= _T_4492_34;
    end
    if (_T_4289_34) begin
      _T_5914 <= _T_4492_34;
    end
    if (_T_4289_35) begin
      _T_5916 <= _T_4492_35;
    end
    if (_T_4289_35) begin
      _T_5918 <= _T_4492_35;
    end
    if (_T_4289_36) begin
      _T_5920 <= _T_4492_36;
    end
    if (_T_4289_36) begin
      _T_5922 <= _T_4492_36;
    end
    if (_T_4289_37) begin
      _T_5924 <= _T_4492_37;
    end
    if (_T_4289_37) begin
      _T_5926 <= _T_4492_37;
    end
    if (_T_4289_38) begin
      _T_5928 <= _T_4492_38;
    end
    if (_T_4289_38) begin
      _T_5930 <= _T_4492_38;
    end
    if (_T_4289_39) begin
      _T_5932 <= _T_4492_39;
    end
    if (_T_4289_39) begin
      _T_5934 <= _T_4492_39;
    end
    if (_T_4289_40) begin
      _T_5936 <= _T_4492_40;
    end
    if (_T_4289_40) begin
      _T_5938 <= _T_4492_40;
    end
    if (_T_4289_41) begin
      _T_5940 <= _T_4492_41;
    end
    if (_T_4289_41) begin
      _T_5942 <= _T_4492_41;
    end
    if (_T_4289_42) begin
      _T_5944 <= _T_4492_42;
    end
    if (_T_4289_42) begin
      _T_5946 <= _T_4492_42;
    end
    if (_T_4289_43) begin
      _T_5948 <= _T_4492_43;
    end
    if (_T_4289_43) begin
      _T_5950 <= _T_4492_43;
    end
    if (_T_4289_44) begin
      _T_5952 <= _T_4492_44;
    end
    if (_T_4289_44) begin
      _T_5954 <= _T_4492_44;
    end
    if (_T_4289_45) begin
      _T_5956 <= _T_4492_45;
    end
    if (_T_4289_45) begin
      _T_5958 <= _T_4492_45;
    end
    if (_T_4289_46) begin
      _T_5960 <= _T_4492_46;
    end
    if (_T_4289_46) begin
      _T_5962 <= _T_4492_46;
    end
    if (_T_4289_47) begin
      _T_5964 <= _T_4492_47;
    end
    if (_T_4289_47) begin
      _T_5966 <= _T_4492_47;
    end
    if (_T_4289_48) begin
      _T_5968 <= _T_4492_48;
    end
    if (_T_4289_48) begin
      _T_5970 <= _T_4492_48;
    end
    if (_T_4289_49) begin
      _T_5972 <= _T_4492_49;
    end
    if (_T_4289_49) begin
      _T_5974 <= _T_4492_49;
    end
    if (_T_4289_50) begin
      _T_5976 <= _T_4492_50;
    end
    if (_T_4289_50) begin
      _T_5978 <= _T_4492_50;
    end
    if (_T_4289_51) begin
      _T_5980 <= _T_4492_51;
    end
    if (_T_4289_51) begin
      _T_5982 <= _T_4492_51;
    end
    if (_T_4289_52) begin
      _T_5984 <= _T_4492_52;
    end
    if (_T_4289_52) begin
      _T_5986 <= _T_4492_52;
    end
    if (_T_4289_53) begin
      _T_5988 <= _T_4492_53;
    end
    if (_T_4289_53) begin
      _T_5990 <= _T_4492_53;
    end
    if (_T_4289_54) begin
      _T_5992 <= _T_4492_54;
    end
    if (_T_4289_54) begin
      _T_5994 <= _T_4492_54;
    end
    if (_T_4289_55) begin
      _T_5996 <= _T_4492_55;
    end
    if (_T_4289_55) begin
      _T_5998 <= _T_4492_55;
    end
    if (_T_4289_56) begin
      _T_6000 <= _T_4492_56;
    end
    if (_T_4289_56) begin
      _T_6002 <= _T_4492_56;
    end
    if (_T_4289_57) begin
      _T_6004 <= _T_4492_57;
    end
    if (_T_4289_57) begin
      _T_6006 <= _T_4492_57;
    end
    if (_T_4289_58) begin
      _T_6008 <= _T_4492_58;
    end
    if (_T_4289_58) begin
      _T_6010 <= _T_4492_58;
    end
    if (_T_4289_59) begin
      _T_6012 <= _T_4492_59;
    end
    if (_T_4289_59) begin
      _T_6014 <= _T_4492_59;
    end
    if (_T_4289_60) begin
      _T_6016 <= _T_4492_60;
    end
    if (_T_4289_60) begin
      _T_6018 <= _T_4492_60;
    end
    if (_T_4289_61) begin
      _T_6020 <= _T_4492_61;
    end
    if (_T_4289_61) begin
      _T_6022 <= _T_4492_61;
    end
    if (_T_4289_62) begin
      _T_6024 <= _T_4492_62;
    end
    if (_T_4289_62) begin
      _T_6026 <= _T_4492_62;
    end
    if (_T_4289_63) begin
      _T_6028 <= _T_4492_63;
    end
    if (_T_4289_63) begin
      _T_6030 <= _T_4492_63;
    end
  end
  always @(posedge io_nvdla_core_ng_clk) begin
    if (reset) begin
      _T_1076 <= 15'h0;
    end else begin
      if (_T_1148) begin
        if (io_sc2cdma_dat_pending_req) begin
          _T_1076 <= 15'h0;
        end else begin
          if (_T_1119) begin
            _T_1076 <= _T_1112;
          end else begin
            _T_1076 <= _T_1103;
          end
        end
      end
    end
  end
endmodule
module NV_NVDLA_slcg( // @[:@23604.2]
  input   io_nvdla_clock_nvdla_core_clk, // @[:@23607.4]
  output  io_nvdla_core_gated_clk // @[:@23607.4]
);
  assign io_nvdla_core_gated_clk = io_nvdla_clock_nvdla_core_clk; // @[slcg.scala 23:31:@23609.4]
endmodule
module NV_soDLA_csc( // @[:@23625.2]
  input          clock, // @[:@23626.4]
  input          reset, // @[:@23627.4]
  input          io_nvdla_clock_nvdla_core_clk, // @[:@23628.4]
  input          io_nvdla_clock_dla_clk_ovr_on_sync, // @[:@23628.4]
  input          io_nvdla_clock_global_clk_ovr_on_sync, // @[:@23628.4]
  input          io_nvdla_clock_tmc2slcg_disable_clock_gating, // @[:@23628.4]
  input          io_nvdla_core_rstn, // @[:@23628.4]
  output         io_sc2cdma_dat_pending_req, // @[:@23628.4]
  output         io_sc2cdma_wt_pending_req, // @[:@23628.4]
  input          io_cdma2sc_dat_pending_ack, // @[:@23628.4]
  input          io_cdma2sc_wt_pending_ack, // @[:@23628.4]
  input          io_cdma2sc_dat_updt_valid, // @[:@23628.4]
  input  [14:0]  io_cdma2sc_dat_updt_bits_entries, // @[:@23628.4]
  input  [13:0]  io_cdma2sc_dat_updt_bits_slices, // @[:@23628.4]
  output         io_sc2cdma_dat_updt_valid, // @[:@23628.4]
  output [14:0]  io_sc2cdma_dat_updt_bits_entries, // @[:@23628.4]
  output [13:0]  io_sc2cdma_dat_updt_bits_slices, // @[:@23628.4]
  input          io_cdma2sc_wt_updt_valid, // @[:@23628.4]
  input  [14:0]  io_cdma2sc_wt_updt_bits_entries, // @[:@23628.4]
  input  [13:0]  io_cdma2sc_wt_updt_bits_kernels, // @[:@23628.4]
  output         io_sc2cdma_wt_updt_valid, // @[:@23628.4]
  output [14:0]  io_sc2cdma_wt_updt_bits_entries, // @[:@23628.4]
  output [13:0]  io_sc2cdma_wt_updt_bits_kernels, // @[:@23628.4]
  output [8:0]   io_sc2cdma_wmb_entries, // @[:@23628.4]
  input  [8:0]   io_cdma2sc_wmb_entries, // @[:@23628.4]
  input          io_accu2sc_credit_size_valid, // @[:@23628.4]
  input  [2:0]   io_accu2sc_credit_size_bits, // @[:@23628.4]
  output         io_csb2csc_req_ready, // @[:@23628.4]
  input          io_csb2csc_req_valid, // @[:@23628.4]
  input  [62:0]  io_csb2csc_req_bits, // @[:@23628.4]
  output         io_csb2csc_resp_valid, // @[:@23628.4]
  output [33:0]  io_csb2csc_resp_bits, // @[:@23628.4]
  output         io_sc2buf_dat_rd_addr_valid, // @[:@23628.4]
  output [12:0]  io_sc2buf_dat_rd_addr_bits, // @[:@23628.4]
  input          io_sc2buf_dat_rd_data_valid, // @[:@23628.4]
  input  [511:0] io_sc2buf_dat_rd_data_bits, // @[:@23628.4]
  output         io_sc2buf_wt_rd_addr_valid, // @[:@23628.4]
  output [12:0]  io_sc2buf_wt_rd_addr_bits, // @[:@23628.4]
  input          io_sc2buf_wt_rd_data_valid, // @[:@23628.4]
  input  [511:0] io_sc2buf_wt_rd_data_bits, // @[:@23628.4]
  output         io_sc2mac_dat_a_valid, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_0, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_1, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_2, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_3, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_4, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_5, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_6, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_7, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_8, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_9, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_10, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_11, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_12, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_13, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_14, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_15, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_16, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_17, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_18, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_19, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_20, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_21, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_22, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_23, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_24, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_25, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_26, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_27, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_28, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_29, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_30, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_31, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_32, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_33, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_34, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_35, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_36, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_37, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_38, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_39, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_40, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_41, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_42, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_43, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_44, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_45, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_46, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_47, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_48, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_49, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_50, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_51, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_52, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_53, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_54, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_55, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_56, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_57, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_58, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_59, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_60, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_61, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_62, // @[:@23628.4]
  output         io_sc2mac_dat_a_bits_mask_63, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_0, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_1, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_2, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_3, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_4, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_5, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_6, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_7, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_8, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_9, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_10, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_11, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_12, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_13, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_14, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_15, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_16, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_17, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_18, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_19, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_20, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_21, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_22, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_23, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_24, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_25, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_26, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_27, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_28, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_29, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_30, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_31, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_32, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_33, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_34, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_35, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_36, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_37, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_38, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_39, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_40, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_41, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_42, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_43, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_44, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_45, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_46, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_47, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_48, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_49, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_50, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_51, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_52, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_53, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_54, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_55, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_56, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_57, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_58, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_59, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_60, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_61, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_62, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_63, // @[:@23628.4]
  output [8:0]   io_sc2mac_dat_a_bits_pd, // @[:@23628.4]
  output         io_sc2mac_dat_b_valid, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_0, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_1, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_2, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_3, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_4, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_5, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_6, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_7, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_8, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_9, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_10, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_11, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_12, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_13, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_14, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_15, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_16, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_17, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_18, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_19, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_20, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_21, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_22, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_23, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_24, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_25, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_26, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_27, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_28, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_29, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_30, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_31, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_32, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_33, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_34, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_35, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_36, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_37, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_38, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_39, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_40, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_41, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_42, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_43, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_44, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_45, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_46, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_47, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_48, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_49, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_50, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_51, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_52, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_53, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_54, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_55, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_56, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_57, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_58, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_59, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_60, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_61, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_62, // @[:@23628.4]
  output         io_sc2mac_dat_b_bits_mask_63, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_0, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_1, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_2, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_3, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_4, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_5, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_6, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_7, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_8, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_9, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_10, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_11, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_12, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_13, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_14, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_15, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_16, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_17, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_18, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_19, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_20, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_21, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_22, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_23, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_24, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_25, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_26, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_27, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_28, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_29, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_30, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_31, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_32, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_33, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_34, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_35, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_36, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_37, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_38, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_39, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_40, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_41, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_42, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_43, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_44, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_45, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_46, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_47, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_48, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_49, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_50, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_51, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_52, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_53, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_54, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_55, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_56, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_57, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_58, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_59, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_60, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_61, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_62, // @[:@23628.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_63, // @[:@23628.4]
  output [8:0]   io_sc2mac_dat_b_bits_pd, // @[:@23628.4]
  output         io_sc2mac_wt_a_valid, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_sel_0, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_sel_1, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_sel_2, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_sel_3, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_sel_4, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_sel_5, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_sel_6, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_sel_7, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_sel_8, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_sel_9, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_sel_10, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_sel_11, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_sel_12, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_sel_13, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_sel_14, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_sel_15, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_0, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_1, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_2, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_3, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_4, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_5, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_6, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_7, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_8, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_9, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_10, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_11, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_12, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_13, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_14, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_15, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_16, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_17, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_18, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_19, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_20, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_21, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_22, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_23, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_24, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_25, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_26, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_27, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_28, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_29, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_30, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_31, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_32, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_33, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_34, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_35, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_36, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_37, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_38, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_39, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_40, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_41, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_42, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_43, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_44, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_45, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_46, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_47, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_48, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_49, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_50, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_51, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_52, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_53, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_54, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_55, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_56, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_57, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_58, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_59, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_60, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_61, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_62, // @[:@23628.4]
  output         io_sc2mac_wt_a_bits_mask_63, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_0, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_1, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_2, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_3, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_4, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_5, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_6, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_7, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_8, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_9, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_10, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_11, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_12, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_13, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_14, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_15, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_16, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_17, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_18, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_19, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_20, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_21, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_22, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_23, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_24, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_25, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_26, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_27, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_28, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_29, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_30, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_31, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_32, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_33, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_34, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_35, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_36, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_37, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_38, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_39, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_40, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_41, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_42, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_43, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_44, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_45, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_46, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_47, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_48, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_49, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_50, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_51, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_52, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_53, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_54, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_55, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_56, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_57, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_58, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_59, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_60, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_61, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_62, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_63, // @[:@23628.4]
  output         io_sc2mac_wt_b_valid, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_sel_0, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_sel_1, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_sel_2, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_sel_3, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_sel_4, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_sel_5, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_sel_6, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_sel_7, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_sel_8, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_sel_9, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_sel_10, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_sel_11, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_sel_12, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_sel_13, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_sel_14, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_sel_15, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_0, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_1, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_2, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_3, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_4, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_5, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_6, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_7, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_8, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_9, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_10, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_11, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_12, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_13, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_14, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_15, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_16, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_17, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_18, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_19, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_20, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_21, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_22, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_23, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_24, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_25, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_26, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_27, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_28, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_29, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_30, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_31, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_32, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_33, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_34, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_35, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_36, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_37, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_38, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_39, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_40, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_41, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_42, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_43, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_44, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_45, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_46, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_47, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_48, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_49, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_50, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_51, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_52, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_53, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_54, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_55, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_56, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_57, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_58, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_59, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_60, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_61, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_62, // @[:@23628.4]
  output         io_sc2mac_wt_b_bits_mask_63, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_0, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_1, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_2, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_3, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_4, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_5, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_6, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_7, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_8, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_9, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_10, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_11, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_12, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_13, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_14, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_15, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_16, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_17, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_18, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_19, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_20, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_21, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_22, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_23, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_24, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_25, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_26, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_27, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_28, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_29, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_30, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_31, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_32, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_33, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_34, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_35, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_36, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_37, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_38, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_39, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_40, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_41, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_42, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_43, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_44, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_45, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_46, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_47, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_48, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_49, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_50, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_51, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_52, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_53, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_54, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_55, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_56, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_57, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_58, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_59, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_60, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_61, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_62, // @[:@23628.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_63, // @[:@23628.4]
  input  [31:0]  io_pwrbus_ram_pd // @[:@23628.4]
);
  wire  NV_NVDLA_CSC_regfile_reset; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire  NV_NVDLA_CSC_regfile_io_nvdla_core_clk; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire  NV_NVDLA_CSC_regfile_io_csb2csc_req_valid; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [62:0] NV_NVDLA_CSC_regfile_io_csb2csc_req_bits; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire  NV_NVDLA_CSC_regfile_io_csb2csc_resp_valid; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [33:0] NV_NVDLA_CSC_regfile_io_csb2csc_resp_bits; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire  NV_NVDLA_CSC_regfile_io_reg2dp_op_en; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [20:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_atomics; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [4:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_data_bank; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [4:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_bank; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [2:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_conv_x_stride_ext; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [2:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_conv_y_stride_ext; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire  NV_NVDLA_CSC_regfile_io_reg2dp_field_datain_format; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [12:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_datain_height_ext; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [12:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_datain_width_ext; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [12:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_datain_channel_ext; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [12:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_dataout_height; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [12:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_dataout_width; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [4:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_x_dilation_ext; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [4:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_y_dilation_ext; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [13:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_entries; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire  NV_NVDLA_CSC_regfile_io_reg2dp_field_conv_mode; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire  NV_NVDLA_CSC_regfile_io_reg2dp_field_data_reuse; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire  NV_NVDLA_CSC_regfile_io_reg2dp_field_skip_data_rls; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire  NV_NVDLA_CSC_regfile_io_reg2dp_field_skip_weight_rls; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire  NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_reuse; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [1:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_y_extension; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [11:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_rls_slices; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [31:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_bytes; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire  NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_format; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [4:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_height_ext; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [4:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_width_ext; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [12:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_channel_ext; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [12:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_kernel; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [27:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_wmb_bytes; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [4:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_pad_left; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [4:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_pad_top; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire [15:0] NV_NVDLA_CSC_regfile_io_reg2dp_field_pad_value; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire  NV_NVDLA_CSC_regfile_io_dp2reg_done; // @[NV_NVDLA_csc.scala 76:27:@23632.4]
  wire  NV_NVDLA_CSC_sg_reset; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_nvdla_core_clk; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_nvdla_core_ng_clk; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_cdma2sc_dat_updt_valid; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire [13:0] NV_NVDLA_CSC_sg_io_cdma2sc_dat_updt_bits_slices; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_sc2cdma_dat_pending_req; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_cdma2sc_dat_pending_ack; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_cdma2sc_wt_updt_valid; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire [13:0] NV_NVDLA_CSC_sg_io_cdma2sc_wt_updt_bits_kernels; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_sc2cdma_wt_pending_req; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_cdma2sc_wt_pending_ack; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire [1:0] NV_NVDLA_CSC_sg_io_sc_state; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_sg2dl_pd_valid; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_sg2dl_reuse_rls; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_sg2wl_pd_valid; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire [17:0] NV_NVDLA_CSC_sg_io_sg2wl_pd_bits; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_sg2wl_reuse_rls; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_accu2sc_credit_size_valid; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire [2:0] NV_NVDLA_CSC_sg_io_accu2sc_credit_size_bits; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_reg2dp_op_en; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_reg2dp_conv_mode; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_reg2dp_data_reuse; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_reg2dp_skip_data_rls; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_reg2dp_weight_reuse; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_reg2dp_skip_weight_rls; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_reg2dp_datain_format; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire [12:0] NV_NVDLA_CSC_sg_io_reg2dp_datain_height_ext; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire [1:0] NV_NVDLA_CSC_sg_io_reg2dp_y_extension; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire [4:0] NV_NVDLA_CSC_sg_io_reg2dp_weight_width_ext; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire [4:0] NV_NVDLA_CSC_sg_io_reg2dp_weight_height_ext; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire [12:0] NV_NVDLA_CSC_sg_io_reg2dp_weight_channel_ext; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire [12:0] NV_NVDLA_CSC_sg_io_reg2dp_weight_kernel; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire [12:0] NV_NVDLA_CSC_sg_io_reg2dp_dataout_width; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire [12:0] NV_NVDLA_CSC_sg_io_reg2dp_dataout_height; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire [4:0] NV_NVDLA_CSC_sg_io_reg2dp_data_bank; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire [4:0] NV_NVDLA_CSC_sg_io_reg2dp_weight_bank; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire [20:0] NV_NVDLA_CSC_sg_io_reg2dp_atomics; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire [11:0] NV_NVDLA_CSC_sg_io_reg2dp_rls_slices; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_sg_io_dp2reg_done; // @[NV_NVDLA_csc.scala 77:22:@23635.4]
  wire  NV_NVDLA_CSC_wl_reset; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_nvdla_core_clk; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_nvdla_core_ng_clk; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sg2wl_pd_valid; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [17:0] NV_NVDLA_CSC_wl_io_sg2wl_pd_bits; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sg2wl_reuse_rls; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [1:0] NV_NVDLA_CSC_wl_io_sc_state; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2cdma_wt_pending_req; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2cdma_wt_updt_valid; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [14:0] NV_NVDLA_CSC_wl_io_sc2cdma_wt_updt_bits_entries; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [8:0] NV_NVDLA_CSC_wl_io_sc2cdma_wmb_entries; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2buf_wt_rd_addr_valid; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [12:0] NV_NVDLA_CSC_wl_io_sc2buf_wt_rd_addr_bits; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2buf_wt_rd_data_valid; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [511:0] NV_NVDLA_CSC_wl_io_sc2buf_wt_rd_data_bits; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_valid; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_0; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_1; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_2; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_3; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_4; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_5; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_6; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_7; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_8; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_9; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_10; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_11; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_12; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_13; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_14; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_15; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_0; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_1; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_2; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_3; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_4; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_5; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_6; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_7; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_8; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_9; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_10; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_11; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_12; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_13; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_14; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_15; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_16; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_17; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_18; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_19; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_20; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_21; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_22; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_23; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_24; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_25; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_26; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_27; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_28; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_29; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_30; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_31; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_32; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_33; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_34; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_35; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_36; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_37; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_38; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_39; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_40; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_41; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_42; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_43; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_44; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_45; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_46; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_47; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_48; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_49; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_50; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_51; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_52; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_53; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_54; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_55; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_56; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_57; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_58; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_59; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_60; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_61; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_62; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_63; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_0; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_1; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_2; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_3; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_4; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_5; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_6; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_7; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_8; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_9; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_10; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_11; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_12; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_13; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_14; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_15; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_16; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_17; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_18; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_19; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_20; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_21; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_22; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_23; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_24; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_25; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_26; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_27; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_28; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_29; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_30; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_31; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_32; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_33; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_34; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_35; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_36; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_37; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_38; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_39; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_40; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_41; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_42; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_43; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_44; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_45; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_46; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_47; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_48; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_49; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_50; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_51; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_52; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_53; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_54; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_55; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_56; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_57; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_58; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_59; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_60; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_61; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_62; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_63; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_valid; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_0; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_1; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_2; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_3; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_4; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_5; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_6; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_7; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_8; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_9; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_10; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_11; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_12; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_13; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_14; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_15; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_0; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_1; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_2; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_3; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_4; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_5; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_6; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_7; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_8; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_9; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_10; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_11; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_12; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_13; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_14; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_15; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_16; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_17; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_18; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_19; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_20; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_21; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_22; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_23; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_24; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_25; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_26; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_27; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_28; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_29; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_30; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_31; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_32; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_33; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_34; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_35; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_36; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_37; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_38; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_39; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_40; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_41; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_42; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_43; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_44; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_45; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_46; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_47; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_48; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_49; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_50; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_51; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_52; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_53; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_54; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_55; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_56; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_57; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_58; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_59; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_60; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_61; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_62; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_63; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_0; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_1; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_2; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_3; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_4; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_5; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_6; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_7; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_8; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_9; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_10; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_11; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_12; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_13; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_14; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_15; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_16; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_17; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_18; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_19; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_20; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_21; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_22; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_23; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_24; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_25; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_26; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_27; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_28; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_29; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_30; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_31; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_32; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_33; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_34; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_35; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_36; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_37; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_38; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_39; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_40; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_41; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_42; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_43; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_44; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_45; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_46; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_47; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_48; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_49; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_50; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_51; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_52; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_53; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_54; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_55; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_56; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_57; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_58; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_59; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_60; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_61; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_62; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [7:0] NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_63; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_reg2dp_op_en; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [1:0] NV_NVDLA_CSC_wl_io_reg2dp_y_extension; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_reg2dp_skip_weight_rls; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_wl_io_reg2dp_weight_format; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [31:0] NV_NVDLA_CSC_wl_io_reg2dp_weight_bytes; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [27:0] NV_NVDLA_CSC_wl_io_reg2dp_wmb_bytes; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [4:0] NV_NVDLA_CSC_wl_io_reg2dp_data_bank; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire [4:0] NV_NVDLA_CSC_wl_io_reg2dp_weight_bank; // @[NV_NVDLA_csc.scala 129:22:@23683.4]
  wire  NV_NVDLA_CSC_dl_reset; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_nvdla_core_clk; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_nvdla_core_ng_clk; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [1:0] NV_NVDLA_CSC_dl_io_sc_state; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sg2dl_pd_valid; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sg2dl_reuse_rls; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2cdma_dat_pending_req; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2cdma_dat_updt_valid; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [14:0] NV_NVDLA_CSC_dl_io_sc2cdma_dat_updt_bits_entries; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [13:0] NV_NVDLA_CSC_dl_io_sc2cdma_dat_updt_bits_slices; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2buf_dat_rd_addr_valid; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [12:0] NV_NVDLA_CSC_dl_io_sc2buf_dat_rd_addr_bits; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2buf_dat_rd_data_valid; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [511:0] NV_NVDLA_CSC_dl_io_sc2buf_dat_rd_data_bits; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_valid; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_0; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_1; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_2; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_3; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_4; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_5; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_6; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_7; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_8; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_9; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_10; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_11; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_12; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_13; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_14; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_15; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_16; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_17; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_18; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_19; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_20; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_21; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_22; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_23; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_24; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_25; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_26; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_27; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_28; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_29; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_30; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_31; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_32; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_33; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_34; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_35; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_36; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_37; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_38; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_39; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_40; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_41; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_42; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_43; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_44; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_45; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_46; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_47; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_48; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_49; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_50; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_51; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_52; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_53; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_54; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_55; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_56; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_57; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_58; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_59; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_60; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_61; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_62; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_63; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_0; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_1; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_2; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_3; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_4; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_5; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_6; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_7; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_8; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_9; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_10; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_11; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_12; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_13; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_14; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_15; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_16; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_17; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_18; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_19; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_20; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_21; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_22; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_23; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_24; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_25; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_26; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_27; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_28; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_29; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_30; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_31; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_32; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_33; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_34; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_35; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_36; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_37; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_38; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_39; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_40; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_41; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_42; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_43; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_44; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_45; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_46; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_47; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_48; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_49; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_50; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_51; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_52; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_53; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_54; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_55; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_56; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_57; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_58; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_59; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_60; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_61; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_62; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_63; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [8:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_pd; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_valid; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_0; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_1; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_2; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_3; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_4; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_5; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_6; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_7; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_8; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_9; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_10; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_11; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_12; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_13; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_14; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_15; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_16; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_17; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_18; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_19; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_20; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_21; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_22; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_23; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_24; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_25; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_26; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_27; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_28; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_29; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_30; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_31; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_32; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_33; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_34; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_35; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_36; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_37; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_38; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_39; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_40; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_41; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_42; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_43; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_44; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_45; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_46; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_47; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_48; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_49; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_50; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_51; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_52; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_53; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_54; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_55; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_56; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_57; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_58; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_59; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_60; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_61; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_62; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_63; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_0; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_1; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_2; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_3; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_4; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_5; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_6; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_7; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_8; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_9; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_10; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_11; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_12; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_13; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_14; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_15; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_16; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_17; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_18; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_19; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_20; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_21; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_22; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_23; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_24; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_25; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_26; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_27; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_28; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_29; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_30; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_31; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_32; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_33; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_34; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_35; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_36; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_37; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_38; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_39; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_40; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_41; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_42; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_43; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_44; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_45; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_46; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_47; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_48; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_49; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_50; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_51; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_52; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_53; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_54; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_55; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_56; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_57; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_58; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_59; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_60; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_61; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_62; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [7:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_63; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [8:0] NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_pd; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_reg2dp_op_en; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_reg2dp_conv_mode; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_reg2dp_datain_format; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_CSC_dl_io_reg2dp_skip_data_rls; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [12:0] NV_NVDLA_CSC_dl_io_reg2dp_datain_channel_ext; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [12:0] NV_NVDLA_CSC_dl_io_reg2dp_datain_height_ext; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [12:0] NV_NVDLA_CSC_dl_io_reg2dp_datain_width_ext; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [1:0] NV_NVDLA_CSC_dl_io_reg2dp_y_extension; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [12:0] NV_NVDLA_CSC_dl_io_reg2dp_weight_channel_ext; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [13:0] NV_NVDLA_CSC_dl_io_reg2dp_entries; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [12:0] NV_NVDLA_CSC_dl_io_reg2dp_dataout_width; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [11:0] NV_NVDLA_CSC_dl_io_reg2dp_rls_slices; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [2:0] NV_NVDLA_CSC_dl_io_reg2dp_conv_x_stride_ext; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [2:0] NV_NVDLA_CSC_dl_io_reg2dp_conv_y_stride_ext; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [4:0] NV_NVDLA_CSC_dl_io_reg2dp_x_dilation_ext; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [4:0] NV_NVDLA_CSC_dl_io_reg2dp_y_dilation_ext; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [4:0] NV_NVDLA_CSC_dl_io_reg2dp_pad_left; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [4:0] NV_NVDLA_CSC_dl_io_reg2dp_pad_top; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [15:0] NV_NVDLA_CSC_dl_io_reg2dp_pad_value; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire [4:0] NV_NVDLA_CSC_dl_io_reg2dp_data_bank; // @[NV_NVDLA_csc.scala 161:22:@24006.4]
  wire  NV_NVDLA_slcg_io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_csc.scala 205:41:@24309.4]
  wire  NV_NVDLA_slcg_io_nvdla_core_gated_clk; // @[NV_NVDLA_csc.scala 205:41:@24309.4]
  wire  NV_NVDLA_slcg_1_io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_csc.scala 205:41:@24312.4]
  wire  NV_NVDLA_slcg_1_io_nvdla_core_gated_clk; // @[NV_NVDLA_csc.scala 205:41:@24312.4]
  wire  NV_NVDLA_slcg_2_io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_csc.scala 205:41:@24315.4]
  wire  NV_NVDLA_slcg_2_io_nvdla_core_gated_clk; // @[NV_NVDLA_csc.scala 205:41:@24315.4]
  NV_NVDLA_CSC_regfile NV_NVDLA_CSC_regfile ( // @[NV_NVDLA_csc.scala 76:27:@23632.4]
    .reset(NV_NVDLA_CSC_regfile_reset),
    .io_nvdla_core_clk(NV_NVDLA_CSC_regfile_io_nvdla_core_clk),
    .io_csb2csc_req_valid(NV_NVDLA_CSC_regfile_io_csb2csc_req_valid),
    .io_csb2csc_req_bits(NV_NVDLA_CSC_regfile_io_csb2csc_req_bits),
    .io_csb2csc_resp_valid(NV_NVDLA_CSC_regfile_io_csb2csc_resp_valid),
    .io_csb2csc_resp_bits(NV_NVDLA_CSC_regfile_io_csb2csc_resp_bits),
    .io_reg2dp_op_en(NV_NVDLA_CSC_regfile_io_reg2dp_op_en),
    .io_reg2dp_field_atomics(NV_NVDLA_CSC_regfile_io_reg2dp_field_atomics),
    .io_reg2dp_field_data_bank(NV_NVDLA_CSC_regfile_io_reg2dp_field_data_bank),
    .io_reg2dp_field_weight_bank(NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_bank),
    .io_reg2dp_field_conv_x_stride_ext(NV_NVDLA_CSC_regfile_io_reg2dp_field_conv_x_stride_ext),
    .io_reg2dp_field_conv_y_stride_ext(NV_NVDLA_CSC_regfile_io_reg2dp_field_conv_y_stride_ext),
    .io_reg2dp_field_datain_format(NV_NVDLA_CSC_regfile_io_reg2dp_field_datain_format),
    .io_reg2dp_field_datain_height_ext(NV_NVDLA_CSC_regfile_io_reg2dp_field_datain_height_ext),
    .io_reg2dp_field_datain_width_ext(NV_NVDLA_CSC_regfile_io_reg2dp_field_datain_width_ext),
    .io_reg2dp_field_datain_channel_ext(NV_NVDLA_CSC_regfile_io_reg2dp_field_datain_channel_ext),
    .io_reg2dp_field_dataout_height(NV_NVDLA_CSC_regfile_io_reg2dp_field_dataout_height),
    .io_reg2dp_field_dataout_width(NV_NVDLA_CSC_regfile_io_reg2dp_field_dataout_width),
    .io_reg2dp_field_x_dilation_ext(NV_NVDLA_CSC_regfile_io_reg2dp_field_x_dilation_ext),
    .io_reg2dp_field_y_dilation_ext(NV_NVDLA_CSC_regfile_io_reg2dp_field_y_dilation_ext),
    .io_reg2dp_field_entries(NV_NVDLA_CSC_regfile_io_reg2dp_field_entries),
    .io_reg2dp_field_conv_mode(NV_NVDLA_CSC_regfile_io_reg2dp_field_conv_mode),
    .io_reg2dp_field_data_reuse(NV_NVDLA_CSC_regfile_io_reg2dp_field_data_reuse),
    .io_reg2dp_field_skip_data_rls(NV_NVDLA_CSC_regfile_io_reg2dp_field_skip_data_rls),
    .io_reg2dp_field_skip_weight_rls(NV_NVDLA_CSC_regfile_io_reg2dp_field_skip_weight_rls),
    .io_reg2dp_field_weight_reuse(NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_reuse),
    .io_reg2dp_field_y_extension(NV_NVDLA_CSC_regfile_io_reg2dp_field_y_extension),
    .io_reg2dp_field_rls_slices(NV_NVDLA_CSC_regfile_io_reg2dp_field_rls_slices),
    .io_reg2dp_field_weight_bytes(NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_bytes),
    .io_reg2dp_field_weight_format(NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_format),
    .io_reg2dp_field_weight_height_ext(NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_height_ext),
    .io_reg2dp_field_weight_width_ext(NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_width_ext),
    .io_reg2dp_field_weight_channel_ext(NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_channel_ext),
    .io_reg2dp_field_weight_kernel(NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_kernel),
    .io_reg2dp_field_wmb_bytes(NV_NVDLA_CSC_regfile_io_reg2dp_field_wmb_bytes),
    .io_reg2dp_field_pad_left(NV_NVDLA_CSC_regfile_io_reg2dp_field_pad_left),
    .io_reg2dp_field_pad_top(NV_NVDLA_CSC_regfile_io_reg2dp_field_pad_top),
    .io_reg2dp_field_pad_value(NV_NVDLA_CSC_regfile_io_reg2dp_field_pad_value),
    .io_dp2reg_done(NV_NVDLA_CSC_regfile_io_dp2reg_done)
  );
  NV_NVDLA_CSC_sg NV_NVDLA_CSC_sg ( // @[NV_NVDLA_csc.scala 77:22:@23635.4]
    .reset(NV_NVDLA_CSC_sg_reset),
    .io_nvdla_core_clk(NV_NVDLA_CSC_sg_io_nvdla_core_clk),
    .io_nvdla_core_ng_clk(NV_NVDLA_CSC_sg_io_nvdla_core_ng_clk),
    .io_cdma2sc_dat_updt_valid(NV_NVDLA_CSC_sg_io_cdma2sc_dat_updt_valid),
    .io_cdma2sc_dat_updt_bits_slices(NV_NVDLA_CSC_sg_io_cdma2sc_dat_updt_bits_slices),
    .io_sc2cdma_dat_pending_req(NV_NVDLA_CSC_sg_io_sc2cdma_dat_pending_req),
    .io_cdma2sc_dat_pending_ack(NV_NVDLA_CSC_sg_io_cdma2sc_dat_pending_ack),
    .io_cdma2sc_wt_updt_valid(NV_NVDLA_CSC_sg_io_cdma2sc_wt_updt_valid),
    .io_cdma2sc_wt_updt_bits_kernels(NV_NVDLA_CSC_sg_io_cdma2sc_wt_updt_bits_kernels),
    .io_sc2cdma_wt_pending_req(NV_NVDLA_CSC_sg_io_sc2cdma_wt_pending_req),
    .io_cdma2sc_wt_pending_ack(NV_NVDLA_CSC_sg_io_cdma2sc_wt_pending_ack),
    .io_sc_state(NV_NVDLA_CSC_sg_io_sc_state),
    .io_sg2dl_pd_valid(NV_NVDLA_CSC_sg_io_sg2dl_pd_valid),
    .io_sg2dl_reuse_rls(NV_NVDLA_CSC_sg_io_sg2dl_reuse_rls),
    .io_sg2wl_pd_valid(NV_NVDLA_CSC_sg_io_sg2wl_pd_valid),
    .io_sg2wl_pd_bits(NV_NVDLA_CSC_sg_io_sg2wl_pd_bits),
    .io_sg2wl_reuse_rls(NV_NVDLA_CSC_sg_io_sg2wl_reuse_rls),
    .io_accu2sc_credit_size_valid(NV_NVDLA_CSC_sg_io_accu2sc_credit_size_valid),
    .io_accu2sc_credit_size_bits(NV_NVDLA_CSC_sg_io_accu2sc_credit_size_bits),
    .io_reg2dp_op_en(NV_NVDLA_CSC_sg_io_reg2dp_op_en),
    .io_reg2dp_conv_mode(NV_NVDLA_CSC_sg_io_reg2dp_conv_mode),
    .io_reg2dp_data_reuse(NV_NVDLA_CSC_sg_io_reg2dp_data_reuse),
    .io_reg2dp_skip_data_rls(NV_NVDLA_CSC_sg_io_reg2dp_skip_data_rls),
    .io_reg2dp_weight_reuse(NV_NVDLA_CSC_sg_io_reg2dp_weight_reuse),
    .io_reg2dp_skip_weight_rls(NV_NVDLA_CSC_sg_io_reg2dp_skip_weight_rls),
    .io_reg2dp_datain_format(NV_NVDLA_CSC_sg_io_reg2dp_datain_format),
    .io_reg2dp_datain_height_ext(NV_NVDLA_CSC_sg_io_reg2dp_datain_height_ext),
    .io_reg2dp_y_extension(NV_NVDLA_CSC_sg_io_reg2dp_y_extension),
    .io_reg2dp_weight_width_ext(NV_NVDLA_CSC_sg_io_reg2dp_weight_width_ext),
    .io_reg2dp_weight_height_ext(NV_NVDLA_CSC_sg_io_reg2dp_weight_height_ext),
    .io_reg2dp_weight_channel_ext(NV_NVDLA_CSC_sg_io_reg2dp_weight_channel_ext),
    .io_reg2dp_weight_kernel(NV_NVDLA_CSC_sg_io_reg2dp_weight_kernel),
    .io_reg2dp_dataout_width(NV_NVDLA_CSC_sg_io_reg2dp_dataout_width),
    .io_reg2dp_dataout_height(NV_NVDLA_CSC_sg_io_reg2dp_dataout_height),
    .io_reg2dp_data_bank(NV_NVDLA_CSC_sg_io_reg2dp_data_bank),
    .io_reg2dp_weight_bank(NV_NVDLA_CSC_sg_io_reg2dp_weight_bank),
    .io_reg2dp_atomics(NV_NVDLA_CSC_sg_io_reg2dp_atomics),
    .io_reg2dp_rls_slices(NV_NVDLA_CSC_sg_io_reg2dp_rls_slices),
    .io_dp2reg_done(NV_NVDLA_CSC_sg_io_dp2reg_done)
  );
  NV_NVDLA_CSC_wl NV_NVDLA_CSC_wl ( // @[NV_NVDLA_csc.scala 129:22:@23683.4]
    .reset(NV_NVDLA_CSC_wl_reset),
    .io_nvdla_core_clk(NV_NVDLA_CSC_wl_io_nvdla_core_clk),
    .io_nvdla_core_ng_clk(NV_NVDLA_CSC_wl_io_nvdla_core_ng_clk),
    .io_sg2wl_pd_valid(NV_NVDLA_CSC_wl_io_sg2wl_pd_valid),
    .io_sg2wl_pd_bits(NV_NVDLA_CSC_wl_io_sg2wl_pd_bits),
    .io_sg2wl_reuse_rls(NV_NVDLA_CSC_wl_io_sg2wl_reuse_rls),
    .io_sc_state(NV_NVDLA_CSC_wl_io_sc_state),
    .io_sc2cdma_wt_pending_req(NV_NVDLA_CSC_wl_io_sc2cdma_wt_pending_req),
    .io_sc2cdma_wt_updt_valid(NV_NVDLA_CSC_wl_io_sc2cdma_wt_updt_valid),
    .io_sc2cdma_wt_updt_bits_entries(NV_NVDLA_CSC_wl_io_sc2cdma_wt_updt_bits_entries),
    .io_sc2cdma_wmb_entries(NV_NVDLA_CSC_wl_io_sc2cdma_wmb_entries),
    .io_sc2buf_wt_rd_addr_valid(NV_NVDLA_CSC_wl_io_sc2buf_wt_rd_addr_valid),
    .io_sc2buf_wt_rd_addr_bits(NV_NVDLA_CSC_wl_io_sc2buf_wt_rd_addr_bits),
    .io_sc2buf_wt_rd_data_valid(NV_NVDLA_CSC_wl_io_sc2buf_wt_rd_data_valid),
    .io_sc2buf_wt_rd_data_bits(NV_NVDLA_CSC_wl_io_sc2buf_wt_rd_data_bits),
    .io_sc2mac_wt_a_valid(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_valid),
    .io_sc2mac_wt_a_bits_sel_0(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_0),
    .io_sc2mac_wt_a_bits_sel_1(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_1),
    .io_sc2mac_wt_a_bits_sel_2(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_2),
    .io_sc2mac_wt_a_bits_sel_3(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_3),
    .io_sc2mac_wt_a_bits_sel_4(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_4),
    .io_sc2mac_wt_a_bits_sel_5(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_5),
    .io_sc2mac_wt_a_bits_sel_6(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_6),
    .io_sc2mac_wt_a_bits_sel_7(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_7),
    .io_sc2mac_wt_a_bits_sel_8(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_8),
    .io_sc2mac_wt_a_bits_sel_9(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_9),
    .io_sc2mac_wt_a_bits_sel_10(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_10),
    .io_sc2mac_wt_a_bits_sel_11(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_11),
    .io_sc2mac_wt_a_bits_sel_12(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_12),
    .io_sc2mac_wt_a_bits_sel_13(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_13),
    .io_sc2mac_wt_a_bits_sel_14(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_14),
    .io_sc2mac_wt_a_bits_sel_15(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_15),
    .io_sc2mac_wt_a_bits_mask_0(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_0),
    .io_sc2mac_wt_a_bits_mask_1(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_1),
    .io_sc2mac_wt_a_bits_mask_2(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_2),
    .io_sc2mac_wt_a_bits_mask_3(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_3),
    .io_sc2mac_wt_a_bits_mask_4(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_4),
    .io_sc2mac_wt_a_bits_mask_5(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_5),
    .io_sc2mac_wt_a_bits_mask_6(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_6),
    .io_sc2mac_wt_a_bits_mask_7(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_7),
    .io_sc2mac_wt_a_bits_mask_8(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_8),
    .io_sc2mac_wt_a_bits_mask_9(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_9),
    .io_sc2mac_wt_a_bits_mask_10(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_10),
    .io_sc2mac_wt_a_bits_mask_11(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_11),
    .io_sc2mac_wt_a_bits_mask_12(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_12),
    .io_sc2mac_wt_a_bits_mask_13(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_13),
    .io_sc2mac_wt_a_bits_mask_14(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_14),
    .io_sc2mac_wt_a_bits_mask_15(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_15),
    .io_sc2mac_wt_a_bits_mask_16(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_16),
    .io_sc2mac_wt_a_bits_mask_17(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_17),
    .io_sc2mac_wt_a_bits_mask_18(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_18),
    .io_sc2mac_wt_a_bits_mask_19(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_19),
    .io_sc2mac_wt_a_bits_mask_20(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_20),
    .io_sc2mac_wt_a_bits_mask_21(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_21),
    .io_sc2mac_wt_a_bits_mask_22(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_22),
    .io_sc2mac_wt_a_bits_mask_23(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_23),
    .io_sc2mac_wt_a_bits_mask_24(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_24),
    .io_sc2mac_wt_a_bits_mask_25(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_25),
    .io_sc2mac_wt_a_bits_mask_26(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_26),
    .io_sc2mac_wt_a_bits_mask_27(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_27),
    .io_sc2mac_wt_a_bits_mask_28(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_28),
    .io_sc2mac_wt_a_bits_mask_29(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_29),
    .io_sc2mac_wt_a_bits_mask_30(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_30),
    .io_sc2mac_wt_a_bits_mask_31(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_31),
    .io_sc2mac_wt_a_bits_mask_32(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_32),
    .io_sc2mac_wt_a_bits_mask_33(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_33),
    .io_sc2mac_wt_a_bits_mask_34(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_34),
    .io_sc2mac_wt_a_bits_mask_35(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_35),
    .io_sc2mac_wt_a_bits_mask_36(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_36),
    .io_sc2mac_wt_a_bits_mask_37(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_37),
    .io_sc2mac_wt_a_bits_mask_38(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_38),
    .io_sc2mac_wt_a_bits_mask_39(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_39),
    .io_sc2mac_wt_a_bits_mask_40(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_40),
    .io_sc2mac_wt_a_bits_mask_41(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_41),
    .io_sc2mac_wt_a_bits_mask_42(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_42),
    .io_sc2mac_wt_a_bits_mask_43(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_43),
    .io_sc2mac_wt_a_bits_mask_44(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_44),
    .io_sc2mac_wt_a_bits_mask_45(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_45),
    .io_sc2mac_wt_a_bits_mask_46(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_46),
    .io_sc2mac_wt_a_bits_mask_47(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_47),
    .io_sc2mac_wt_a_bits_mask_48(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_48),
    .io_sc2mac_wt_a_bits_mask_49(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_49),
    .io_sc2mac_wt_a_bits_mask_50(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_50),
    .io_sc2mac_wt_a_bits_mask_51(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_51),
    .io_sc2mac_wt_a_bits_mask_52(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_52),
    .io_sc2mac_wt_a_bits_mask_53(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_53),
    .io_sc2mac_wt_a_bits_mask_54(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_54),
    .io_sc2mac_wt_a_bits_mask_55(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_55),
    .io_sc2mac_wt_a_bits_mask_56(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_56),
    .io_sc2mac_wt_a_bits_mask_57(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_57),
    .io_sc2mac_wt_a_bits_mask_58(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_58),
    .io_sc2mac_wt_a_bits_mask_59(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_59),
    .io_sc2mac_wt_a_bits_mask_60(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_60),
    .io_sc2mac_wt_a_bits_mask_61(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_61),
    .io_sc2mac_wt_a_bits_mask_62(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_62),
    .io_sc2mac_wt_a_bits_mask_63(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_63),
    .io_sc2mac_wt_a_bits_data_0(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_0),
    .io_sc2mac_wt_a_bits_data_1(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_1),
    .io_sc2mac_wt_a_bits_data_2(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_2),
    .io_sc2mac_wt_a_bits_data_3(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_3),
    .io_sc2mac_wt_a_bits_data_4(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_4),
    .io_sc2mac_wt_a_bits_data_5(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_5),
    .io_sc2mac_wt_a_bits_data_6(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_6),
    .io_sc2mac_wt_a_bits_data_7(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_7),
    .io_sc2mac_wt_a_bits_data_8(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_8),
    .io_sc2mac_wt_a_bits_data_9(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_9),
    .io_sc2mac_wt_a_bits_data_10(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_10),
    .io_sc2mac_wt_a_bits_data_11(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_11),
    .io_sc2mac_wt_a_bits_data_12(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_12),
    .io_sc2mac_wt_a_bits_data_13(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_13),
    .io_sc2mac_wt_a_bits_data_14(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_14),
    .io_sc2mac_wt_a_bits_data_15(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_15),
    .io_sc2mac_wt_a_bits_data_16(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_16),
    .io_sc2mac_wt_a_bits_data_17(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_17),
    .io_sc2mac_wt_a_bits_data_18(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_18),
    .io_sc2mac_wt_a_bits_data_19(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_19),
    .io_sc2mac_wt_a_bits_data_20(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_20),
    .io_sc2mac_wt_a_bits_data_21(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_21),
    .io_sc2mac_wt_a_bits_data_22(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_22),
    .io_sc2mac_wt_a_bits_data_23(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_23),
    .io_sc2mac_wt_a_bits_data_24(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_24),
    .io_sc2mac_wt_a_bits_data_25(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_25),
    .io_sc2mac_wt_a_bits_data_26(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_26),
    .io_sc2mac_wt_a_bits_data_27(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_27),
    .io_sc2mac_wt_a_bits_data_28(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_28),
    .io_sc2mac_wt_a_bits_data_29(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_29),
    .io_sc2mac_wt_a_bits_data_30(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_30),
    .io_sc2mac_wt_a_bits_data_31(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_31),
    .io_sc2mac_wt_a_bits_data_32(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_32),
    .io_sc2mac_wt_a_bits_data_33(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_33),
    .io_sc2mac_wt_a_bits_data_34(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_34),
    .io_sc2mac_wt_a_bits_data_35(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_35),
    .io_sc2mac_wt_a_bits_data_36(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_36),
    .io_sc2mac_wt_a_bits_data_37(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_37),
    .io_sc2mac_wt_a_bits_data_38(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_38),
    .io_sc2mac_wt_a_bits_data_39(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_39),
    .io_sc2mac_wt_a_bits_data_40(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_40),
    .io_sc2mac_wt_a_bits_data_41(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_41),
    .io_sc2mac_wt_a_bits_data_42(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_42),
    .io_sc2mac_wt_a_bits_data_43(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_43),
    .io_sc2mac_wt_a_bits_data_44(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_44),
    .io_sc2mac_wt_a_bits_data_45(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_45),
    .io_sc2mac_wt_a_bits_data_46(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_46),
    .io_sc2mac_wt_a_bits_data_47(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_47),
    .io_sc2mac_wt_a_bits_data_48(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_48),
    .io_sc2mac_wt_a_bits_data_49(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_49),
    .io_sc2mac_wt_a_bits_data_50(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_50),
    .io_sc2mac_wt_a_bits_data_51(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_51),
    .io_sc2mac_wt_a_bits_data_52(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_52),
    .io_sc2mac_wt_a_bits_data_53(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_53),
    .io_sc2mac_wt_a_bits_data_54(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_54),
    .io_sc2mac_wt_a_bits_data_55(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_55),
    .io_sc2mac_wt_a_bits_data_56(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_56),
    .io_sc2mac_wt_a_bits_data_57(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_57),
    .io_sc2mac_wt_a_bits_data_58(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_58),
    .io_sc2mac_wt_a_bits_data_59(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_59),
    .io_sc2mac_wt_a_bits_data_60(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_60),
    .io_sc2mac_wt_a_bits_data_61(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_61),
    .io_sc2mac_wt_a_bits_data_62(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_62),
    .io_sc2mac_wt_a_bits_data_63(NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_63),
    .io_sc2mac_wt_b_valid(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_valid),
    .io_sc2mac_wt_b_bits_sel_0(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_0),
    .io_sc2mac_wt_b_bits_sel_1(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_1),
    .io_sc2mac_wt_b_bits_sel_2(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_2),
    .io_sc2mac_wt_b_bits_sel_3(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_3),
    .io_sc2mac_wt_b_bits_sel_4(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_4),
    .io_sc2mac_wt_b_bits_sel_5(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_5),
    .io_sc2mac_wt_b_bits_sel_6(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_6),
    .io_sc2mac_wt_b_bits_sel_7(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_7),
    .io_sc2mac_wt_b_bits_sel_8(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_8),
    .io_sc2mac_wt_b_bits_sel_9(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_9),
    .io_sc2mac_wt_b_bits_sel_10(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_10),
    .io_sc2mac_wt_b_bits_sel_11(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_11),
    .io_sc2mac_wt_b_bits_sel_12(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_12),
    .io_sc2mac_wt_b_bits_sel_13(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_13),
    .io_sc2mac_wt_b_bits_sel_14(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_14),
    .io_sc2mac_wt_b_bits_sel_15(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_15),
    .io_sc2mac_wt_b_bits_mask_0(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_0),
    .io_sc2mac_wt_b_bits_mask_1(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_1),
    .io_sc2mac_wt_b_bits_mask_2(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_2),
    .io_sc2mac_wt_b_bits_mask_3(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_3),
    .io_sc2mac_wt_b_bits_mask_4(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_4),
    .io_sc2mac_wt_b_bits_mask_5(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_5),
    .io_sc2mac_wt_b_bits_mask_6(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_6),
    .io_sc2mac_wt_b_bits_mask_7(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_7),
    .io_sc2mac_wt_b_bits_mask_8(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_8),
    .io_sc2mac_wt_b_bits_mask_9(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_9),
    .io_sc2mac_wt_b_bits_mask_10(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_10),
    .io_sc2mac_wt_b_bits_mask_11(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_11),
    .io_sc2mac_wt_b_bits_mask_12(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_12),
    .io_sc2mac_wt_b_bits_mask_13(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_13),
    .io_sc2mac_wt_b_bits_mask_14(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_14),
    .io_sc2mac_wt_b_bits_mask_15(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_15),
    .io_sc2mac_wt_b_bits_mask_16(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_16),
    .io_sc2mac_wt_b_bits_mask_17(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_17),
    .io_sc2mac_wt_b_bits_mask_18(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_18),
    .io_sc2mac_wt_b_bits_mask_19(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_19),
    .io_sc2mac_wt_b_bits_mask_20(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_20),
    .io_sc2mac_wt_b_bits_mask_21(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_21),
    .io_sc2mac_wt_b_bits_mask_22(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_22),
    .io_sc2mac_wt_b_bits_mask_23(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_23),
    .io_sc2mac_wt_b_bits_mask_24(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_24),
    .io_sc2mac_wt_b_bits_mask_25(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_25),
    .io_sc2mac_wt_b_bits_mask_26(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_26),
    .io_sc2mac_wt_b_bits_mask_27(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_27),
    .io_sc2mac_wt_b_bits_mask_28(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_28),
    .io_sc2mac_wt_b_bits_mask_29(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_29),
    .io_sc2mac_wt_b_bits_mask_30(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_30),
    .io_sc2mac_wt_b_bits_mask_31(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_31),
    .io_sc2mac_wt_b_bits_mask_32(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_32),
    .io_sc2mac_wt_b_bits_mask_33(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_33),
    .io_sc2mac_wt_b_bits_mask_34(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_34),
    .io_sc2mac_wt_b_bits_mask_35(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_35),
    .io_sc2mac_wt_b_bits_mask_36(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_36),
    .io_sc2mac_wt_b_bits_mask_37(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_37),
    .io_sc2mac_wt_b_bits_mask_38(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_38),
    .io_sc2mac_wt_b_bits_mask_39(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_39),
    .io_sc2mac_wt_b_bits_mask_40(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_40),
    .io_sc2mac_wt_b_bits_mask_41(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_41),
    .io_sc2mac_wt_b_bits_mask_42(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_42),
    .io_sc2mac_wt_b_bits_mask_43(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_43),
    .io_sc2mac_wt_b_bits_mask_44(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_44),
    .io_sc2mac_wt_b_bits_mask_45(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_45),
    .io_sc2mac_wt_b_bits_mask_46(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_46),
    .io_sc2mac_wt_b_bits_mask_47(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_47),
    .io_sc2mac_wt_b_bits_mask_48(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_48),
    .io_sc2mac_wt_b_bits_mask_49(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_49),
    .io_sc2mac_wt_b_bits_mask_50(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_50),
    .io_sc2mac_wt_b_bits_mask_51(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_51),
    .io_sc2mac_wt_b_bits_mask_52(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_52),
    .io_sc2mac_wt_b_bits_mask_53(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_53),
    .io_sc2mac_wt_b_bits_mask_54(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_54),
    .io_sc2mac_wt_b_bits_mask_55(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_55),
    .io_sc2mac_wt_b_bits_mask_56(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_56),
    .io_sc2mac_wt_b_bits_mask_57(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_57),
    .io_sc2mac_wt_b_bits_mask_58(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_58),
    .io_sc2mac_wt_b_bits_mask_59(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_59),
    .io_sc2mac_wt_b_bits_mask_60(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_60),
    .io_sc2mac_wt_b_bits_mask_61(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_61),
    .io_sc2mac_wt_b_bits_mask_62(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_62),
    .io_sc2mac_wt_b_bits_mask_63(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_63),
    .io_sc2mac_wt_b_bits_data_0(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_0),
    .io_sc2mac_wt_b_bits_data_1(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_1),
    .io_sc2mac_wt_b_bits_data_2(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_2),
    .io_sc2mac_wt_b_bits_data_3(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_3),
    .io_sc2mac_wt_b_bits_data_4(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_4),
    .io_sc2mac_wt_b_bits_data_5(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_5),
    .io_sc2mac_wt_b_bits_data_6(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_6),
    .io_sc2mac_wt_b_bits_data_7(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_7),
    .io_sc2mac_wt_b_bits_data_8(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_8),
    .io_sc2mac_wt_b_bits_data_9(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_9),
    .io_sc2mac_wt_b_bits_data_10(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_10),
    .io_sc2mac_wt_b_bits_data_11(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_11),
    .io_sc2mac_wt_b_bits_data_12(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_12),
    .io_sc2mac_wt_b_bits_data_13(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_13),
    .io_sc2mac_wt_b_bits_data_14(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_14),
    .io_sc2mac_wt_b_bits_data_15(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_15),
    .io_sc2mac_wt_b_bits_data_16(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_16),
    .io_sc2mac_wt_b_bits_data_17(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_17),
    .io_sc2mac_wt_b_bits_data_18(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_18),
    .io_sc2mac_wt_b_bits_data_19(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_19),
    .io_sc2mac_wt_b_bits_data_20(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_20),
    .io_sc2mac_wt_b_bits_data_21(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_21),
    .io_sc2mac_wt_b_bits_data_22(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_22),
    .io_sc2mac_wt_b_bits_data_23(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_23),
    .io_sc2mac_wt_b_bits_data_24(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_24),
    .io_sc2mac_wt_b_bits_data_25(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_25),
    .io_sc2mac_wt_b_bits_data_26(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_26),
    .io_sc2mac_wt_b_bits_data_27(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_27),
    .io_sc2mac_wt_b_bits_data_28(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_28),
    .io_sc2mac_wt_b_bits_data_29(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_29),
    .io_sc2mac_wt_b_bits_data_30(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_30),
    .io_sc2mac_wt_b_bits_data_31(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_31),
    .io_sc2mac_wt_b_bits_data_32(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_32),
    .io_sc2mac_wt_b_bits_data_33(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_33),
    .io_sc2mac_wt_b_bits_data_34(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_34),
    .io_sc2mac_wt_b_bits_data_35(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_35),
    .io_sc2mac_wt_b_bits_data_36(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_36),
    .io_sc2mac_wt_b_bits_data_37(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_37),
    .io_sc2mac_wt_b_bits_data_38(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_38),
    .io_sc2mac_wt_b_bits_data_39(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_39),
    .io_sc2mac_wt_b_bits_data_40(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_40),
    .io_sc2mac_wt_b_bits_data_41(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_41),
    .io_sc2mac_wt_b_bits_data_42(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_42),
    .io_sc2mac_wt_b_bits_data_43(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_43),
    .io_sc2mac_wt_b_bits_data_44(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_44),
    .io_sc2mac_wt_b_bits_data_45(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_45),
    .io_sc2mac_wt_b_bits_data_46(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_46),
    .io_sc2mac_wt_b_bits_data_47(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_47),
    .io_sc2mac_wt_b_bits_data_48(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_48),
    .io_sc2mac_wt_b_bits_data_49(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_49),
    .io_sc2mac_wt_b_bits_data_50(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_50),
    .io_sc2mac_wt_b_bits_data_51(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_51),
    .io_sc2mac_wt_b_bits_data_52(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_52),
    .io_sc2mac_wt_b_bits_data_53(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_53),
    .io_sc2mac_wt_b_bits_data_54(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_54),
    .io_sc2mac_wt_b_bits_data_55(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_55),
    .io_sc2mac_wt_b_bits_data_56(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_56),
    .io_sc2mac_wt_b_bits_data_57(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_57),
    .io_sc2mac_wt_b_bits_data_58(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_58),
    .io_sc2mac_wt_b_bits_data_59(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_59),
    .io_sc2mac_wt_b_bits_data_60(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_60),
    .io_sc2mac_wt_b_bits_data_61(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_61),
    .io_sc2mac_wt_b_bits_data_62(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_62),
    .io_sc2mac_wt_b_bits_data_63(NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_63),
    .io_reg2dp_op_en(NV_NVDLA_CSC_wl_io_reg2dp_op_en),
    .io_reg2dp_y_extension(NV_NVDLA_CSC_wl_io_reg2dp_y_extension),
    .io_reg2dp_skip_weight_rls(NV_NVDLA_CSC_wl_io_reg2dp_skip_weight_rls),
    .io_reg2dp_weight_format(NV_NVDLA_CSC_wl_io_reg2dp_weight_format),
    .io_reg2dp_weight_bytes(NV_NVDLA_CSC_wl_io_reg2dp_weight_bytes),
    .io_reg2dp_wmb_bytes(NV_NVDLA_CSC_wl_io_reg2dp_wmb_bytes),
    .io_reg2dp_data_bank(NV_NVDLA_CSC_wl_io_reg2dp_data_bank),
    .io_reg2dp_weight_bank(NV_NVDLA_CSC_wl_io_reg2dp_weight_bank)
  );
  NV_NVDLA_CSC_dl NV_NVDLA_CSC_dl ( // @[NV_NVDLA_csc.scala 161:22:@24006.4]
    .reset(NV_NVDLA_CSC_dl_reset),
    .io_nvdla_core_clk(NV_NVDLA_CSC_dl_io_nvdla_core_clk),
    .io_nvdla_core_ng_clk(NV_NVDLA_CSC_dl_io_nvdla_core_ng_clk),
    .io_sc_state(NV_NVDLA_CSC_dl_io_sc_state),
    .io_sg2dl_pd_valid(NV_NVDLA_CSC_dl_io_sg2dl_pd_valid),
    .io_sg2dl_reuse_rls(NV_NVDLA_CSC_dl_io_sg2dl_reuse_rls),
    .io_sc2cdma_dat_pending_req(NV_NVDLA_CSC_dl_io_sc2cdma_dat_pending_req),
    .io_sc2cdma_dat_updt_valid(NV_NVDLA_CSC_dl_io_sc2cdma_dat_updt_valid),
    .io_sc2cdma_dat_updt_bits_entries(NV_NVDLA_CSC_dl_io_sc2cdma_dat_updt_bits_entries),
    .io_sc2cdma_dat_updt_bits_slices(NV_NVDLA_CSC_dl_io_sc2cdma_dat_updt_bits_slices),
    .io_sc2buf_dat_rd_addr_valid(NV_NVDLA_CSC_dl_io_sc2buf_dat_rd_addr_valid),
    .io_sc2buf_dat_rd_addr_bits(NV_NVDLA_CSC_dl_io_sc2buf_dat_rd_addr_bits),
    .io_sc2buf_dat_rd_data_valid(NV_NVDLA_CSC_dl_io_sc2buf_dat_rd_data_valid),
    .io_sc2buf_dat_rd_data_bits(NV_NVDLA_CSC_dl_io_sc2buf_dat_rd_data_bits),
    .io_sc2mac_dat_a_valid(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_valid),
    .io_sc2mac_dat_a_bits_mask_0(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_0),
    .io_sc2mac_dat_a_bits_mask_1(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_1),
    .io_sc2mac_dat_a_bits_mask_2(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_2),
    .io_sc2mac_dat_a_bits_mask_3(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_3),
    .io_sc2mac_dat_a_bits_mask_4(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_4),
    .io_sc2mac_dat_a_bits_mask_5(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_5),
    .io_sc2mac_dat_a_bits_mask_6(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_6),
    .io_sc2mac_dat_a_bits_mask_7(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_7),
    .io_sc2mac_dat_a_bits_mask_8(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_8),
    .io_sc2mac_dat_a_bits_mask_9(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_9),
    .io_sc2mac_dat_a_bits_mask_10(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_10),
    .io_sc2mac_dat_a_bits_mask_11(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_11),
    .io_sc2mac_dat_a_bits_mask_12(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_12),
    .io_sc2mac_dat_a_bits_mask_13(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_13),
    .io_sc2mac_dat_a_bits_mask_14(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_14),
    .io_sc2mac_dat_a_bits_mask_15(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_15),
    .io_sc2mac_dat_a_bits_mask_16(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_16),
    .io_sc2mac_dat_a_bits_mask_17(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_17),
    .io_sc2mac_dat_a_bits_mask_18(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_18),
    .io_sc2mac_dat_a_bits_mask_19(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_19),
    .io_sc2mac_dat_a_bits_mask_20(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_20),
    .io_sc2mac_dat_a_bits_mask_21(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_21),
    .io_sc2mac_dat_a_bits_mask_22(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_22),
    .io_sc2mac_dat_a_bits_mask_23(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_23),
    .io_sc2mac_dat_a_bits_mask_24(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_24),
    .io_sc2mac_dat_a_bits_mask_25(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_25),
    .io_sc2mac_dat_a_bits_mask_26(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_26),
    .io_sc2mac_dat_a_bits_mask_27(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_27),
    .io_sc2mac_dat_a_bits_mask_28(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_28),
    .io_sc2mac_dat_a_bits_mask_29(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_29),
    .io_sc2mac_dat_a_bits_mask_30(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_30),
    .io_sc2mac_dat_a_bits_mask_31(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_31),
    .io_sc2mac_dat_a_bits_mask_32(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_32),
    .io_sc2mac_dat_a_bits_mask_33(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_33),
    .io_sc2mac_dat_a_bits_mask_34(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_34),
    .io_sc2mac_dat_a_bits_mask_35(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_35),
    .io_sc2mac_dat_a_bits_mask_36(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_36),
    .io_sc2mac_dat_a_bits_mask_37(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_37),
    .io_sc2mac_dat_a_bits_mask_38(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_38),
    .io_sc2mac_dat_a_bits_mask_39(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_39),
    .io_sc2mac_dat_a_bits_mask_40(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_40),
    .io_sc2mac_dat_a_bits_mask_41(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_41),
    .io_sc2mac_dat_a_bits_mask_42(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_42),
    .io_sc2mac_dat_a_bits_mask_43(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_43),
    .io_sc2mac_dat_a_bits_mask_44(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_44),
    .io_sc2mac_dat_a_bits_mask_45(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_45),
    .io_sc2mac_dat_a_bits_mask_46(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_46),
    .io_sc2mac_dat_a_bits_mask_47(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_47),
    .io_sc2mac_dat_a_bits_mask_48(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_48),
    .io_sc2mac_dat_a_bits_mask_49(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_49),
    .io_sc2mac_dat_a_bits_mask_50(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_50),
    .io_sc2mac_dat_a_bits_mask_51(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_51),
    .io_sc2mac_dat_a_bits_mask_52(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_52),
    .io_sc2mac_dat_a_bits_mask_53(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_53),
    .io_sc2mac_dat_a_bits_mask_54(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_54),
    .io_sc2mac_dat_a_bits_mask_55(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_55),
    .io_sc2mac_dat_a_bits_mask_56(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_56),
    .io_sc2mac_dat_a_bits_mask_57(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_57),
    .io_sc2mac_dat_a_bits_mask_58(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_58),
    .io_sc2mac_dat_a_bits_mask_59(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_59),
    .io_sc2mac_dat_a_bits_mask_60(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_60),
    .io_sc2mac_dat_a_bits_mask_61(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_61),
    .io_sc2mac_dat_a_bits_mask_62(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_62),
    .io_sc2mac_dat_a_bits_mask_63(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_63),
    .io_sc2mac_dat_a_bits_data_0(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_0),
    .io_sc2mac_dat_a_bits_data_1(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_1),
    .io_sc2mac_dat_a_bits_data_2(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_2),
    .io_sc2mac_dat_a_bits_data_3(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_3),
    .io_sc2mac_dat_a_bits_data_4(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_4),
    .io_sc2mac_dat_a_bits_data_5(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_5),
    .io_sc2mac_dat_a_bits_data_6(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_6),
    .io_sc2mac_dat_a_bits_data_7(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_7),
    .io_sc2mac_dat_a_bits_data_8(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_8),
    .io_sc2mac_dat_a_bits_data_9(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_9),
    .io_sc2mac_dat_a_bits_data_10(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_10),
    .io_sc2mac_dat_a_bits_data_11(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_11),
    .io_sc2mac_dat_a_bits_data_12(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_12),
    .io_sc2mac_dat_a_bits_data_13(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_13),
    .io_sc2mac_dat_a_bits_data_14(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_14),
    .io_sc2mac_dat_a_bits_data_15(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_15),
    .io_sc2mac_dat_a_bits_data_16(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_16),
    .io_sc2mac_dat_a_bits_data_17(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_17),
    .io_sc2mac_dat_a_bits_data_18(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_18),
    .io_sc2mac_dat_a_bits_data_19(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_19),
    .io_sc2mac_dat_a_bits_data_20(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_20),
    .io_sc2mac_dat_a_bits_data_21(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_21),
    .io_sc2mac_dat_a_bits_data_22(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_22),
    .io_sc2mac_dat_a_bits_data_23(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_23),
    .io_sc2mac_dat_a_bits_data_24(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_24),
    .io_sc2mac_dat_a_bits_data_25(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_25),
    .io_sc2mac_dat_a_bits_data_26(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_26),
    .io_sc2mac_dat_a_bits_data_27(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_27),
    .io_sc2mac_dat_a_bits_data_28(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_28),
    .io_sc2mac_dat_a_bits_data_29(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_29),
    .io_sc2mac_dat_a_bits_data_30(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_30),
    .io_sc2mac_dat_a_bits_data_31(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_31),
    .io_sc2mac_dat_a_bits_data_32(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_32),
    .io_sc2mac_dat_a_bits_data_33(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_33),
    .io_sc2mac_dat_a_bits_data_34(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_34),
    .io_sc2mac_dat_a_bits_data_35(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_35),
    .io_sc2mac_dat_a_bits_data_36(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_36),
    .io_sc2mac_dat_a_bits_data_37(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_37),
    .io_sc2mac_dat_a_bits_data_38(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_38),
    .io_sc2mac_dat_a_bits_data_39(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_39),
    .io_sc2mac_dat_a_bits_data_40(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_40),
    .io_sc2mac_dat_a_bits_data_41(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_41),
    .io_sc2mac_dat_a_bits_data_42(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_42),
    .io_sc2mac_dat_a_bits_data_43(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_43),
    .io_sc2mac_dat_a_bits_data_44(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_44),
    .io_sc2mac_dat_a_bits_data_45(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_45),
    .io_sc2mac_dat_a_bits_data_46(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_46),
    .io_sc2mac_dat_a_bits_data_47(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_47),
    .io_sc2mac_dat_a_bits_data_48(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_48),
    .io_sc2mac_dat_a_bits_data_49(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_49),
    .io_sc2mac_dat_a_bits_data_50(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_50),
    .io_sc2mac_dat_a_bits_data_51(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_51),
    .io_sc2mac_dat_a_bits_data_52(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_52),
    .io_sc2mac_dat_a_bits_data_53(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_53),
    .io_sc2mac_dat_a_bits_data_54(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_54),
    .io_sc2mac_dat_a_bits_data_55(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_55),
    .io_sc2mac_dat_a_bits_data_56(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_56),
    .io_sc2mac_dat_a_bits_data_57(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_57),
    .io_sc2mac_dat_a_bits_data_58(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_58),
    .io_sc2mac_dat_a_bits_data_59(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_59),
    .io_sc2mac_dat_a_bits_data_60(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_60),
    .io_sc2mac_dat_a_bits_data_61(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_61),
    .io_sc2mac_dat_a_bits_data_62(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_62),
    .io_sc2mac_dat_a_bits_data_63(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_63),
    .io_sc2mac_dat_a_bits_pd(NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_pd),
    .io_sc2mac_dat_b_valid(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_valid),
    .io_sc2mac_dat_b_bits_mask_0(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_0),
    .io_sc2mac_dat_b_bits_mask_1(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_1),
    .io_sc2mac_dat_b_bits_mask_2(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_2),
    .io_sc2mac_dat_b_bits_mask_3(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_3),
    .io_sc2mac_dat_b_bits_mask_4(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_4),
    .io_sc2mac_dat_b_bits_mask_5(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_5),
    .io_sc2mac_dat_b_bits_mask_6(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_6),
    .io_sc2mac_dat_b_bits_mask_7(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_7),
    .io_sc2mac_dat_b_bits_mask_8(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_8),
    .io_sc2mac_dat_b_bits_mask_9(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_9),
    .io_sc2mac_dat_b_bits_mask_10(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_10),
    .io_sc2mac_dat_b_bits_mask_11(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_11),
    .io_sc2mac_dat_b_bits_mask_12(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_12),
    .io_sc2mac_dat_b_bits_mask_13(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_13),
    .io_sc2mac_dat_b_bits_mask_14(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_14),
    .io_sc2mac_dat_b_bits_mask_15(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_15),
    .io_sc2mac_dat_b_bits_mask_16(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_16),
    .io_sc2mac_dat_b_bits_mask_17(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_17),
    .io_sc2mac_dat_b_bits_mask_18(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_18),
    .io_sc2mac_dat_b_bits_mask_19(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_19),
    .io_sc2mac_dat_b_bits_mask_20(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_20),
    .io_sc2mac_dat_b_bits_mask_21(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_21),
    .io_sc2mac_dat_b_bits_mask_22(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_22),
    .io_sc2mac_dat_b_bits_mask_23(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_23),
    .io_sc2mac_dat_b_bits_mask_24(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_24),
    .io_sc2mac_dat_b_bits_mask_25(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_25),
    .io_sc2mac_dat_b_bits_mask_26(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_26),
    .io_sc2mac_dat_b_bits_mask_27(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_27),
    .io_sc2mac_dat_b_bits_mask_28(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_28),
    .io_sc2mac_dat_b_bits_mask_29(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_29),
    .io_sc2mac_dat_b_bits_mask_30(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_30),
    .io_sc2mac_dat_b_bits_mask_31(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_31),
    .io_sc2mac_dat_b_bits_mask_32(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_32),
    .io_sc2mac_dat_b_bits_mask_33(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_33),
    .io_sc2mac_dat_b_bits_mask_34(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_34),
    .io_sc2mac_dat_b_bits_mask_35(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_35),
    .io_sc2mac_dat_b_bits_mask_36(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_36),
    .io_sc2mac_dat_b_bits_mask_37(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_37),
    .io_sc2mac_dat_b_bits_mask_38(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_38),
    .io_sc2mac_dat_b_bits_mask_39(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_39),
    .io_sc2mac_dat_b_bits_mask_40(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_40),
    .io_sc2mac_dat_b_bits_mask_41(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_41),
    .io_sc2mac_dat_b_bits_mask_42(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_42),
    .io_sc2mac_dat_b_bits_mask_43(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_43),
    .io_sc2mac_dat_b_bits_mask_44(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_44),
    .io_sc2mac_dat_b_bits_mask_45(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_45),
    .io_sc2mac_dat_b_bits_mask_46(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_46),
    .io_sc2mac_dat_b_bits_mask_47(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_47),
    .io_sc2mac_dat_b_bits_mask_48(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_48),
    .io_sc2mac_dat_b_bits_mask_49(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_49),
    .io_sc2mac_dat_b_bits_mask_50(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_50),
    .io_sc2mac_dat_b_bits_mask_51(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_51),
    .io_sc2mac_dat_b_bits_mask_52(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_52),
    .io_sc2mac_dat_b_bits_mask_53(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_53),
    .io_sc2mac_dat_b_bits_mask_54(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_54),
    .io_sc2mac_dat_b_bits_mask_55(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_55),
    .io_sc2mac_dat_b_bits_mask_56(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_56),
    .io_sc2mac_dat_b_bits_mask_57(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_57),
    .io_sc2mac_dat_b_bits_mask_58(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_58),
    .io_sc2mac_dat_b_bits_mask_59(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_59),
    .io_sc2mac_dat_b_bits_mask_60(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_60),
    .io_sc2mac_dat_b_bits_mask_61(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_61),
    .io_sc2mac_dat_b_bits_mask_62(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_62),
    .io_sc2mac_dat_b_bits_mask_63(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_63),
    .io_sc2mac_dat_b_bits_data_0(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_0),
    .io_sc2mac_dat_b_bits_data_1(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_1),
    .io_sc2mac_dat_b_bits_data_2(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_2),
    .io_sc2mac_dat_b_bits_data_3(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_3),
    .io_sc2mac_dat_b_bits_data_4(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_4),
    .io_sc2mac_dat_b_bits_data_5(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_5),
    .io_sc2mac_dat_b_bits_data_6(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_6),
    .io_sc2mac_dat_b_bits_data_7(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_7),
    .io_sc2mac_dat_b_bits_data_8(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_8),
    .io_sc2mac_dat_b_bits_data_9(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_9),
    .io_sc2mac_dat_b_bits_data_10(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_10),
    .io_sc2mac_dat_b_bits_data_11(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_11),
    .io_sc2mac_dat_b_bits_data_12(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_12),
    .io_sc2mac_dat_b_bits_data_13(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_13),
    .io_sc2mac_dat_b_bits_data_14(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_14),
    .io_sc2mac_dat_b_bits_data_15(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_15),
    .io_sc2mac_dat_b_bits_data_16(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_16),
    .io_sc2mac_dat_b_bits_data_17(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_17),
    .io_sc2mac_dat_b_bits_data_18(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_18),
    .io_sc2mac_dat_b_bits_data_19(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_19),
    .io_sc2mac_dat_b_bits_data_20(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_20),
    .io_sc2mac_dat_b_bits_data_21(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_21),
    .io_sc2mac_dat_b_bits_data_22(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_22),
    .io_sc2mac_dat_b_bits_data_23(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_23),
    .io_sc2mac_dat_b_bits_data_24(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_24),
    .io_sc2mac_dat_b_bits_data_25(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_25),
    .io_sc2mac_dat_b_bits_data_26(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_26),
    .io_sc2mac_dat_b_bits_data_27(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_27),
    .io_sc2mac_dat_b_bits_data_28(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_28),
    .io_sc2mac_dat_b_bits_data_29(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_29),
    .io_sc2mac_dat_b_bits_data_30(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_30),
    .io_sc2mac_dat_b_bits_data_31(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_31),
    .io_sc2mac_dat_b_bits_data_32(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_32),
    .io_sc2mac_dat_b_bits_data_33(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_33),
    .io_sc2mac_dat_b_bits_data_34(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_34),
    .io_sc2mac_dat_b_bits_data_35(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_35),
    .io_sc2mac_dat_b_bits_data_36(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_36),
    .io_sc2mac_dat_b_bits_data_37(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_37),
    .io_sc2mac_dat_b_bits_data_38(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_38),
    .io_sc2mac_dat_b_bits_data_39(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_39),
    .io_sc2mac_dat_b_bits_data_40(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_40),
    .io_sc2mac_dat_b_bits_data_41(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_41),
    .io_sc2mac_dat_b_bits_data_42(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_42),
    .io_sc2mac_dat_b_bits_data_43(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_43),
    .io_sc2mac_dat_b_bits_data_44(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_44),
    .io_sc2mac_dat_b_bits_data_45(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_45),
    .io_sc2mac_dat_b_bits_data_46(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_46),
    .io_sc2mac_dat_b_bits_data_47(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_47),
    .io_sc2mac_dat_b_bits_data_48(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_48),
    .io_sc2mac_dat_b_bits_data_49(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_49),
    .io_sc2mac_dat_b_bits_data_50(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_50),
    .io_sc2mac_dat_b_bits_data_51(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_51),
    .io_sc2mac_dat_b_bits_data_52(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_52),
    .io_sc2mac_dat_b_bits_data_53(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_53),
    .io_sc2mac_dat_b_bits_data_54(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_54),
    .io_sc2mac_dat_b_bits_data_55(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_55),
    .io_sc2mac_dat_b_bits_data_56(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_56),
    .io_sc2mac_dat_b_bits_data_57(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_57),
    .io_sc2mac_dat_b_bits_data_58(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_58),
    .io_sc2mac_dat_b_bits_data_59(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_59),
    .io_sc2mac_dat_b_bits_data_60(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_60),
    .io_sc2mac_dat_b_bits_data_61(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_61),
    .io_sc2mac_dat_b_bits_data_62(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_62),
    .io_sc2mac_dat_b_bits_data_63(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_63),
    .io_sc2mac_dat_b_bits_pd(NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_pd),
    .io_reg2dp_op_en(NV_NVDLA_CSC_dl_io_reg2dp_op_en),
    .io_reg2dp_conv_mode(NV_NVDLA_CSC_dl_io_reg2dp_conv_mode),
    .io_reg2dp_datain_format(NV_NVDLA_CSC_dl_io_reg2dp_datain_format),
    .io_reg2dp_skip_data_rls(NV_NVDLA_CSC_dl_io_reg2dp_skip_data_rls),
    .io_reg2dp_datain_channel_ext(NV_NVDLA_CSC_dl_io_reg2dp_datain_channel_ext),
    .io_reg2dp_datain_height_ext(NV_NVDLA_CSC_dl_io_reg2dp_datain_height_ext),
    .io_reg2dp_datain_width_ext(NV_NVDLA_CSC_dl_io_reg2dp_datain_width_ext),
    .io_reg2dp_y_extension(NV_NVDLA_CSC_dl_io_reg2dp_y_extension),
    .io_reg2dp_weight_channel_ext(NV_NVDLA_CSC_dl_io_reg2dp_weight_channel_ext),
    .io_reg2dp_entries(NV_NVDLA_CSC_dl_io_reg2dp_entries),
    .io_reg2dp_dataout_width(NV_NVDLA_CSC_dl_io_reg2dp_dataout_width),
    .io_reg2dp_rls_slices(NV_NVDLA_CSC_dl_io_reg2dp_rls_slices),
    .io_reg2dp_conv_x_stride_ext(NV_NVDLA_CSC_dl_io_reg2dp_conv_x_stride_ext),
    .io_reg2dp_conv_y_stride_ext(NV_NVDLA_CSC_dl_io_reg2dp_conv_y_stride_ext),
    .io_reg2dp_x_dilation_ext(NV_NVDLA_CSC_dl_io_reg2dp_x_dilation_ext),
    .io_reg2dp_y_dilation_ext(NV_NVDLA_CSC_dl_io_reg2dp_y_dilation_ext),
    .io_reg2dp_pad_left(NV_NVDLA_CSC_dl_io_reg2dp_pad_left),
    .io_reg2dp_pad_top(NV_NVDLA_CSC_dl_io_reg2dp_pad_top),
    .io_reg2dp_pad_value(NV_NVDLA_CSC_dl_io_reg2dp_pad_value),
    .io_reg2dp_data_bank(NV_NVDLA_CSC_dl_io_reg2dp_data_bank)
  );
  NV_NVDLA_slcg NV_NVDLA_slcg ( // @[NV_NVDLA_csc.scala 205:41:@24309.4]
    .io_nvdla_clock_nvdla_core_clk(NV_NVDLA_slcg_io_nvdla_clock_nvdla_core_clk),
    .io_nvdla_core_gated_clk(NV_NVDLA_slcg_io_nvdla_core_gated_clk)
  );
  NV_NVDLA_slcg NV_NVDLA_slcg_1 ( // @[NV_NVDLA_csc.scala 205:41:@24312.4]
    .io_nvdla_clock_nvdla_core_clk(NV_NVDLA_slcg_1_io_nvdla_clock_nvdla_core_clk),
    .io_nvdla_core_gated_clk(NV_NVDLA_slcg_1_io_nvdla_core_gated_clk)
  );
  NV_NVDLA_slcg NV_NVDLA_slcg_2 ( // @[NV_NVDLA_csc.scala 205:41:@24315.4]
    .io_nvdla_clock_nvdla_core_clk(NV_NVDLA_slcg_2_io_nvdla_clock_nvdla_core_clk),
    .io_nvdla_core_gated_clk(NV_NVDLA_slcg_2_io_nvdla_core_gated_clk)
  );
  assign io_sc2cdma_dat_pending_req = NV_NVDLA_CSC_sg_io_sc2cdma_dat_pending_req; // @[NV_NVDLA_csc.scala 98:32:@23658.4]
  assign io_sc2cdma_wt_pending_req = NV_NVDLA_CSC_sg_io_sc2cdma_wt_pending_req; // @[NV_NVDLA_csc.scala 99:31:@23659.4]
  assign io_sc2cdma_dat_updt_valid = NV_NVDLA_CSC_dl_io_sc2cdma_dat_updt_valid; // @[NV_NVDLA_csc.scala 169:25:@24021.4]
  assign io_sc2cdma_dat_updt_bits_entries = NV_NVDLA_CSC_dl_io_sc2cdma_dat_updt_bits_entries; // @[NV_NVDLA_csc.scala 169:25:@24020.4]
  assign io_sc2cdma_dat_updt_bits_slices = NV_NVDLA_CSC_dl_io_sc2cdma_dat_updt_bits_slices; // @[NV_NVDLA_csc.scala 169:25:@24019.4]
  assign io_sc2cdma_wt_updt_valid = NV_NVDLA_CSC_wl_io_sc2cdma_wt_updt_valid; // @[NV_NVDLA_csc.scala 138:24:@23698.4]
  assign io_sc2cdma_wt_updt_bits_entries = NV_NVDLA_CSC_wl_io_sc2cdma_wt_updt_bits_entries; // @[NV_NVDLA_csc.scala 138:24:@23697.4]
  assign io_sc2cdma_wt_updt_bits_kernels = 14'h0; // @[NV_NVDLA_csc.scala 138:24:@23696.4]
  assign io_sc2cdma_wmb_entries = NV_NVDLA_CSC_wl_io_sc2cdma_wmb_entries; // @[NV_NVDLA_csc.scala 141:28:@23704.4]
  assign io_csb2csc_req_ready = 1'h1; // @[NV_NVDLA_csc.scala 80:26:@23643.4]
  assign io_csb2csc_resp_valid = NV_NVDLA_CSC_regfile_io_csb2csc_resp_valid; // @[NV_NVDLA_csc.scala 80:26:@23640.4]
  assign io_csb2csc_resp_bits = NV_NVDLA_CSC_regfile_io_csb2csc_resp_bits; // @[NV_NVDLA_csc.scala 80:26:@23639.4]
  assign io_sc2buf_dat_rd_addr_valid = NV_NVDLA_CSC_dl_io_sc2buf_dat_rd_addr_valid; // @[NV_NVDLA_csc.scala 170:22:@24025.4]
  assign io_sc2buf_dat_rd_addr_bits = NV_NVDLA_CSC_dl_io_sc2buf_dat_rd_addr_bits; // @[NV_NVDLA_csc.scala 170:22:@24024.4]
  assign io_sc2buf_wt_rd_addr_valid = NV_NVDLA_CSC_wl_io_sc2buf_wt_rd_addr_valid; // @[NV_NVDLA_csc.scala 139:21:@23702.4]
  assign io_sc2buf_wt_rd_addr_bits = NV_NVDLA_CSC_wl_io_sc2buf_wt_rd_addr_bits; // @[NV_NVDLA_csc.scala 139:21:@23701.4]
  assign io_sc2mac_dat_a_valid = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_valid; // @[NV_NVDLA_csc.scala 171:21:@24155.4]
  assign io_sc2mac_dat_a_bits_mask_0 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_0; // @[NV_NVDLA_csc.scala 171:21:@24091.4]
  assign io_sc2mac_dat_a_bits_mask_1 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_1; // @[NV_NVDLA_csc.scala 171:21:@24092.4]
  assign io_sc2mac_dat_a_bits_mask_2 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_2; // @[NV_NVDLA_csc.scala 171:21:@24093.4]
  assign io_sc2mac_dat_a_bits_mask_3 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_3; // @[NV_NVDLA_csc.scala 171:21:@24094.4]
  assign io_sc2mac_dat_a_bits_mask_4 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_4; // @[NV_NVDLA_csc.scala 171:21:@24095.4]
  assign io_sc2mac_dat_a_bits_mask_5 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_5; // @[NV_NVDLA_csc.scala 171:21:@24096.4]
  assign io_sc2mac_dat_a_bits_mask_6 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_6; // @[NV_NVDLA_csc.scala 171:21:@24097.4]
  assign io_sc2mac_dat_a_bits_mask_7 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_7; // @[NV_NVDLA_csc.scala 171:21:@24098.4]
  assign io_sc2mac_dat_a_bits_mask_8 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_8; // @[NV_NVDLA_csc.scala 171:21:@24099.4]
  assign io_sc2mac_dat_a_bits_mask_9 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_9; // @[NV_NVDLA_csc.scala 171:21:@24100.4]
  assign io_sc2mac_dat_a_bits_mask_10 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_10; // @[NV_NVDLA_csc.scala 171:21:@24101.4]
  assign io_sc2mac_dat_a_bits_mask_11 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_11; // @[NV_NVDLA_csc.scala 171:21:@24102.4]
  assign io_sc2mac_dat_a_bits_mask_12 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_12; // @[NV_NVDLA_csc.scala 171:21:@24103.4]
  assign io_sc2mac_dat_a_bits_mask_13 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_13; // @[NV_NVDLA_csc.scala 171:21:@24104.4]
  assign io_sc2mac_dat_a_bits_mask_14 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_14; // @[NV_NVDLA_csc.scala 171:21:@24105.4]
  assign io_sc2mac_dat_a_bits_mask_15 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_15; // @[NV_NVDLA_csc.scala 171:21:@24106.4]
  assign io_sc2mac_dat_a_bits_mask_16 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_16; // @[NV_NVDLA_csc.scala 171:21:@24107.4]
  assign io_sc2mac_dat_a_bits_mask_17 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_17; // @[NV_NVDLA_csc.scala 171:21:@24108.4]
  assign io_sc2mac_dat_a_bits_mask_18 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_18; // @[NV_NVDLA_csc.scala 171:21:@24109.4]
  assign io_sc2mac_dat_a_bits_mask_19 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_19; // @[NV_NVDLA_csc.scala 171:21:@24110.4]
  assign io_sc2mac_dat_a_bits_mask_20 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_20; // @[NV_NVDLA_csc.scala 171:21:@24111.4]
  assign io_sc2mac_dat_a_bits_mask_21 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_21; // @[NV_NVDLA_csc.scala 171:21:@24112.4]
  assign io_sc2mac_dat_a_bits_mask_22 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_22; // @[NV_NVDLA_csc.scala 171:21:@24113.4]
  assign io_sc2mac_dat_a_bits_mask_23 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_23; // @[NV_NVDLA_csc.scala 171:21:@24114.4]
  assign io_sc2mac_dat_a_bits_mask_24 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_24; // @[NV_NVDLA_csc.scala 171:21:@24115.4]
  assign io_sc2mac_dat_a_bits_mask_25 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_25; // @[NV_NVDLA_csc.scala 171:21:@24116.4]
  assign io_sc2mac_dat_a_bits_mask_26 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_26; // @[NV_NVDLA_csc.scala 171:21:@24117.4]
  assign io_sc2mac_dat_a_bits_mask_27 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_27; // @[NV_NVDLA_csc.scala 171:21:@24118.4]
  assign io_sc2mac_dat_a_bits_mask_28 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_28; // @[NV_NVDLA_csc.scala 171:21:@24119.4]
  assign io_sc2mac_dat_a_bits_mask_29 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_29; // @[NV_NVDLA_csc.scala 171:21:@24120.4]
  assign io_sc2mac_dat_a_bits_mask_30 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_30; // @[NV_NVDLA_csc.scala 171:21:@24121.4]
  assign io_sc2mac_dat_a_bits_mask_31 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_31; // @[NV_NVDLA_csc.scala 171:21:@24122.4]
  assign io_sc2mac_dat_a_bits_mask_32 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_32; // @[NV_NVDLA_csc.scala 171:21:@24123.4]
  assign io_sc2mac_dat_a_bits_mask_33 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_33; // @[NV_NVDLA_csc.scala 171:21:@24124.4]
  assign io_sc2mac_dat_a_bits_mask_34 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_34; // @[NV_NVDLA_csc.scala 171:21:@24125.4]
  assign io_sc2mac_dat_a_bits_mask_35 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_35; // @[NV_NVDLA_csc.scala 171:21:@24126.4]
  assign io_sc2mac_dat_a_bits_mask_36 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_36; // @[NV_NVDLA_csc.scala 171:21:@24127.4]
  assign io_sc2mac_dat_a_bits_mask_37 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_37; // @[NV_NVDLA_csc.scala 171:21:@24128.4]
  assign io_sc2mac_dat_a_bits_mask_38 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_38; // @[NV_NVDLA_csc.scala 171:21:@24129.4]
  assign io_sc2mac_dat_a_bits_mask_39 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_39; // @[NV_NVDLA_csc.scala 171:21:@24130.4]
  assign io_sc2mac_dat_a_bits_mask_40 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_40; // @[NV_NVDLA_csc.scala 171:21:@24131.4]
  assign io_sc2mac_dat_a_bits_mask_41 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_41; // @[NV_NVDLA_csc.scala 171:21:@24132.4]
  assign io_sc2mac_dat_a_bits_mask_42 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_42; // @[NV_NVDLA_csc.scala 171:21:@24133.4]
  assign io_sc2mac_dat_a_bits_mask_43 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_43; // @[NV_NVDLA_csc.scala 171:21:@24134.4]
  assign io_sc2mac_dat_a_bits_mask_44 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_44; // @[NV_NVDLA_csc.scala 171:21:@24135.4]
  assign io_sc2mac_dat_a_bits_mask_45 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_45; // @[NV_NVDLA_csc.scala 171:21:@24136.4]
  assign io_sc2mac_dat_a_bits_mask_46 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_46; // @[NV_NVDLA_csc.scala 171:21:@24137.4]
  assign io_sc2mac_dat_a_bits_mask_47 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_47; // @[NV_NVDLA_csc.scala 171:21:@24138.4]
  assign io_sc2mac_dat_a_bits_mask_48 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_48; // @[NV_NVDLA_csc.scala 171:21:@24139.4]
  assign io_sc2mac_dat_a_bits_mask_49 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_49; // @[NV_NVDLA_csc.scala 171:21:@24140.4]
  assign io_sc2mac_dat_a_bits_mask_50 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_50; // @[NV_NVDLA_csc.scala 171:21:@24141.4]
  assign io_sc2mac_dat_a_bits_mask_51 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_51; // @[NV_NVDLA_csc.scala 171:21:@24142.4]
  assign io_sc2mac_dat_a_bits_mask_52 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_52; // @[NV_NVDLA_csc.scala 171:21:@24143.4]
  assign io_sc2mac_dat_a_bits_mask_53 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_53; // @[NV_NVDLA_csc.scala 171:21:@24144.4]
  assign io_sc2mac_dat_a_bits_mask_54 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_54; // @[NV_NVDLA_csc.scala 171:21:@24145.4]
  assign io_sc2mac_dat_a_bits_mask_55 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_55; // @[NV_NVDLA_csc.scala 171:21:@24146.4]
  assign io_sc2mac_dat_a_bits_mask_56 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_56; // @[NV_NVDLA_csc.scala 171:21:@24147.4]
  assign io_sc2mac_dat_a_bits_mask_57 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_57; // @[NV_NVDLA_csc.scala 171:21:@24148.4]
  assign io_sc2mac_dat_a_bits_mask_58 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_58; // @[NV_NVDLA_csc.scala 171:21:@24149.4]
  assign io_sc2mac_dat_a_bits_mask_59 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_59; // @[NV_NVDLA_csc.scala 171:21:@24150.4]
  assign io_sc2mac_dat_a_bits_mask_60 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_60; // @[NV_NVDLA_csc.scala 171:21:@24151.4]
  assign io_sc2mac_dat_a_bits_mask_61 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_61; // @[NV_NVDLA_csc.scala 171:21:@24152.4]
  assign io_sc2mac_dat_a_bits_mask_62 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_62; // @[NV_NVDLA_csc.scala 171:21:@24153.4]
  assign io_sc2mac_dat_a_bits_mask_63 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_mask_63; // @[NV_NVDLA_csc.scala 171:21:@24154.4]
  assign io_sc2mac_dat_a_bits_data_0 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_0; // @[NV_NVDLA_csc.scala 171:21:@24027.4]
  assign io_sc2mac_dat_a_bits_data_1 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_1; // @[NV_NVDLA_csc.scala 171:21:@24028.4]
  assign io_sc2mac_dat_a_bits_data_2 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_2; // @[NV_NVDLA_csc.scala 171:21:@24029.4]
  assign io_sc2mac_dat_a_bits_data_3 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_3; // @[NV_NVDLA_csc.scala 171:21:@24030.4]
  assign io_sc2mac_dat_a_bits_data_4 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_4; // @[NV_NVDLA_csc.scala 171:21:@24031.4]
  assign io_sc2mac_dat_a_bits_data_5 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_5; // @[NV_NVDLA_csc.scala 171:21:@24032.4]
  assign io_sc2mac_dat_a_bits_data_6 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_6; // @[NV_NVDLA_csc.scala 171:21:@24033.4]
  assign io_sc2mac_dat_a_bits_data_7 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_7; // @[NV_NVDLA_csc.scala 171:21:@24034.4]
  assign io_sc2mac_dat_a_bits_data_8 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_8; // @[NV_NVDLA_csc.scala 171:21:@24035.4]
  assign io_sc2mac_dat_a_bits_data_9 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_9; // @[NV_NVDLA_csc.scala 171:21:@24036.4]
  assign io_sc2mac_dat_a_bits_data_10 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_10; // @[NV_NVDLA_csc.scala 171:21:@24037.4]
  assign io_sc2mac_dat_a_bits_data_11 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_11; // @[NV_NVDLA_csc.scala 171:21:@24038.4]
  assign io_sc2mac_dat_a_bits_data_12 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_12; // @[NV_NVDLA_csc.scala 171:21:@24039.4]
  assign io_sc2mac_dat_a_bits_data_13 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_13; // @[NV_NVDLA_csc.scala 171:21:@24040.4]
  assign io_sc2mac_dat_a_bits_data_14 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_14; // @[NV_NVDLA_csc.scala 171:21:@24041.4]
  assign io_sc2mac_dat_a_bits_data_15 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_15; // @[NV_NVDLA_csc.scala 171:21:@24042.4]
  assign io_sc2mac_dat_a_bits_data_16 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_16; // @[NV_NVDLA_csc.scala 171:21:@24043.4]
  assign io_sc2mac_dat_a_bits_data_17 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_17; // @[NV_NVDLA_csc.scala 171:21:@24044.4]
  assign io_sc2mac_dat_a_bits_data_18 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_18; // @[NV_NVDLA_csc.scala 171:21:@24045.4]
  assign io_sc2mac_dat_a_bits_data_19 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_19; // @[NV_NVDLA_csc.scala 171:21:@24046.4]
  assign io_sc2mac_dat_a_bits_data_20 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_20; // @[NV_NVDLA_csc.scala 171:21:@24047.4]
  assign io_sc2mac_dat_a_bits_data_21 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_21; // @[NV_NVDLA_csc.scala 171:21:@24048.4]
  assign io_sc2mac_dat_a_bits_data_22 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_22; // @[NV_NVDLA_csc.scala 171:21:@24049.4]
  assign io_sc2mac_dat_a_bits_data_23 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_23; // @[NV_NVDLA_csc.scala 171:21:@24050.4]
  assign io_sc2mac_dat_a_bits_data_24 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_24; // @[NV_NVDLA_csc.scala 171:21:@24051.4]
  assign io_sc2mac_dat_a_bits_data_25 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_25; // @[NV_NVDLA_csc.scala 171:21:@24052.4]
  assign io_sc2mac_dat_a_bits_data_26 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_26; // @[NV_NVDLA_csc.scala 171:21:@24053.4]
  assign io_sc2mac_dat_a_bits_data_27 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_27; // @[NV_NVDLA_csc.scala 171:21:@24054.4]
  assign io_sc2mac_dat_a_bits_data_28 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_28; // @[NV_NVDLA_csc.scala 171:21:@24055.4]
  assign io_sc2mac_dat_a_bits_data_29 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_29; // @[NV_NVDLA_csc.scala 171:21:@24056.4]
  assign io_sc2mac_dat_a_bits_data_30 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_30; // @[NV_NVDLA_csc.scala 171:21:@24057.4]
  assign io_sc2mac_dat_a_bits_data_31 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_31; // @[NV_NVDLA_csc.scala 171:21:@24058.4]
  assign io_sc2mac_dat_a_bits_data_32 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_32; // @[NV_NVDLA_csc.scala 171:21:@24059.4]
  assign io_sc2mac_dat_a_bits_data_33 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_33; // @[NV_NVDLA_csc.scala 171:21:@24060.4]
  assign io_sc2mac_dat_a_bits_data_34 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_34; // @[NV_NVDLA_csc.scala 171:21:@24061.4]
  assign io_sc2mac_dat_a_bits_data_35 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_35; // @[NV_NVDLA_csc.scala 171:21:@24062.4]
  assign io_sc2mac_dat_a_bits_data_36 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_36; // @[NV_NVDLA_csc.scala 171:21:@24063.4]
  assign io_sc2mac_dat_a_bits_data_37 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_37; // @[NV_NVDLA_csc.scala 171:21:@24064.4]
  assign io_sc2mac_dat_a_bits_data_38 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_38; // @[NV_NVDLA_csc.scala 171:21:@24065.4]
  assign io_sc2mac_dat_a_bits_data_39 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_39; // @[NV_NVDLA_csc.scala 171:21:@24066.4]
  assign io_sc2mac_dat_a_bits_data_40 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_40; // @[NV_NVDLA_csc.scala 171:21:@24067.4]
  assign io_sc2mac_dat_a_bits_data_41 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_41; // @[NV_NVDLA_csc.scala 171:21:@24068.4]
  assign io_sc2mac_dat_a_bits_data_42 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_42; // @[NV_NVDLA_csc.scala 171:21:@24069.4]
  assign io_sc2mac_dat_a_bits_data_43 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_43; // @[NV_NVDLA_csc.scala 171:21:@24070.4]
  assign io_sc2mac_dat_a_bits_data_44 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_44; // @[NV_NVDLA_csc.scala 171:21:@24071.4]
  assign io_sc2mac_dat_a_bits_data_45 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_45; // @[NV_NVDLA_csc.scala 171:21:@24072.4]
  assign io_sc2mac_dat_a_bits_data_46 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_46; // @[NV_NVDLA_csc.scala 171:21:@24073.4]
  assign io_sc2mac_dat_a_bits_data_47 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_47; // @[NV_NVDLA_csc.scala 171:21:@24074.4]
  assign io_sc2mac_dat_a_bits_data_48 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_48; // @[NV_NVDLA_csc.scala 171:21:@24075.4]
  assign io_sc2mac_dat_a_bits_data_49 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_49; // @[NV_NVDLA_csc.scala 171:21:@24076.4]
  assign io_sc2mac_dat_a_bits_data_50 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_50; // @[NV_NVDLA_csc.scala 171:21:@24077.4]
  assign io_sc2mac_dat_a_bits_data_51 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_51; // @[NV_NVDLA_csc.scala 171:21:@24078.4]
  assign io_sc2mac_dat_a_bits_data_52 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_52; // @[NV_NVDLA_csc.scala 171:21:@24079.4]
  assign io_sc2mac_dat_a_bits_data_53 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_53; // @[NV_NVDLA_csc.scala 171:21:@24080.4]
  assign io_sc2mac_dat_a_bits_data_54 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_54; // @[NV_NVDLA_csc.scala 171:21:@24081.4]
  assign io_sc2mac_dat_a_bits_data_55 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_55; // @[NV_NVDLA_csc.scala 171:21:@24082.4]
  assign io_sc2mac_dat_a_bits_data_56 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_56; // @[NV_NVDLA_csc.scala 171:21:@24083.4]
  assign io_sc2mac_dat_a_bits_data_57 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_57; // @[NV_NVDLA_csc.scala 171:21:@24084.4]
  assign io_sc2mac_dat_a_bits_data_58 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_58; // @[NV_NVDLA_csc.scala 171:21:@24085.4]
  assign io_sc2mac_dat_a_bits_data_59 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_59; // @[NV_NVDLA_csc.scala 171:21:@24086.4]
  assign io_sc2mac_dat_a_bits_data_60 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_60; // @[NV_NVDLA_csc.scala 171:21:@24087.4]
  assign io_sc2mac_dat_a_bits_data_61 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_61; // @[NV_NVDLA_csc.scala 171:21:@24088.4]
  assign io_sc2mac_dat_a_bits_data_62 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_62; // @[NV_NVDLA_csc.scala 171:21:@24089.4]
  assign io_sc2mac_dat_a_bits_data_63 = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_data_63; // @[NV_NVDLA_csc.scala 171:21:@24090.4]
  assign io_sc2mac_dat_a_bits_pd = NV_NVDLA_CSC_dl_io_sc2mac_dat_a_bits_pd; // @[NV_NVDLA_csc.scala 171:21:@24026.4]
  assign io_sc2mac_dat_b_valid = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_valid; // @[NV_NVDLA_csc.scala 172:21:@24285.4]
  assign io_sc2mac_dat_b_bits_mask_0 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_0; // @[NV_NVDLA_csc.scala 172:21:@24221.4]
  assign io_sc2mac_dat_b_bits_mask_1 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_1; // @[NV_NVDLA_csc.scala 172:21:@24222.4]
  assign io_sc2mac_dat_b_bits_mask_2 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_2; // @[NV_NVDLA_csc.scala 172:21:@24223.4]
  assign io_sc2mac_dat_b_bits_mask_3 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_3; // @[NV_NVDLA_csc.scala 172:21:@24224.4]
  assign io_sc2mac_dat_b_bits_mask_4 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_4; // @[NV_NVDLA_csc.scala 172:21:@24225.4]
  assign io_sc2mac_dat_b_bits_mask_5 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_5; // @[NV_NVDLA_csc.scala 172:21:@24226.4]
  assign io_sc2mac_dat_b_bits_mask_6 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_6; // @[NV_NVDLA_csc.scala 172:21:@24227.4]
  assign io_sc2mac_dat_b_bits_mask_7 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_7; // @[NV_NVDLA_csc.scala 172:21:@24228.4]
  assign io_sc2mac_dat_b_bits_mask_8 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_8; // @[NV_NVDLA_csc.scala 172:21:@24229.4]
  assign io_sc2mac_dat_b_bits_mask_9 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_9; // @[NV_NVDLA_csc.scala 172:21:@24230.4]
  assign io_sc2mac_dat_b_bits_mask_10 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_10; // @[NV_NVDLA_csc.scala 172:21:@24231.4]
  assign io_sc2mac_dat_b_bits_mask_11 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_11; // @[NV_NVDLA_csc.scala 172:21:@24232.4]
  assign io_sc2mac_dat_b_bits_mask_12 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_12; // @[NV_NVDLA_csc.scala 172:21:@24233.4]
  assign io_sc2mac_dat_b_bits_mask_13 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_13; // @[NV_NVDLA_csc.scala 172:21:@24234.4]
  assign io_sc2mac_dat_b_bits_mask_14 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_14; // @[NV_NVDLA_csc.scala 172:21:@24235.4]
  assign io_sc2mac_dat_b_bits_mask_15 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_15; // @[NV_NVDLA_csc.scala 172:21:@24236.4]
  assign io_sc2mac_dat_b_bits_mask_16 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_16; // @[NV_NVDLA_csc.scala 172:21:@24237.4]
  assign io_sc2mac_dat_b_bits_mask_17 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_17; // @[NV_NVDLA_csc.scala 172:21:@24238.4]
  assign io_sc2mac_dat_b_bits_mask_18 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_18; // @[NV_NVDLA_csc.scala 172:21:@24239.4]
  assign io_sc2mac_dat_b_bits_mask_19 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_19; // @[NV_NVDLA_csc.scala 172:21:@24240.4]
  assign io_sc2mac_dat_b_bits_mask_20 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_20; // @[NV_NVDLA_csc.scala 172:21:@24241.4]
  assign io_sc2mac_dat_b_bits_mask_21 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_21; // @[NV_NVDLA_csc.scala 172:21:@24242.4]
  assign io_sc2mac_dat_b_bits_mask_22 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_22; // @[NV_NVDLA_csc.scala 172:21:@24243.4]
  assign io_sc2mac_dat_b_bits_mask_23 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_23; // @[NV_NVDLA_csc.scala 172:21:@24244.4]
  assign io_sc2mac_dat_b_bits_mask_24 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_24; // @[NV_NVDLA_csc.scala 172:21:@24245.4]
  assign io_sc2mac_dat_b_bits_mask_25 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_25; // @[NV_NVDLA_csc.scala 172:21:@24246.4]
  assign io_sc2mac_dat_b_bits_mask_26 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_26; // @[NV_NVDLA_csc.scala 172:21:@24247.4]
  assign io_sc2mac_dat_b_bits_mask_27 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_27; // @[NV_NVDLA_csc.scala 172:21:@24248.4]
  assign io_sc2mac_dat_b_bits_mask_28 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_28; // @[NV_NVDLA_csc.scala 172:21:@24249.4]
  assign io_sc2mac_dat_b_bits_mask_29 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_29; // @[NV_NVDLA_csc.scala 172:21:@24250.4]
  assign io_sc2mac_dat_b_bits_mask_30 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_30; // @[NV_NVDLA_csc.scala 172:21:@24251.4]
  assign io_sc2mac_dat_b_bits_mask_31 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_31; // @[NV_NVDLA_csc.scala 172:21:@24252.4]
  assign io_sc2mac_dat_b_bits_mask_32 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_32; // @[NV_NVDLA_csc.scala 172:21:@24253.4]
  assign io_sc2mac_dat_b_bits_mask_33 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_33; // @[NV_NVDLA_csc.scala 172:21:@24254.4]
  assign io_sc2mac_dat_b_bits_mask_34 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_34; // @[NV_NVDLA_csc.scala 172:21:@24255.4]
  assign io_sc2mac_dat_b_bits_mask_35 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_35; // @[NV_NVDLA_csc.scala 172:21:@24256.4]
  assign io_sc2mac_dat_b_bits_mask_36 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_36; // @[NV_NVDLA_csc.scala 172:21:@24257.4]
  assign io_sc2mac_dat_b_bits_mask_37 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_37; // @[NV_NVDLA_csc.scala 172:21:@24258.4]
  assign io_sc2mac_dat_b_bits_mask_38 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_38; // @[NV_NVDLA_csc.scala 172:21:@24259.4]
  assign io_sc2mac_dat_b_bits_mask_39 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_39; // @[NV_NVDLA_csc.scala 172:21:@24260.4]
  assign io_sc2mac_dat_b_bits_mask_40 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_40; // @[NV_NVDLA_csc.scala 172:21:@24261.4]
  assign io_sc2mac_dat_b_bits_mask_41 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_41; // @[NV_NVDLA_csc.scala 172:21:@24262.4]
  assign io_sc2mac_dat_b_bits_mask_42 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_42; // @[NV_NVDLA_csc.scala 172:21:@24263.4]
  assign io_sc2mac_dat_b_bits_mask_43 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_43; // @[NV_NVDLA_csc.scala 172:21:@24264.4]
  assign io_sc2mac_dat_b_bits_mask_44 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_44; // @[NV_NVDLA_csc.scala 172:21:@24265.4]
  assign io_sc2mac_dat_b_bits_mask_45 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_45; // @[NV_NVDLA_csc.scala 172:21:@24266.4]
  assign io_sc2mac_dat_b_bits_mask_46 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_46; // @[NV_NVDLA_csc.scala 172:21:@24267.4]
  assign io_sc2mac_dat_b_bits_mask_47 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_47; // @[NV_NVDLA_csc.scala 172:21:@24268.4]
  assign io_sc2mac_dat_b_bits_mask_48 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_48; // @[NV_NVDLA_csc.scala 172:21:@24269.4]
  assign io_sc2mac_dat_b_bits_mask_49 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_49; // @[NV_NVDLA_csc.scala 172:21:@24270.4]
  assign io_sc2mac_dat_b_bits_mask_50 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_50; // @[NV_NVDLA_csc.scala 172:21:@24271.4]
  assign io_sc2mac_dat_b_bits_mask_51 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_51; // @[NV_NVDLA_csc.scala 172:21:@24272.4]
  assign io_sc2mac_dat_b_bits_mask_52 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_52; // @[NV_NVDLA_csc.scala 172:21:@24273.4]
  assign io_sc2mac_dat_b_bits_mask_53 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_53; // @[NV_NVDLA_csc.scala 172:21:@24274.4]
  assign io_sc2mac_dat_b_bits_mask_54 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_54; // @[NV_NVDLA_csc.scala 172:21:@24275.4]
  assign io_sc2mac_dat_b_bits_mask_55 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_55; // @[NV_NVDLA_csc.scala 172:21:@24276.4]
  assign io_sc2mac_dat_b_bits_mask_56 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_56; // @[NV_NVDLA_csc.scala 172:21:@24277.4]
  assign io_sc2mac_dat_b_bits_mask_57 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_57; // @[NV_NVDLA_csc.scala 172:21:@24278.4]
  assign io_sc2mac_dat_b_bits_mask_58 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_58; // @[NV_NVDLA_csc.scala 172:21:@24279.4]
  assign io_sc2mac_dat_b_bits_mask_59 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_59; // @[NV_NVDLA_csc.scala 172:21:@24280.4]
  assign io_sc2mac_dat_b_bits_mask_60 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_60; // @[NV_NVDLA_csc.scala 172:21:@24281.4]
  assign io_sc2mac_dat_b_bits_mask_61 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_61; // @[NV_NVDLA_csc.scala 172:21:@24282.4]
  assign io_sc2mac_dat_b_bits_mask_62 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_62; // @[NV_NVDLA_csc.scala 172:21:@24283.4]
  assign io_sc2mac_dat_b_bits_mask_63 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_mask_63; // @[NV_NVDLA_csc.scala 172:21:@24284.4]
  assign io_sc2mac_dat_b_bits_data_0 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_0; // @[NV_NVDLA_csc.scala 172:21:@24157.4]
  assign io_sc2mac_dat_b_bits_data_1 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_1; // @[NV_NVDLA_csc.scala 172:21:@24158.4]
  assign io_sc2mac_dat_b_bits_data_2 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_2; // @[NV_NVDLA_csc.scala 172:21:@24159.4]
  assign io_sc2mac_dat_b_bits_data_3 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_3; // @[NV_NVDLA_csc.scala 172:21:@24160.4]
  assign io_sc2mac_dat_b_bits_data_4 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_4; // @[NV_NVDLA_csc.scala 172:21:@24161.4]
  assign io_sc2mac_dat_b_bits_data_5 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_5; // @[NV_NVDLA_csc.scala 172:21:@24162.4]
  assign io_sc2mac_dat_b_bits_data_6 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_6; // @[NV_NVDLA_csc.scala 172:21:@24163.4]
  assign io_sc2mac_dat_b_bits_data_7 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_7; // @[NV_NVDLA_csc.scala 172:21:@24164.4]
  assign io_sc2mac_dat_b_bits_data_8 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_8; // @[NV_NVDLA_csc.scala 172:21:@24165.4]
  assign io_sc2mac_dat_b_bits_data_9 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_9; // @[NV_NVDLA_csc.scala 172:21:@24166.4]
  assign io_sc2mac_dat_b_bits_data_10 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_10; // @[NV_NVDLA_csc.scala 172:21:@24167.4]
  assign io_sc2mac_dat_b_bits_data_11 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_11; // @[NV_NVDLA_csc.scala 172:21:@24168.4]
  assign io_sc2mac_dat_b_bits_data_12 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_12; // @[NV_NVDLA_csc.scala 172:21:@24169.4]
  assign io_sc2mac_dat_b_bits_data_13 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_13; // @[NV_NVDLA_csc.scala 172:21:@24170.4]
  assign io_sc2mac_dat_b_bits_data_14 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_14; // @[NV_NVDLA_csc.scala 172:21:@24171.4]
  assign io_sc2mac_dat_b_bits_data_15 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_15; // @[NV_NVDLA_csc.scala 172:21:@24172.4]
  assign io_sc2mac_dat_b_bits_data_16 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_16; // @[NV_NVDLA_csc.scala 172:21:@24173.4]
  assign io_sc2mac_dat_b_bits_data_17 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_17; // @[NV_NVDLA_csc.scala 172:21:@24174.4]
  assign io_sc2mac_dat_b_bits_data_18 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_18; // @[NV_NVDLA_csc.scala 172:21:@24175.4]
  assign io_sc2mac_dat_b_bits_data_19 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_19; // @[NV_NVDLA_csc.scala 172:21:@24176.4]
  assign io_sc2mac_dat_b_bits_data_20 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_20; // @[NV_NVDLA_csc.scala 172:21:@24177.4]
  assign io_sc2mac_dat_b_bits_data_21 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_21; // @[NV_NVDLA_csc.scala 172:21:@24178.4]
  assign io_sc2mac_dat_b_bits_data_22 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_22; // @[NV_NVDLA_csc.scala 172:21:@24179.4]
  assign io_sc2mac_dat_b_bits_data_23 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_23; // @[NV_NVDLA_csc.scala 172:21:@24180.4]
  assign io_sc2mac_dat_b_bits_data_24 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_24; // @[NV_NVDLA_csc.scala 172:21:@24181.4]
  assign io_sc2mac_dat_b_bits_data_25 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_25; // @[NV_NVDLA_csc.scala 172:21:@24182.4]
  assign io_sc2mac_dat_b_bits_data_26 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_26; // @[NV_NVDLA_csc.scala 172:21:@24183.4]
  assign io_sc2mac_dat_b_bits_data_27 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_27; // @[NV_NVDLA_csc.scala 172:21:@24184.4]
  assign io_sc2mac_dat_b_bits_data_28 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_28; // @[NV_NVDLA_csc.scala 172:21:@24185.4]
  assign io_sc2mac_dat_b_bits_data_29 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_29; // @[NV_NVDLA_csc.scala 172:21:@24186.4]
  assign io_sc2mac_dat_b_bits_data_30 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_30; // @[NV_NVDLA_csc.scala 172:21:@24187.4]
  assign io_sc2mac_dat_b_bits_data_31 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_31; // @[NV_NVDLA_csc.scala 172:21:@24188.4]
  assign io_sc2mac_dat_b_bits_data_32 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_32; // @[NV_NVDLA_csc.scala 172:21:@24189.4]
  assign io_sc2mac_dat_b_bits_data_33 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_33; // @[NV_NVDLA_csc.scala 172:21:@24190.4]
  assign io_sc2mac_dat_b_bits_data_34 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_34; // @[NV_NVDLA_csc.scala 172:21:@24191.4]
  assign io_sc2mac_dat_b_bits_data_35 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_35; // @[NV_NVDLA_csc.scala 172:21:@24192.4]
  assign io_sc2mac_dat_b_bits_data_36 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_36; // @[NV_NVDLA_csc.scala 172:21:@24193.4]
  assign io_sc2mac_dat_b_bits_data_37 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_37; // @[NV_NVDLA_csc.scala 172:21:@24194.4]
  assign io_sc2mac_dat_b_bits_data_38 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_38; // @[NV_NVDLA_csc.scala 172:21:@24195.4]
  assign io_sc2mac_dat_b_bits_data_39 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_39; // @[NV_NVDLA_csc.scala 172:21:@24196.4]
  assign io_sc2mac_dat_b_bits_data_40 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_40; // @[NV_NVDLA_csc.scala 172:21:@24197.4]
  assign io_sc2mac_dat_b_bits_data_41 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_41; // @[NV_NVDLA_csc.scala 172:21:@24198.4]
  assign io_sc2mac_dat_b_bits_data_42 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_42; // @[NV_NVDLA_csc.scala 172:21:@24199.4]
  assign io_sc2mac_dat_b_bits_data_43 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_43; // @[NV_NVDLA_csc.scala 172:21:@24200.4]
  assign io_sc2mac_dat_b_bits_data_44 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_44; // @[NV_NVDLA_csc.scala 172:21:@24201.4]
  assign io_sc2mac_dat_b_bits_data_45 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_45; // @[NV_NVDLA_csc.scala 172:21:@24202.4]
  assign io_sc2mac_dat_b_bits_data_46 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_46; // @[NV_NVDLA_csc.scala 172:21:@24203.4]
  assign io_sc2mac_dat_b_bits_data_47 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_47; // @[NV_NVDLA_csc.scala 172:21:@24204.4]
  assign io_sc2mac_dat_b_bits_data_48 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_48; // @[NV_NVDLA_csc.scala 172:21:@24205.4]
  assign io_sc2mac_dat_b_bits_data_49 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_49; // @[NV_NVDLA_csc.scala 172:21:@24206.4]
  assign io_sc2mac_dat_b_bits_data_50 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_50; // @[NV_NVDLA_csc.scala 172:21:@24207.4]
  assign io_sc2mac_dat_b_bits_data_51 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_51; // @[NV_NVDLA_csc.scala 172:21:@24208.4]
  assign io_sc2mac_dat_b_bits_data_52 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_52; // @[NV_NVDLA_csc.scala 172:21:@24209.4]
  assign io_sc2mac_dat_b_bits_data_53 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_53; // @[NV_NVDLA_csc.scala 172:21:@24210.4]
  assign io_sc2mac_dat_b_bits_data_54 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_54; // @[NV_NVDLA_csc.scala 172:21:@24211.4]
  assign io_sc2mac_dat_b_bits_data_55 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_55; // @[NV_NVDLA_csc.scala 172:21:@24212.4]
  assign io_sc2mac_dat_b_bits_data_56 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_56; // @[NV_NVDLA_csc.scala 172:21:@24213.4]
  assign io_sc2mac_dat_b_bits_data_57 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_57; // @[NV_NVDLA_csc.scala 172:21:@24214.4]
  assign io_sc2mac_dat_b_bits_data_58 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_58; // @[NV_NVDLA_csc.scala 172:21:@24215.4]
  assign io_sc2mac_dat_b_bits_data_59 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_59; // @[NV_NVDLA_csc.scala 172:21:@24216.4]
  assign io_sc2mac_dat_b_bits_data_60 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_60; // @[NV_NVDLA_csc.scala 172:21:@24217.4]
  assign io_sc2mac_dat_b_bits_data_61 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_61; // @[NV_NVDLA_csc.scala 172:21:@24218.4]
  assign io_sc2mac_dat_b_bits_data_62 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_62; // @[NV_NVDLA_csc.scala 172:21:@24219.4]
  assign io_sc2mac_dat_b_bits_data_63 = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_data_63; // @[NV_NVDLA_csc.scala 172:21:@24220.4]
  assign io_sc2mac_dat_b_bits_pd = NV_NVDLA_CSC_dl_io_sc2mac_dat_b_bits_pd; // @[NV_NVDLA_csc.scala 172:21:@24156.4]
  assign io_sc2mac_wt_a_valid = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_valid; // @[NV_NVDLA_csc.scala 142:20:@23849.4]
  assign io_sc2mac_wt_a_bits_sel_0 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_0; // @[NV_NVDLA_csc.scala 142:20:@23833.4]
  assign io_sc2mac_wt_a_bits_sel_1 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_1; // @[NV_NVDLA_csc.scala 142:20:@23834.4]
  assign io_sc2mac_wt_a_bits_sel_2 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_2; // @[NV_NVDLA_csc.scala 142:20:@23835.4]
  assign io_sc2mac_wt_a_bits_sel_3 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_3; // @[NV_NVDLA_csc.scala 142:20:@23836.4]
  assign io_sc2mac_wt_a_bits_sel_4 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_4; // @[NV_NVDLA_csc.scala 142:20:@23837.4]
  assign io_sc2mac_wt_a_bits_sel_5 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_5; // @[NV_NVDLA_csc.scala 142:20:@23838.4]
  assign io_sc2mac_wt_a_bits_sel_6 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_6; // @[NV_NVDLA_csc.scala 142:20:@23839.4]
  assign io_sc2mac_wt_a_bits_sel_7 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_7; // @[NV_NVDLA_csc.scala 142:20:@23840.4]
  assign io_sc2mac_wt_a_bits_sel_8 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_8; // @[NV_NVDLA_csc.scala 142:20:@23841.4]
  assign io_sc2mac_wt_a_bits_sel_9 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_9; // @[NV_NVDLA_csc.scala 142:20:@23842.4]
  assign io_sc2mac_wt_a_bits_sel_10 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_10; // @[NV_NVDLA_csc.scala 142:20:@23843.4]
  assign io_sc2mac_wt_a_bits_sel_11 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_11; // @[NV_NVDLA_csc.scala 142:20:@23844.4]
  assign io_sc2mac_wt_a_bits_sel_12 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_12; // @[NV_NVDLA_csc.scala 142:20:@23845.4]
  assign io_sc2mac_wt_a_bits_sel_13 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_13; // @[NV_NVDLA_csc.scala 142:20:@23846.4]
  assign io_sc2mac_wt_a_bits_sel_14 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_14; // @[NV_NVDLA_csc.scala 142:20:@23847.4]
  assign io_sc2mac_wt_a_bits_sel_15 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_sel_15; // @[NV_NVDLA_csc.scala 142:20:@23848.4]
  assign io_sc2mac_wt_a_bits_mask_0 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_0; // @[NV_NVDLA_csc.scala 142:20:@23769.4]
  assign io_sc2mac_wt_a_bits_mask_1 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_1; // @[NV_NVDLA_csc.scala 142:20:@23770.4]
  assign io_sc2mac_wt_a_bits_mask_2 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_2; // @[NV_NVDLA_csc.scala 142:20:@23771.4]
  assign io_sc2mac_wt_a_bits_mask_3 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_3; // @[NV_NVDLA_csc.scala 142:20:@23772.4]
  assign io_sc2mac_wt_a_bits_mask_4 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_4; // @[NV_NVDLA_csc.scala 142:20:@23773.4]
  assign io_sc2mac_wt_a_bits_mask_5 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_5; // @[NV_NVDLA_csc.scala 142:20:@23774.4]
  assign io_sc2mac_wt_a_bits_mask_6 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_6; // @[NV_NVDLA_csc.scala 142:20:@23775.4]
  assign io_sc2mac_wt_a_bits_mask_7 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_7; // @[NV_NVDLA_csc.scala 142:20:@23776.4]
  assign io_sc2mac_wt_a_bits_mask_8 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_8; // @[NV_NVDLA_csc.scala 142:20:@23777.4]
  assign io_sc2mac_wt_a_bits_mask_9 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_9; // @[NV_NVDLA_csc.scala 142:20:@23778.4]
  assign io_sc2mac_wt_a_bits_mask_10 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_10; // @[NV_NVDLA_csc.scala 142:20:@23779.4]
  assign io_sc2mac_wt_a_bits_mask_11 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_11; // @[NV_NVDLA_csc.scala 142:20:@23780.4]
  assign io_sc2mac_wt_a_bits_mask_12 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_12; // @[NV_NVDLA_csc.scala 142:20:@23781.4]
  assign io_sc2mac_wt_a_bits_mask_13 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_13; // @[NV_NVDLA_csc.scala 142:20:@23782.4]
  assign io_sc2mac_wt_a_bits_mask_14 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_14; // @[NV_NVDLA_csc.scala 142:20:@23783.4]
  assign io_sc2mac_wt_a_bits_mask_15 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_15; // @[NV_NVDLA_csc.scala 142:20:@23784.4]
  assign io_sc2mac_wt_a_bits_mask_16 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_16; // @[NV_NVDLA_csc.scala 142:20:@23785.4]
  assign io_sc2mac_wt_a_bits_mask_17 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_17; // @[NV_NVDLA_csc.scala 142:20:@23786.4]
  assign io_sc2mac_wt_a_bits_mask_18 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_18; // @[NV_NVDLA_csc.scala 142:20:@23787.4]
  assign io_sc2mac_wt_a_bits_mask_19 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_19; // @[NV_NVDLA_csc.scala 142:20:@23788.4]
  assign io_sc2mac_wt_a_bits_mask_20 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_20; // @[NV_NVDLA_csc.scala 142:20:@23789.4]
  assign io_sc2mac_wt_a_bits_mask_21 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_21; // @[NV_NVDLA_csc.scala 142:20:@23790.4]
  assign io_sc2mac_wt_a_bits_mask_22 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_22; // @[NV_NVDLA_csc.scala 142:20:@23791.4]
  assign io_sc2mac_wt_a_bits_mask_23 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_23; // @[NV_NVDLA_csc.scala 142:20:@23792.4]
  assign io_sc2mac_wt_a_bits_mask_24 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_24; // @[NV_NVDLA_csc.scala 142:20:@23793.4]
  assign io_sc2mac_wt_a_bits_mask_25 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_25; // @[NV_NVDLA_csc.scala 142:20:@23794.4]
  assign io_sc2mac_wt_a_bits_mask_26 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_26; // @[NV_NVDLA_csc.scala 142:20:@23795.4]
  assign io_sc2mac_wt_a_bits_mask_27 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_27; // @[NV_NVDLA_csc.scala 142:20:@23796.4]
  assign io_sc2mac_wt_a_bits_mask_28 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_28; // @[NV_NVDLA_csc.scala 142:20:@23797.4]
  assign io_sc2mac_wt_a_bits_mask_29 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_29; // @[NV_NVDLA_csc.scala 142:20:@23798.4]
  assign io_sc2mac_wt_a_bits_mask_30 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_30; // @[NV_NVDLA_csc.scala 142:20:@23799.4]
  assign io_sc2mac_wt_a_bits_mask_31 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_31; // @[NV_NVDLA_csc.scala 142:20:@23800.4]
  assign io_sc2mac_wt_a_bits_mask_32 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_32; // @[NV_NVDLA_csc.scala 142:20:@23801.4]
  assign io_sc2mac_wt_a_bits_mask_33 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_33; // @[NV_NVDLA_csc.scala 142:20:@23802.4]
  assign io_sc2mac_wt_a_bits_mask_34 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_34; // @[NV_NVDLA_csc.scala 142:20:@23803.4]
  assign io_sc2mac_wt_a_bits_mask_35 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_35; // @[NV_NVDLA_csc.scala 142:20:@23804.4]
  assign io_sc2mac_wt_a_bits_mask_36 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_36; // @[NV_NVDLA_csc.scala 142:20:@23805.4]
  assign io_sc2mac_wt_a_bits_mask_37 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_37; // @[NV_NVDLA_csc.scala 142:20:@23806.4]
  assign io_sc2mac_wt_a_bits_mask_38 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_38; // @[NV_NVDLA_csc.scala 142:20:@23807.4]
  assign io_sc2mac_wt_a_bits_mask_39 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_39; // @[NV_NVDLA_csc.scala 142:20:@23808.4]
  assign io_sc2mac_wt_a_bits_mask_40 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_40; // @[NV_NVDLA_csc.scala 142:20:@23809.4]
  assign io_sc2mac_wt_a_bits_mask_41 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_41; // @[NV_NVDLA_csc.scala 142:20:@23810.4]
  assign io_sc2mac_wt_a_bits_mask_42 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_42; // @[NV_NVDLA_csc.scala 142:20:@23811.4]
  assign io_sc2mac_wt_a_bits_mask_43 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_43; // @[NV_NVDLA_csc.scala 142:20:@23812.4]
  assign io_sc2mac_wt_a_bits_mask_44 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_44; // @[NV_NVDLA_csc.scala 142:20:@23813.4]
  assign io_sc2mac_wt_a_bits_mask_45 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_45; // @[NV_NVDLA_csc.scala 142:20:@23814.4]
  assign io_sc2mac_wt_a_bits_mask_46 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_46; // @[NV_NVDLA_csc.scala 142:20:@23815.4]
  assign io_sc2mac_wt_a_bits_mask_47 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_47; // @[NV_NVDLA_csc.scala 142:20:@23816.4]
  assign io_sc2mac_wt_a_bits_mask_48 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_48; // @[NV_NVDLA_csc.scala 142:20:@23817.4]
  assign io_sc2mac_wt_a_bits_mask_49 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_49; // @[NV_NVDLA_csc.scala 142:20:@23818.4]
  assign io_sc2mac_wt_a_bits_mask_50 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_50; // @[NV_NVDLA_csc.scala 142:20:@23819.4]
  assign io_sc2mac_wt_a_bits_mask_51 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_51; // @[NV_NVDLA_csc.scala 142:20:@23820.4]
  assign io_sc2mac_wt_a_bits_mask_52 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_52; // @[NV_NVDLA_csc.scala 142:20:@23821.4]
  assign io_sc2mac_wt_a_bits_mask_53 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_53; // @[NV_NVDLA_csc.scala 142:20:@23822.4]
  assign io_sc2mac_wt_a_bits_mask_54 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_54; // @[NV_NVDLA_csc.scala 142:20:@23823.4]
  assign io_sc2mac_wt_a_bits_mask_55 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_55; // @[NV_NVDLA_csc.scala 142:20:@23824.4]
  assign io_sc2mac_wt_a_bits_mask_56 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_56; // @[NV_NVDLA_csc.scala 142:20:@23825.4]
  assign io_sc2mac_wt_a_bits_mask_57 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_57; // @[NV_NVDLA_csc.scala 142:20:@23826.4]
  assign io_sc2mac_wt_a_bits_mask_58 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_58; // @[NV_NVDLA_csc.scala 142:20:@23827.4]
  assign io_sc2mac_wt_a_bits_mask_59 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_59; // @[NV_NVDLA_csc.scala 142:20:@23828.4]
  assign io_sc2mac_wt_a_bits_mask_60 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_60; // @[NV_NVDLA_csc.scala 142:20:@23829.4]
  assign io_sc2mac_wt_a_bits_mask_61 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_61; // @[NV_NVDLA_csc.scala 142:20:@23830.4]
  assign io_sc2mac_wt_a_bits_mask_62 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_62; // @[NV_NVDLA_csc.scala 142:20:@23831.4]
  assign io_sc2mac_wt_a_bits_mask_63 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_mask_63; // @[NV_NVDLA_csc.scala 142:20:@23832.4]
  assign io_sc2mac_wt_a_bits_data_0 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_0; // @[NV_NVDLA_csc.scala 142:20:@23705.4]
  assign io_sc2mac_wt_a_bits_data_1 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_1; // @[NV_NVDLA_csc.scala 142:20:@23706.4]
  assign io_sc2mac_wt_a_bits_data_2 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_2; // @[NV_NVDLA_csc.scala 142:20:@23707.4]
  assign io_sc2mac_wt_a_bits_data_3 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_3; // @[NV_NVDLA_csc.scala 142:20:@23708.4]
  assign io_sc2mac_wt_a_bits_data_4 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_4; // @[NV_NVDLA_csc.scala 142:20:@23709.4]
  assign io_sc2mac_wt_a_bits_data_5 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_5; // @[NV_NVDLA_csc.scala 142:20:@23710.4]
  assign io_sc2mac_wt_a_bits_data_6 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_6; // @[NV_NVDLA_csc.scala 142:20:@23711.4]
  assign io_sc2mac_wt_a_bits_data_7 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_7; // @[NV_NVDLA_csc.scala 142:20:@23712.4]
  assign io_sc2mac_wt_a_bits_data_8 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_8; // @[NV_NVDLA_csc.scala 142:20:@23713.4]
  assign io_sc2mac_wt_a_bits_data_9 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_9; // @[NV_NVDLA_csc.scala 142:20:@23714.4]
  assign io_sc2mac_wt_a_bits_data_10 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_10; // @[NV_NVDLA_csc.scala 142:20:@23715.4]
  assign io_sc2mac_wt_a_bits_data_11 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_11; // @[NV_NVDLA_csc.scala 142:20:@23716.4]
  assign io_sc2mac_wt_a_bits_data_12 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_12; // @[NV_NVDLA_csc.scala 142:20:@23717.4]
  assign io_sc2mac_wt_a_bits_data_13 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_13; // @[NV_NVDLA_csc.scala 142:20:@23718.4]
  assign io_sc2mac_wt_a_bits_data_14 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_14; // @[NV_NVDLA_csc.scala 142:20:@23719.4]
  assign io_sc2mac_wt_a_bits_data_15 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_15; // @[NV_NVDLA_csc.scala 142:20:@23720.4]
  assign io_sc2mac_wt_a_bits_data_16 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_16; // @[NV_NVDLA_csc.scala 142:20:@23721.4]
  assign io_sc2mac_wt_a_bits_data_17 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_17; // @[NV_NVDLA_csc.scala 142:20:@23722.4]
  assign io_sc2mac_wt_a_bits_data_18 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_18; // @[NV_NVDLA_csc.scala 142:20:@23723.4]
  assign io_sc2mac_wt_a_bits_data_19 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_19; // @[NV_NVDLA_csc.scala 142:20:@23724.4]
  assign io_sc2mac_wt_a_bits_data_20 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_20; // @[NV_NVDLA_csc.scala 142:20:@23725.4]
  assign io_sc2mac_wt_a_bits_data_21 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_21; // @[NV_NVDLA_csc.scala 142:20:@23726.4]
  assign io_sc2mac_wt_a_bits_data_22 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_22; // @[NV_NVDLA_csc.scala 142:20:@23727.4]
  assign io_sc2mac_wt_a_bits_data_23 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_23; // @[NV_NVDLA_csc.scala 142:20:@23728.4]
  assign io_sc2mac_wt_a_bits_data_24 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_24; // @[NV_NVDLA_csc.scala 142:20:@23729.4]
  assign io_sc2mac_wt_a_bits_data_25 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_25; // @[NV_NVDLA_csc.scala 142:20:@23730.4]
  assign io_sc2mac_wt_a_bits_data_26 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_26; // @[NV_NVDLA_csc.scala 142:20:@23731.4]
  assign io_sc2mac_wt_a_bits_data_27 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_27; // @[NV_NVDLA_csc.scala 142:20:@23732.4]
  assign io_sc2mac_wt_a_bits_data_28 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_28; // @[NV_NVDLA_csc.scala 142:20:@23733.4]
  assign io_sc2mac_wt_a_bits_data_29 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_29; // @[NV_NVDLA_csc.scala 142:20:@23734.4]
  assign io_sc2mac_wt_a_bits_data_30 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_30; // @[NV_NVDLA_csc.scala 142:20:@23735.4]
  assign io_sc2mac_wt_a_bits_data_31 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_31; // @[NV_NVDLA_csc.scala 142:20:@23736.4]
  assign io_sc2mac_wt_a_bits_data_32 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_32; // @[NV_NVDLA_csc.scala 142:20:@23737.4]
  assign io_sc2mac_wt_a_bits_data_33 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_33; // @[NV_NVDLA_csc.scala 142:20:@23738.4]
  assign io_sc2mac_wt_a_bits_data_34 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_34; // @[NV_NVDLA_csc.scala 142:20:@23739.4]
  assign io_sc2mac_wt_a_bits_data_35 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_35; // @[NV_NVDLA_csc.scala 142:20:@23740.4]
  assign io_sc2mac_wt_a_bits_data_36 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_36; // @[NV_NVDLA_csc.scala 142:20:@23741.4]
  assign io_sc2mac_wt_a_bits_data_37 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_37; // @[NV_NVDLA_csc.scala 142:20:@23742.4]
  assign io_sc2mac_wt_a_bits_data_38 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_38; // @[NV_NVDLA_csc.scala 142:20:@23743.4]
  assign io_sc2mac_wt_a_bits_data_39 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_39; // @[NV_NVDLA_csc.scala 142:20:@23744.4]
  assign io_sc2mac_wt_a_bits_data_40 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_40; // @[NV_NVDLA_csc.scala 142:20:@23745.4]
  assign io_sc2mac_wt_a_bits_data_41 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_41; // @[NV_NVDLA_csc.scala 142:20:@23746.4]
  assign io_sc2mac_wt_a_bits_data_42 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_42; // @[NV_NVDLA_csc.scala 142:20:@23747.4]
  assign io_sc2mac_wt_a_bits_data_43 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_43; // @[NV_NVDLA_csc.scala 142:20:@23748.4]
  assign io_sc2mac_wt_a_bits_data_44 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_44; // @[NV_NVDLA_csc.scala 142:20:@23749.4]
  assign io_sc2mac_wt_a_bits_data_45 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_45; // @[NV_NVDLA_csc.scala 142:20:@23750.4]
  assign io_sc2mac_wt_a_bits_data_46 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_46; // @[NV_NVDLA_csc.scala 142:20:@23751.4]
  assign io_sc2mac_wt_a_bits_data_47 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_47; // @[NV_NVDLA_csc.scala 142:20:@23752.4]
  assign io_sc2mac_wt_a_bits_data_48 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_48; // @[NV_NVDLA_csc.scala 142:20:@23753.4]
  assign io_sc2mac_wt_a_bits_data_49 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_49; // @[NV_NVDLA_csc.scala 142:20:@23754.4]
  assign io_sc2mac_wt_a_bits_data_50 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_50; // @[NV_NVDLA_csc.scala 142:20:@23755.4]
  assign io_sc2mac_wt_a_bits_data_51 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_51; // @[NV_NVDLA_csc.scala 142:20:@23756.4]
  assign io_sc2mac_wt_a_bits_data_52 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_52; // @[NV_NVDLA_csc.scala 142:20:@23757.4]
  assign io_sc2mac_wt_a_bits_data_53 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_53; // @[NV_NVDLA_csc.scala 142:20:@23758.4]
  assign io_sc2mac_wt_a_bits_data_54 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_54; // @[NV_NVDLA_csc.scala 142:20:@23759.4]
  assign io_sc2mac_wt_a_bits_data_55 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_55; // @[NV_NVDLA_csc.scala 142:20:@23760.4]
  assign io_sc2mac_wt_a_bits_data_56 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_56; // @[NV_NVDLA_csc.scala 142:20:@23761.4]
  assign io_sc2mac_wt_a_bits_data_57 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_57; // @[NV_NVDLA_csc.scala 142:20:@23762.4]
  assign io_sc2mac_wt_a_bits_data_58 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_58; // @[NV_NVDLA_csc.scala 142:20:@23763.4]
  assign io_sc2mac_wt_a_bits_data_59 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_59; // @[NV_NVDLA_csc.scala 142:20:@23764.4]
  assign io_sc2mac_wt_a_bits_data_60 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_60; // @[NV_NVDLA_csc.scala 142:20:@23765.4]
  assign io_sc2mac_wt_a_bits_data_61 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_61; // @[NV_NVDLA_csc.scala 142:20:@23766.4]
  assign io_sc2mac_wt_a_bits_data_62 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_62; // @[NV_NVDLA_csc.scala 142:20:@23767.4]
  assign io_sc2mac_wt_a_bits_data_63 = NV_NVDLA_CSC_wl_io_sc2mac_wt_a_bits_data_63; // @[NV_NVDLA_csc.scala 142:20:@23768.4]
  assign io_sc2mac_wt_b_valid = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_valid; // @[NV_NVDLA_csc.scala 143:20:@23994.4]
  assign io_sc2mac_wt_b_bits_sel_0 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_0; // @[NV_NVDLA_csc.scala 143:20:@23978.4]
  assign io_sc2mac_wt_b_bits_sel_1 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_1; // @[NV_NVDLA_csc.scala 143:20:@23979.4]
  assign io_sc2mac_wt_b_bits_sel_2 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_2; // @[NV_NVDLA_csc.scala 143:20:@23980.4]
  assign io_sc2mac_wt_b_bits_sel_3 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_3; // @[NV_NVDLA_csc.scala 143:20:@23981.4]
  assign io_sc2mac_wt_b_bits_sel_4 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_4; // @[NV_NVDLA_csc.scala 143:20:@23982.4]
  assign io_sc2mac_wt_b_bits_sel_5 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_5; // @[NV_NVDLA_csc.scala 143:20:@23983.4]
  assign io_sc2mac_wt_b_bits_sel_6 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_6; // @[NV_NVDLA_csc.scala 143:20:@23984.4]
  assign io_sc2mac_wt_b_bits_sel_7 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_7; // @[NV_NVDLA_csc.scala 143:20:@23985.4]
  assign io_sc2mac_wt_b_bits_sel_8 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_8; // @[NV_NVDLA_csc.scala 143:20:@23986.4]
  assign io_sc2mac_wt_b_bits_sel_9 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_9; // @[NV_NVDLA_csc.scala 143:20:@23987.4]
  assign io_sc2mac_wt_b_bits_sel_10 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_10; // @[NV_NVDLA_csc.scala 143:20:@23988.4]
  assign io_sc2mac_wt_b_bits_sel_11 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_11; // @[NV_NVDLA_csc.scala 143:20:@23989.4]
  assign io_sc2mac_wt_b_bits_sel_12 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_12; // @[NV_NVDLA_csc.scala 143:20:@23990.4]
  assign io_sc2mac_wt_b_bits_sel_13 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_13; // @[NV_NVDLA_csc.scala 143:20:@23991.4]
  assign io_sc2mac_wt_b_bits_sel_14 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_14; // @[NV_NVDLA_csc.scala 143:20:@23992.4]
  assign io_sc2mac_wt_b_bits_sel_15 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_sel_15; // @[NV_NVDLA_csc.scala 143:20:@23993.4]
  assign io_sc2mac_wt_b_bits_mask_0 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_0; // @[NV_NVDLA_csc.scala 143:20:@23914.4]
  assign io_sc2mac_wt_b_bits_mask_1 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_1; // @[NV_NVDLA_csc.scala 143:20:@23915.4]
  assign io_sc2mac_wt_b_bits_mask_2 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_2; // @[NV_NVDLA_csc.scala 143:20:@23916.4]
  assign io_sc2mac_wt_b_bits_mask_3 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_3; // @[NV_NVDLA_csc.scala 143:20:@23917.4]
  assign io_sc2mac_wt_b_bits_mask_4 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_4; // @[NV_NVDLA_csc.scala 143:20:@23918.4]
  assign io_sc2mac_wt_b_bits_mask_5 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_5; // @[NV_NVDLA_csc.scala 143:20:@23919.4]
  assign io_sc2mac_wt_b_bits_mask_6 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_6; // @[NV_NVDLA_csc.scala 143:20:@23920.4]
  assign io_sc2mac_wt_b_bits_mask_7 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_7; // @[NV_NVDLA_csc.scala 143:20:@23921.4]
  assign io_sc2mac_wt_b_bits_mask_8 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_8; // @[NV_NVDLA_csc.scala 143:20:@23922.4]
  assign io_sc2mac_wt_b_bits_mask_9 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_9; // @[NV_NVDLA_csc.scala 143:20:@23923.4]
  assign io_sc2mac_wt_b_bits_mask_10 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_10; // @[NV_NVDLA_csc.scala 143:20:@23924.4]
  assign io_sc2mac_wt_b_bits_mask_11 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_11; // @[NV_NVDLA_csc.scala 143:20:@23925.4]
  assign io_sc2mac_wt_b_bits_mask_12 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_12; // @[NV_NVDLA_csc.scala 143:20:@23926.4]
  assign io_sc2mac_wt_b_bits_mask_13 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_13; // @[NV_NVDLA_csc.scala 143:20:@23927.4]
  assign io_sc2mac_wt_b_bits_mask_14 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_14; // @[NV_NVDLA_csc.scala 143:20:@23928.4]
  assign io_sc2mac_wt_b_bits_mask_15 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_15; // @[NV_NVDLA_csc.scala 143:20:@23929.4]
  assign io_sc2mac_wt_b_bits_mask_16 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_16; // @[NV_NVDLA_csc.scala 143:20:@23930.4]
  assign io_sc2mac_wt_b_bits_mask_17 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_17; // @[NV_NVDLA_csc.scala 143:20:@23931.4]
  assign io_sc2mac_wt_b_bits_mask_18 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_18; // @[NV_NVDLA_csc.scala 143:20:@23932.4]
  assign io_sc2mac_wt_b_bits_mask_19 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_19; // @[NV_NVDLA_csc.scala 143:20:@23933.4]
  assign io_sc2mac_wt_b_bits_mask_20 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_20; // @[NV_NVDLA_csc.scala 143:20:@23934.4]
  assign io_sc2mac_wt_b_bits_mask_21 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_21; // @[NV_NVDLA_csc.scala 143:20:@23935.4]
  assign io_sc2mac_wt_b_bits_mask_22 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_22; // @[NV_NVDLA_csc.scala 143:20:@23936.4]
  assign io_sc2mac_wt_b_bits_mask_23 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_23; // @[NV_NVDLA_csc.scala 143:20:@23937.4]
  assign io_sc2mac_wt_b_bits_mask_24 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_24; // @[NV_NVDLA_csc.scala 143:20:@23938.4]
  assign io_sc2mac_wt_b_bits_mask_25 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_25; // @[NV_NVDLA_csc.scala 143:20:@23939.4]
  assign io_sc2mac_wt_b_bits_mask_26 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_26; // @[NV_NVDLA_csc.scala 143:20:@23940.4]
  assign io_sc2mac_wt_b_bits_mask_27 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_27; // @[NV_NVDLA_csc.scala 143:20:@23941.4]
  assign io_sc2mac_wt_b_bits_mask_28 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_28; // @[NV_NVDLA_csc.scala 143:20:@23942.4]
  assign io_sc2mac_wt_b_bits_mask_29 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_29; // @[NV_NVDLA_csc.scala 143:20:@23943.4]
  assign io_sc2mac_wt_b_bits_mask_30 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_30; // @[NV_NVDLA_csc.scala 143:20:@23944.4]
  assign io_sc2mac_wt_b_bits_mask_31 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_31; // @[NV_NVDLA_csc.scala 143:20:@23945.4]
  assign io_sc2mac_wt_b_bits_mask_32 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_32; // @[NV_NVDLA_csc.scala 143:20:@23946.4]
  assign io_sc2mac_wt_b_bits_mask_33 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_33; // @[NV_NVDLA_csc.scala 143:20:@23947.4]
  assign io_sc2mac_wt_b_bits_mask_34 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_34; // @[NV_NVDLA_csc.scala 143:20:@23948.4]
  assign io_sc2mac_wt_b_bits_mask_35 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_35; // @[NV_NVDLA_csc.scala 143:20:@23949.4]
  assign io_sc2mac_wt_b_bits_mask_36 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_36; // @[NV_NVDLA_csc.scala 143:20:@23950.4]
  assign io_sc2mac_wt_b_bits_mask_37 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_37; // @[NV_NVDLA_csc.scala 143:20:@23951.4]
  assign io_sc2mac_wt_b_bits_mask_38 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_38; // @[NV_NVDLA_csc.scala 143:20:@23952.4]
  assign io_sc2mac_wt_b_bits_mask_39 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_39; // @[NV_NVDLA_csc.scala 143:20:@23953.4]
  assign io_sc2mac_wt_b_bits_mask_40 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_40; // @[NV_NVDLA_csc.scala 143:20:@23954.4]
  assign io_sc2mac_wt_b_bits_mask_41 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_41; // @[NV_NVDLA_csc.scala 143:20:@23955.4]
  assign io_sc2mac_wt_b_bits_mask_42 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_42; // @[NV_NVDLA_csc.scala 143:20:@23956.4]
  assign io_sc2mac_wt_b_bits_mask_43 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_43; // @[NV_NVDLA_csc.scala 143:20:@23957.4]
  assign io_sc2mac_wt_b_bits_mask_44 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_44; // @[NV_NVDLA_csc.scala 143:20:@23958.4]
  assign io_sc2mac_wt_b_bits_mask_45 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_45; // @[NV_NVDLA_csc.scala 143:20:@23959.4]
  assign io_sc2mac_wt_b_bits_mask_46 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_46; // @[NV_NVDLA_csc.scala 143:20:@23960.4]
  assign io_sc2mac_wt_b_bits_mask_47 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_47; // @[NV_NVDLA_csc.scala 143:20:@23961.4]
  assign io_sc2mac_wt_b_bits_mask_48 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_48; // @[NV_NVDLA_csc.scala 143:20:@23962.4]
  assign io_sc2mac_wt_b_bits_mask_49 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_49; // @[NV_NVDLA_csc.scala 143:20:@23963.4]
  assign io_sc2mac_wt_b_bits_mask_50 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_50; // @[NV_NVDLA_csc.scala 143:20:@23964.4]
  assign io_sc2mac_wt_b_bits_mask_51 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_51; // @[NV_NVDLA_csc.scala 143:20:@23965.4]
  assign io_sc2mac_wt_b_bits_mask_52 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_52; // @[NV_NVDLA_csc.scala 143:20:@23966.4]
  assign io_sc2mac_wt_b_bits_mask_53 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_53; // @[NV_NVDLA_csc.scala 143:20:@23967.4]
  assign io_sc2mac_wt_b_bits_mask_54 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_54; // @[NV_NVDLA_csc.scala 143:20:@23968.4]
  assign io_sc2mac_wt_b_bits_mask_55 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_55; // @[NV_NVDLA_csc.scala 143:20:@23969.4]
  assign io_sc2mac_wt_b_bits_mask_56 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_56; // @[NV_NVDLA_csc.scala 143:20:@23970.4]
  assign io_sc2mac_wt_b_bits_mask_57 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_57; // @[NV_NVDLA_csc.scala 143:20:@23971.4]
  assign io_sc2mac_wt_b_bits_mask_58 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_58; // @[NV_NVDLA_csc.scala 143:20:@23972.4]
  assign io_sc2mac_wt_b_bits_mask_59 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_59; // @[NV_NVDLA_csc.scala 143:20:@23973.4]
  assign io_sc2mac_wt_b_bits_mask_60 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_60; // @[NV_NVDLA_csc.scala 143:20:@23974.4]
  assign io_sc2mac_wt_b_bits_mask_61 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_61; // @[NV_NVDLA_csc.scala 143:20:@23975.4]
  assign io_sc2mac_wt_b_bits_mask_62 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_62; // @[NV_NVDLA_csc.scala 143:20:@23976.4]
  assign io_sc2mac_wt_b_bits_mask_63 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_mask_63; // @[NV_NVDLA_csc.scala 143:20:@23977.4]
  assign io_sc2mac_wt_b_bits_data_0 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_0; // @[NV_NVDLA_csc.scala 143:20:@23850.4]
  assign io_sc2mac_wt_b_bits_data_1 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_1; // @[NV_NVDLA_csc.scala 143:20:@23851.4]
  assign io_sc2mac_wt_b_bits_data_2 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_2; // @[NV_NVDLA_csc.scala 143:20:@23852.4]
  assign io_sc2mac_wt_b_bits_data_3 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_3; // @[NV_NVDLA_csc.scala 143:20:@23853.4]
  assign io_sc2mac_wt_b_bits_data_4 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_4; // @[NV_NVDLA_csc.scala 143:20:@23854.4]
  assign io_sc2mac_wt_b_bits_data_5 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_5; // @[NV_NVDLA_csc.scala 143:20:@23855.4]
  assign io_sc2mac_wt_b_bits_data_6 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_6; // @[NV_NVDLA_csc.scala 143:20:@23856.4]
  assign io_sc2mac_wt_b_bits_data_7 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_7; // @[NV_NVDLA_csc.scala 143:20:@23857.4]
  assign io_sc2mac_wt_b_bits_data_8 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_8; // @[NV_NVDLA_csc.scala 143:20:@23858.4]
  assign io_sc2mac_wt_b_bits_data_9 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_9; // @[NV_NVDLA_csc.scala 143:20:@23859.4]
  assign io_sc2mac_wt_b_bits_data_10 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_10; // @[NV_NVDLA_csc.scala 143:20:@23860.4]
  assign io_sc2mac_wt_b_bits_data_11 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_11; // @[NV_NVDLA_csc.scala 143:20:@23861.4]
  assign io_sc2mac_wt_b_bits_data_12 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_12; // @[NV_NVDLA_csc.scala 143:20:@23862.4]
  assign io_sc2mac_wt_b_bits_data_13 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_13; // @[NV_NVDLA_csc.scala 143:20:@23863.4]
  assign io_sc2mac_wt_b_bits_data_14 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_14; // @[NV_NVDLA_csc.scala 143:20:@23864.4]
  assign io_sc2mac_wt_b_bits_data_15 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_15; // @[NV_NVDLA_csc.scala 143:20:@23865.4]
  assign io_sc2mac_wt_b_bits_data_16 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_16; // @[NV_NVDLA_csc.scala 143:20:@23866.4]
  assign io_sc2mac_wt_b_bits_data_17 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_17; // @[NV_NVDLA_csc.scala 143:20:@23867.4]
  assign io_sc2mac_wt_b_bits_data_18 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_18; // @[NV_NVDLA_csc.scala 143:20:@23868.4]
  assign io_sc2mac_wt_b_bits_data_19 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_19; // @[NV_NVDLA_csc.scala 143:20:@23869.4]
  assign io_sc2mac_wt_b_bits_data_20 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_20; // @[NV_NVDLA_csc.scala 143:20:@23870.4]
  assign io_sc2mac_wt_b_bits_data_21 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_21; // @[NV_NVDLA_csc.scala 143:20:@23871.4]
  assign io_sc2mac_wt_b_bits_data_22 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_22; // @[NV_NVDLA_csc.scala 143:20:@23872.4]
  assign io_sc2mac_wt_b_bits_data_23 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_23; // @[NV_NVDLA_csc.scala 143:20:@23873.4]
  assign io_sc2mac_wt_b_bits_data_24 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_24; // @[NV_NVDLA_csc.scala 143:20:@23874.4]
  assign io_sc2mac_wt_b_bits_data_25 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_25; // @[NV_NVDLA_csc.scala 143:20:@23875.4]
  assign io_sc2mac_wt_b_bits_data_26 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_26; // @[NV_NVDLA_csc.scala 143:20:@23876.4]
  assign io_sc2mac_wt_b_bits_data_27 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_27; // @[NV_NVDLA_csc.scala 143:20:@23877.4]
  assign io_sc2mac_wt_b_bits_data_28 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_28; // @[NV_NVDLA_csc.scala 143:20:@23878.4]
  assign io_sc2mac_wt_b_bits_data_29 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_29; // @[NV_NVDLA_csc.scala 143:20:@23879.4]
  assign io_sc2mac_wt_b_bits_data_30 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_30; // @[NV_NVDLA_csc.scala 143:20:@23880.4]
  assign io_sc2mac_wt_b_bits_data_31 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_31; // @[NV_NVDLA_csc.scala 143:20:@23881.4]
  assign io_sc2mac_wt_b_bits_data_32 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_32; // @[NV_NVDLA_csc.scala 143:20:@23882.4]
  assign io_sc2mac_wt_b_bits_data_33 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_33; // @[NV_NVDLA_csc.scala 143:20:@23883.4]
  assign io_sc2mac_wt_b_bits_data_34 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_34; // @[NV_NVDLA_csc.scala 143:20:@23884.4]
  assign io_sc2mac_wt_b_bits_data_35 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_35; // @[NV_NVDLA_csc.scala 143:20:@23885.4]
  assign io_sc2mac_wt_b_bits_data_36 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_36; // @[NV_NVDLA_csc.scala 143:20:@23886.4]
  assign io_sc2mac_wt_b_bits_data_37 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_37; // @[NV_NVDLA_csc.scala 143:20:@23887.4]
  assign io_sc2mac_wt_b_bits_data_38 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_38; // @[NV_NVDLA_csc.scala 143:20:@23888.4]
  assign io_sc2mac_wt_b_bits_data_39 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_39; // @[NV_NVDLA_csc.scala 143:20:@23889.4]
  assign io_sc2mac_wt_b_bits_data_40 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_40; // @[NV_NVDLA_csc.scala 143:20:@23890.4]
  assign io_sc2mac_wt_b_bits_data_41 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_41; // @[NV_NVDLA_csc.scala 143:20:@23891.4]
  assign io_sc2mac_wt_b_bits_data_42 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_42; // @[NV_NVDLA_csc.scala 143:20:@23892.4]
  assign io_sc2mac_wt_b_bits_data_43 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_43; // @[NV_NVDLA_csc.scala 143:20:@23893.4]
  assign io_sc2mac_wt_b_bits_data_44 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_44; // @[NV_NVDLA_csc.scala 143:20:@23894.4]
  assign io_sc2mac_wt_b_bits_data_45 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_45; // @[NV_NVDLA_csc.scala 143:20:@23895.4]
  assign io_sc2mac_wt_b_bits_data_46 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_46; // @[NV_NVDLA_csc.scala 143:20:@23896.4]
  assign io_sc2mac_wt_b_bits_data_47 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_47; // @[NV_NVDLA_csc.scala 143:20:@23897.4]
  assign io_sc2mac_wt_b_bits_data_48 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_48; // @[NV_NVDLA_csc.scala 143:20:@23898.4]
  assign io_sc2mac_wt_b_bits_data_49 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_49; // @[NV_NVDLA_csc.scala 143:20:@23899.4]
  assign io_sc2mac_wt_b_bits_data_50 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_50; // @[NV_NVDLA_csc.scala 143:20:@23900.4]
  assign io_sc2mac_wt_b_bits_data_51 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_51; // @[NV_NVDLA_csc.scala 143:20:@23901.4]
  assign io_sc2mac_wt_b_bits_data_52 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_52; // @[NV_NVDLA_csc.scala 143:20:@23902.4]
  assign io_sc2mac_wt_b_bits_data_53 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_53; // @[NV_NVDLA_csc.scala 143:20:@23903.4]
  assign io_sc2mac_wt_b_bits_data_54 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_54; // @[NV_NVDLA_csc.scala 143:20:@23904.4]
  assign io_sc2mac_wt_b_bits_data_55 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_55; // @[NV_NVDLA_csc.scala 143:20:@23905.4]
  assign io_sc2mac_wt_b_bits_data_56 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_56; // @[NV_NVDLA_csc.scala 143:20:@23906.4]
  assign io_sc2mac_wt_b_bits_data_57 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_57; // @[NV_NVDLA_csc.scala 143:20:@23907.4]
  assign io_sc2mac_wt_b_bits_data_58 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_58; // @[NV_NVDLA_csc.scala 143:20:@23908.4]
  assign io_sc2mac_wt_b_bits_data_59 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_59; // @[NV_NVDLA_csc.scala 143:20:@23909.4]
  assign io_sc2mac_wt_b_bits_data_60 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_60; // @[NV_NVDLA_csc.scala 143:20:@23910.4]
  assign io_sc2mac_wt_b_bits_data_61 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_61; // @[NV_NVDLA_csc.scala 143:20:@23911.4]
  assign io_sc2mac_wt_b_bits_data_62 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_62; // @[NV_NVDLA_csc.scala 143:20:@23912.4]
  assign io_sc2mac_wt_b_bits_data_63 = NV_NVDLA_CSC_wl_io_sc2mac_wt_b_bits_data_63; // @[NV_NVDLA_csc.scala 143:20:@23913.4]
  assign NV_NVDLA_CSC_regfile_reset = io_nvdla_core_rstn == 1'h0; // @[:@23634.4]
  assign NV_NVDLA_CSC_regfile_io_nvdla_core_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_csc.scala 79:33:@23638.4]
  assign NV_NVDLA_CSC_regfile_io_csb2csc_req_valid = io_csb2csc_req_valid; // @[NV_NVDLA_csc.scala 80:26:@23642.4]
  assign NV_NVDLA_CSC_regfile_io_csb2csc_req_bits = io_csb2csc_req_bits; // @[NV_NVDLA_csc.scala 80:26:@23641.4]
  assign NV_NVDLA_CSC_regfile_io_dp2reg_done = NV_NVDLA_CSC_sg_io_dp2reg_done; // @[NV_NVDLA_csc.scala 82:30:@23644.4]
  assign NV_NVDLA_CSC_sg_reset = io_nvdla_core_rstn == 1'h0; // @[:@23637.4]
  assign NV_NVDLA_CSC_sg_io_nvdla_core_clk = NV_NVDLA_slcg_io_nvdla_core_gated_clk; // @[NV_NVDLA_csc.scala 90:28:@23646.4]
  assign NV_NVDLA_CSC_sg_io_nvdla_core_ng_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_csc.scala 89:31:@23645.4]
  assign NV_NVDLA_CSC_sg_io_cdma2sc_dat_updt_valid = io_cdma2sc_dat_updt_valid; // @[NV_NVDLA_csc.scala 93:30:@23650.4]
  assign NV_NVDLA_CSC_sg_io_cdma2sc_dat_updt_bits_slices = io_cdma2sc_dat_updt_bits_slices; // @[NV_NVDLA_csc.scala 93:30:@23648.4]
  assign NV_NVDLA_CSC_sg_io_cdma2sc_dat_pending_ack = io_cdma2sc_dat_pending_ack; // @[NV_NVDLA_csc.scala 96:37:@23656.4]
  assign NV_NVDLA_CSC_sg_io_cdma2sc_wt_updt_valid = io_cdma2sc_wt_updt_valid; // @[NV_NVDLA_csc.scala 94:29:@23653.4]
  assign NV_NVDLA_CSC_sg_io_cdma2sc_wt_updt_bits_kernels = io_cdma2sc_wt_updt_bits_kernels; // @[NV_NVDLA_csc.scala 94:29:@23651.4]
  assign NV_NVDLA_CSC_sg_io_cdma2sc_wt_pending_ack = io_cdma2sc_wt_pending_ack; // @[NV_NVDLA_csc.scala 97:36:@23657.4]
  assign NV_NVDLA_CSC_sg_io_accu2sc_credit_size_valid = io_accu2sc_credit_size_valid; // @[NV_NVDLA_csc.scala 95:33:@23655.4]
  assign NV_NVDLA_CSC_sg_io_accu2sc_credit_size_bits = io_accu2sc_credit_size_bits; // @[NV_NVDLA_csc.scala 95:33:@23654.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_op_en = NV_NVDLA_CSC_regfile_io_reg2dp_op_en; // @[NV_NVDLA_csc.scala 101:26:@23660.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_conv_mode = NV_NVDLA_CSC_regfile_io_reg2dp_field_conv_mode; // @[NV_NVDLA_csc.scala 102:30:@23661.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_data_reuse = NV_NVDLA_CSC_regfile_io_reg2dp_field_data_reuse; // @[NV_NVDLA_csc.scala 104:31:@23663.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_skip_data_rls = NV_NVDLA_CSC_regfile_io_reg2dp_field_skip_data_rls; // @[NV_NVDLA_csc.scala 105:34:@23664.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_weight_reuse = NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_reuse; // @[NV_NVDLA_csc.scala 106:33:@23665.4 NV_NVDLA_csc.scala 108:33:@23667.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_skip_weight_rls = NV_NVDLA_CSC_regfile_io_reg2dp_field_skip_weight_rls; // @[NV_NVDLA_csc.scala 107:36:@23666.4 NV_NVDLA_csc.scala 109:36:@23668.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_datain_format = NV_NVDLA_CSC_regfile_io_reg2dp_field_datain_format; // @[NV_NVDLA_csc.scala 111:34:@23670.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_datain_height_ext = NV_NVDLA_CSC_regfile_io_reg2dp_field_datain_height_ext; // @[NV_NVDLA_csc.scala 112:38:@23671.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_y_extension = NV_NVDLA_CSC_regfile_io_reg2dp_field_y_extension; // @[NV_NVDLA_csc.scala 113:32:@23672.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_weight_width_ext = NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_width_ext; // @[NV_NVDLA_csc.scala 114:37:@23673.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_weight_height_ext = NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_height_ext; // @[NV_NVDLA_csc.scala 115:38:@23674.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_weight_channel_ext = NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_channel_ext; // @[NV_NVDLA_csc.scala 116:39:@23675.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_weight_kernel = NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_kernel; // @[NV_NVDLA_csc.scala 117:34:@23676.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_dataout_width = NV_NVDLA_CSC_regfile_io_reg2dp_field_dataout_width; // @[NV_NVDLA_csc.scala 118:34:@23677.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_dataout_height = NV_NVDLA_CSC_regfile_io_reg2dp_field_dataout_height; // @[NV_NVDLA_csc.scala 119:35:@23678.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_data_bank = NV_NVDLA_CSC_regfile_io_reg2dp_field_data_bank; // @[NV_NVDLA_csc.scala 120:30:@23679.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_weight_bank = NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_bank; // @[NV_NVDLA_csc.scala 121:32:@23680.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_atomics = NV_NVDLA_CSC_regfile_io_reg2dp_field_atomics; // @[NV_NVDLA_csc.scala 122:28:@23681.4]
  assign NV_NVDLA_CSC_sg_io_reg2dp_rls_slices = NV_NVDLA_CSC_regfile_io_reg2dp_field_rls_slices; // @[NV_NVDLA_csc.scala 123:31:@23682.4]
  assign NV_NVDLA_CSC_wl_reset = io_nvdla_core_rstn == 1'h0; // @[:@23685.4]
  assign NV_NVDLA_CSC_wl_io_nvdla_core_clk = NV_NVDLA_slcg_1_io_nvdla_core_gated_clk; // @[NV_NVDLA_csc.scala 132:28:@23687.4]
  assign NV_NVDLA_CSC_wl_io_nvdla_core_ng_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_csc.scala 131:31:@23686.4]
  assign NV_NVDLA_CSC_wl_io_sg2wl_pd_valid = NV_NVDLA_CSC_sg_io_sg2wl_pd_valid; // @[NV_NVDLA_csc.scala 134:19:@23690.4]
  assign NV_NVDLA_CSC_wl_io_sg2wl_pd_bits = NV_NVDLA_CSC_sg_io_sg2wl_pd_bits; // @[NV_NVDLA_csc.scala 134:19:@23689.4]
  assign NV_NVDLA_CSC_wl_io_sg2wl_reuse_rls = NV_NVDLA_CSC_sg_io_sg2wl_reuse_rls; // @[NV_NVDLA_csc.scala 134:19:@23688.4]
  assign NV_NVDLA_CSC_wl_io_sc_state = NV_NVDLA_CSC_sg_io_sc_state; // @[NV_NVDLA_csc.scala 135:22:@23691.4]
  assign NV_NVDLA_CSC_wl_io_sc2cdma_wt_pending_req = io_sc2cdma_wt_pending_req; // @[NV_NVDLA_csc.scala 136:36:@23692.4]
  assign NV_NVDLA_CSC_wl_io_sc2buf_wt_rd_data_valid = io_sc2buf_wt_rd_data_valid; // @[NV_NVDLA_csc.scala 139:21:@23700.4]
  assign NV_NVDLA_CSC_wl_io_sc2buf_wt_rd_data_bits = io_sc2buf_wt_rd_data_bits; // @[NV_NVDLA_csc.scala 139:21:@23699.4]
  assign NV_NVDLA_CSC_wl_io_reg2dp_op_en = NV_NVDLA_CSC_regfile_io_reg2dp_op_en; // @[NV_NVDLA_csc.scala 145:26:@23995.4]
  assign NV_NVDLA_CSC_wl_io_reg2dp_y_extension = NV_NVDLA_CSC_regfile_io_reg2dp_field_y_extension; // @[NV_NVDLA_csc.scala 148:32:@23998.4]
  assign NV_NVDLA_CSC_wl_io_reg2dp_skip_weight_rls = NV_NVDLA_CSC_regfile_io_reg2dp_field_skip_weight_rls; // @[NV_NVDLA_csc.scala 150:36:@24000.4]
  assign NV_NVDLA_CSC_wl_io_reg2dp_weight_format = NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_format; // @[NV_NVDLA_csc.scala 151:34:@24001.4]
  assign NV_NVDLA_CSC_wl_io_reg2dp_weight_bytes = NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_bytes; // @[NV_NVDLA_csc.scala 152:33:@24002.4]
  assign NV_NVDLA_CSC_wl_io_reg2dp_wmb_bytes = NV_NVDLA_CSC_regfile_io_reg2dp_field_wmb_bytes; // @[NV_NVDLA_csc.scala 153:30:@24003.4]
  assign NV_NVDLA_CSC_wl_io_reg2dp_data_bank = NV_NVDLA_CSC_regfile_io_reg2dp_field_data_bank; // @[NV_NVDLA_csc.scala 154:30:@24004.4]
  assign NV_NVDLA_CSC_wl_io_reg2dp_weight_bank = NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_bank; // @[NV_NVDLA_csc.scala 155:32:@24005.4]
  assign NV_NVDLA_CSC_dl_reset = io_nvdla_core_rstn == 1'h0; // @[:@24008.4]
  assign NV_NVDLA_CSC_dl_io_nvdla_core_clk = NV_NVDLA_slcg_2_io_nvdla_core_gated_clk; // @[NV_NVDLA_csc.scala 164:28:@24010.4]
  assign NV_NVDLA_CSC_dl_io_nvdla_core_ng_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_csc.scala 163:31:@24009.4]
  assign NV_NVDLA_CSC_dl_io_sc_state = NV_NVDLA_CSC_sg_io_sc_state; // @[NV_NVDLA_csc.scala 166:22:@24014.4]
  assign NV_NVDLA_CSC_dl_io_sg2dl_pd_valid = NV_NVDLA_CSC_sg_io_sg2dl_pd_valid; // @[NV_NVDLA_csc.scala 165:19:@24013.4]
  assign NV_NVDLA_CSC_dl_io_sg2dl_reuse_rls = NV_NVDLA_CSC_sg_io_sg2dl_reuse_rls; // @[NV_NVDLA_csc.scala 165:19:@24011.4]
  assign NV_NVDLA_CSC_dl_io_sc2cdma_dat_pending_req = io_sc2cdma_dat_pending_req; // @[NV_NVDLA_csc.scala 167:37:@24015.4]
  assign NV_NVDLA_CSC_dl_io_sc2buf_dat_rd_data_valid = io_sc2buf_dat_rd_data_valid; // @[NV_NVDLA_csc.scala 170:22:@24023.4]
  assign NV_NVDLA_CSC_dl_io_sc2buf_dat_rd_data_bits = io_sc2buf_dat_rd_data_bits; // @[NV_NVDLA_csc.scala 170:22:@24022.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_op_en = NV_NVDLA_CSC_regfile_io_reg2dp_op_en; // @[NV_NVDLA_csc.scala 174:26:@24286.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_conv_mode = NV_NVDLA_CSC_regfile_io_reg2dp_field_conv_mode; // @[NV_NVDLA_csc.scala 175:30:@24287.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_datain_format = NV_NVDLA_CSC_regfile_io_reg2dp_field_datain_format; // @[NV_NVDLA_csc.scala 178:34:@24290.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_skip_data_rls = NV_NVDLA_CSC_regfile_io_reg2dp_field_skip_data_rls; // @[NV_NVDLA_csc.scala 179:34:@24291.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_datain_channel_ext = NV_NVDLA_CSC_regfile_io_reg2dp_field_datain_channel_ext; // @[NV_NVDLA_csc.scala 180:39:@24292.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_datain_height_ext = NV_NVDLA_CSC_regfile_io_reg2dp_field_datain_height_ext; // @[NV_NVDLA_csc.scala 181:38:@24293.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_datain_width_ext = NV_NVDLA_CSC_regfile_io_reg2dp_field_datain_width_ext; // @[NV_NVDLA_csc.scala 182:37:@24294.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_y_extension = NV_NVDLA_CSC_regfile_io_reg2dp_field_y_extension; // @[NV_NVDLA_csc.scala 183:32:@24295.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_weight_channel_ext = NV_NVDLA_CSC_regfile_io_reg2dp_field_weight_channel_ext; // @[NV_NVDLA_csc.scala 184:39:@24296.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_entries = NV_NVDLA_CSC_regfile_io_reg2dp_field_entries; // @[NV_NVDLA_csc.scala 185:28:@24297.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_dataout_width = NV_NVDLA_CSC_regfile_io_reg2dp_field_dataout_width; // @[NV_NVDLA_csc.scala 186:34:@24298.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_rls_slices = NV_NVDLA_CSC_regfile_io_reg2dp_field_rls_slices; // @[NV_NVDLA_csc.scala 187:31:@24299.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_conv_x_stride_ext = NV_NVDLA_CSC_regfile_io_reg2dp_field_conv_x_stride_ext; // @[NV_NVDLA_csc.scala 188:38:@24300.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_conv_y_stride_ext = NV_NVDLA_CSC_regfile_io_reg2dp_field_conv_y_stride_ext; // @[NV_NVDLA_csc.scala 189:38:@24301.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_x_dilation_ext = NV_NVDLA_CSC_regfile_io_reg2dp_field_x_dilation_ext; // @[NV_NVDLA_csc.scala 190:35:@24302.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_y_dilation_ext = NV_NVDLA_CSC_regfile_io_reg2dp_field_y_dilation_ext; // @[NV_NVDLA_csc.scala 191:35:@24303.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_pad_left = NV_NVDLA_CSC_regfile_io_reg2dp_field_pad_left; // @[NV_NVDLA_csc.scala 192:29:@24304.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_pad_top = NV_NVDLA_CSC_regfile_io_reg2dp_field_pad_top; // @[NV_NVDLA_csc.scala 193:28:@24305.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_pad_value = NV_NVDLA_CSC_regfile_io_reg2dp_field_pad_value; // @[NV_NVDLA_csc.scala 194:30:@24306.4]
  assign NV_NVDLA_CSC_dl_io_reg2dp_data_bank = NV_NVDLA_CSC_regfile_io_reg2dp_field_data_bank; // @[NV_NVDLA_csc.scala 195:30:@24307.4]
  assign NV_NVDLA_slcg_io_nvdla_clock_nvdla_core_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_csc.scala 208:37:@24321.4]
  assign NV_NVDLA_slcg_1_io_nvdla_clock_nvdla_core_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_csc.scala 208:37:@24328.4]
  assign NV_NVDLA_slcg_2_io_nvdla_clock_nvdla_core_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_csc.scala 208:37:@24335.4]
endmodule
