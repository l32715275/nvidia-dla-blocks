// ================================================================
// NVDLA Open Source Project
//
// Copyright(c) 2016 - 2017 NVIDIA Corporation. Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with
// this distribution for more information.
// ================================================================
// File Name: NV_NVDLA_CMAC_CORE_mac.v
// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================
// File Name: NV_NVDLA_CMAC.h
module NV_NVDLA_CMAC_CORE_mac (
   nvdla_core_clk //|< i
  ,nvdla_wg_clk //|< i
  ,nvdla_core_rstn //|< i
  ,cfg_is_wg //|< i
  ,cfg_reg_en //|< i
  ,dat_actv_data //|< i
  ,dat_actv_nz //|< i
  ,dat_actv_pvld //|< i
  ,wt_actv_data //|< i
  ,wt_actv_nz //|< i
  ,wt_actv_pvld //|< i
  ,mac_out_data //|> o
  ,mac_out_pvld //|> o
  );
input nvdla_core_clk;
input nvdla_wg_clk;
input nvdla_core_rstn;
input cfg_is_wg;
input cfg_reg_en;
input [64*8 -1:0] dat_actv_data;
input [64 -1:0] dat_actv_nz;
input [64 -1:0] dat_actv_pvld;
input [64*8 -1:0] wt_actv_data;
input [64 -1:0] wt_actv_nz;
input [64 -1:0] wt_actv_pvld;
output [22 -1:0] mac_out_data;
output mac_out_pvld;

NV_NVDLA_CMAC_CORE_mac_dft NV_NVDLA_CMAC_CORE_mac_dft(
    .io_mac_out_valid(mac_out_pvld),
    .io_mac_out_bits(mac_out_data),
    .io_nvdla_core_clk(nvdla_core_clk),
    .io_nvdla_core_rstn(nvdla_core_rstn),
    .io_dat_actv_0_bits_data(dat_actv_data[7:0]),
    .io_dat_actv_1_bits_data(dat_actv_data[15:8]),
    .io_dat_actv_2_bits_data(dat_actv_data[23:16]),
    .io_dat_actv_3_bits_data(dat_actv_data[31:24]),
    .io_dat_actv_4_bits_data(dat_actv_data[39:32]),
    .io_dat_actv_5_bits_data(dat_actv_data[47:40]),
    .io_dat_actv_6_bits_data(dat_actv_data[55:48]),
    .io_dat_actv_7_bits_data(dat_actv_data[63:56]),
    .io_dat_actv_8_bits_data(dat_actv_data[71:64]),
    .io_dat_actv_9_bits_data(dat_actv_data[79:72]),
    .io_dat_actv_10_bits_data(dat_actv_data[87:80]),
    .io_dat_actv_11_bits_data(dat_actv_data[95:88]),
    .io_dat_actv_12_bits_data(dat_actv_data[103:96]),
    .io_dat_actv_13_bits_data(dat_actv_data[111:104]),
    .io_dat_actv_14_bits_data(dat_actv_data[119:112]),
    .io_dat_actv_15_bits_data(dat_actv_data[127:120]),
    .io_dat_actv_16_bits_data(dat_actv_data[135:128]),
    .io_dat_actv_17_bits_data(dat_actv_data[143:136]),
    .io_dat_actv_18_bits_data(dat_actv_data[151:144]),
    .io_dat_actv_19_bits_data(dat_actv_data[159:152]),
    .io_dat_actv_20_bits_data(dat_actv_data[167:160]),
    .io_dat_actv_21_bits_data(dat_actv_data[175:168]),
    .io_dat_actv_22_bits_data(dat_actv_data[183:176]),
    .io_dat_actv_23_bits_data(dat_actv_data[191:184]),
    .io_dat_actv_24_bits_data(dat_actv_data[199:192]),
    .io_dat_actv_25_bits_data(dat_actv_data[207:200]),
    .io_dat_actv_26_bits_data(dat_actv_data[215:208]),
    .io_dat_actv_27_bits_data(dat_actv_data[223:216]),
    .io_dat_actv_28_bits_data(dat_actv_data[231:224]),
    .io_dat_actv_29_bits_data(dat_actv_data[239:232]),
    .io_dat_actv_30_bits_data(dat_actv_data[247:240]),
    .io_dat_actv_31_bits_data(dat_actv_data[255:248]),
    .io_dat_actv_32_bits_data(dat_actv_data[263:256]),
    .io_dat_actv_33_bits_data(dat_actv_data[271:264]),
    .io_dat_actv_34_bits_data(dat_actv_data[279:272]),
    .io_dat_actv_35_bits_data(dat_actv_data[287:280]),
    .io_dat_actv_36_bits_data(dat_actv_data[295:288]),
    .io_dat_actv_37_bits_data(dat_actv_data[303:296]),
    .io_dat_actv_38_bits_data(dat_actv_data[311:304]),
    .io_dat_actv_39_bits_data(dat_actv_data[319:312]),
    .io_dat_actv_40_bits_data(dat_actv_data[327:320]),
    .io_dat_actv_41_bits_data(dat_actv_data[335:328]),
    .io_dat_actv_42_bits_data(dat_actv_data[343:336]),
    .io_dat_actv_43_bits_data(dat_actv_data[351:344]),
    .io_dat_actv_44_bits_data(dat_actv_data[359:352]),
    .io_dat_actv_45_bits_data(dat_actv_data[367:360]),
    .io_dat_actv_46_bits_data(dat_actv_data[375:368]),
    .io_dat_actv_47_bits_data(dat_actv_data[383:376]),
    .io_dat_actv_48_bits_data(dat_actv_data[391:384]),
    .io_dat_actv_49_bits_data(dat_actv_data[399:392]),
    .io_dat_actv_50_bits_data(dat_actv_data[407:400]),
    .io_dat_actv_51_bits_data(dat_actv_data[415:408]),
    .io_dat_actv_52_bits_data(dat_actv_data[423:416]),
    .io_dat_actv_53_bits_data(dat_actv_data[431:424]),
    .io_dat_actv_54_bits_data(dat_actv_data[439:432]),
    .io_dat_actv_55_bits_data(dat_actv_data[447:440]),
    .io_dat_actv_56_bits_data(dat_actv_data[455:448]),
    .io_dat_actv_57_bits_data(dat_actv_data[463:456]),
    .io_dat_actv_58_bits_data(dat_actv_data[471:464]),
    .io_dat_actv_59_bits_data(dat_actv_data[479:472]),
    .io_dat_actv_60_bits_data(dat_actv_data[487:480]),
    .io_dat_actv_61_bits_data(dat_actv_data[495:488]),
    .io_dat_actv_62_bits_data(dat_actv_data[503:496]),
    .io_dat_actv_63_bits_data(dat_actv_data[511:504]),
    .io_dat_actv_0_bits_nz(dat_actv_nz[0]),
    .io_dat_actv_1_bits_nz(dat_actv_nz[1]),
    .io_dat_actv_2_bits_nz(dat_actv_nz[2]),
    .io_dat_actv_3_bits_nz(dat_actv_nz[3]),
    .io_dat_actv_4_bits_nz(dat_actv_nz[4]),
    .io_dat_actv_5_bits_nz(dat_actv_nz[5]),
    .io_dat_actv_6_bits_nz(dat_actv_nz[6]),
    .io_dat_actv_7_bits_nz(dat_actv_nz[7]),
    .io_dat_actv_8_bits_nz(dat_actv_nz[8]),
    .io_dat_actv_9_bits_nz(dat_actv_nz[9]),
    .io_dat_actv_10_bits_nz(dat_actv_nz[10]),
    .io_dat_actv_11_bits_nz(dat_actv_nz[11]),
    .io_dat_actv_12_bits_nz(dat_actv_nz[12]),
    .io_dat_actv_13_bits_nz(dat_actv_nz[13]),
    .io_dat_actv_14_bits_nz(dat_actv_nz[14]),
    .io_dat_actv_15_bits_nz(dat_actv_nz[15]),
    .io_dat_actv_16_bits_nz(dat_actv_nz[16]),
    .io_dat_actv_17_bits_nz(dat_actv_nz[17]),
    .io_dat_actv_18_bits_nz(dat_actv_nz[18]),
    .io_dat_actv_19_bits_nz(dat_actv_nz[19]),
    .io_dat_actv_20_bits_nz(dat_actv_nz[20]),
    .io_dat_actv_21_bits_nz(dat_actv_nz[21]),
    .io_dat_actv_22_bits_nz(dat_actv_nz[22]),
    .io_dat_actv_23_bits_nz(dat_actv_nz[23]),
    .io_dat_actv_24_bits_nz(dat_actv_nz[24]),
    .io_dat_actv_25_bits_nz(dat_actv_nz[25]),
    .io_dat_actv_26_bits_nz(dat_actv_nz[26]),
    .io_dat_actv_27_bits_nz(dat_actv_nz[27]),
    .io_dat_actv_28_bits_nz(dat_actv_nz[28]),
    .io_dat_actv_29_bits_nz(dat_actv_nz[29]),
    .io_dat_actv_30_bits_nz(dat_actv_nz[30]),
    .io_dat_actv_31_bits_nz(dat_actv_nz[31]),
    .io_dat_actv_32_bits_nz(dat_actv_nz[32]),
    .io_dat_actv_33_bits_nz(dat_actv_nz[33]),
    .io_dat_actv_34_bits_nz(dat_actv_nz[34]),
    .io_dat_actv_35_bits_nz(dat_actv_nz[35]),
    .io_dat_actv_36_bits_nz(dat_actv_nz[36]),
    .io_dat_actv_37_bits_nz(dat_actv_nz[37]),
    .io_dat_actv_38_bits_nz(dat_actv_nz[38]),
    .io_dat_actv_39_bits_nz(dat_actv_nz[39]),
    .io_dat_actv_40_bits_nz(dat_actv_nz[40]),
    .io_dat_actv_41_bits_nz(dat_actv_nz[41]),
    .io_dat_actv_42_bits_nz(dat_actv_nz[42]),
    .io_dat_actv_43_bits_nz(dat_actv_nz[43]),
    .io_dat_actv_44_bits_nz(dat_actv_nz[44]),
    .io_dat_actv_45_bits_nz(dat_actv_nz[45]),
    .io_dat_actv_46_bits_nz(dat_actv_nz[46]),
    .io_dat_actv_47_bits_nz(dat_actv_nz[47]),
    .io_dat_actv_48_bits_nz(dat_actv_nz[48]),
    .io_dat_actv_49_bits_nz(dat_actv_nz[49]),
    .io_dat_actv_50_bits_nz(dat_actv_nz[50]),
    .io_dat_actv_51_bits_nz(dat_actv_nz[51]),
    .io_dat_actv_52_bits_nz(dat_actv_nz[52]),
    .io_dat_actv_53_bits_nz(dat_actv_nz[53]),
    .io_dat_actv_54_bits_nz(dat_actv_nz[54]),
    .io_dat_actv_55_bits_nz(dat_actv_nz[55]),
    .io_dat_actv_56_bits_nz(dat_actv_nz[56]),
    .io_dat_actv_57_bits_nz(dat_actv_nz[57]),
    .io_dat_actv_58_bits_nz(dat_actv_nz[58]),
    .io_dat_actv_59_bits_nz(dat_actv_nz[59]),
    .io_dat_actv_60_bits_nz(dat_actv_nz[60]),
    .io_dat_actv_61_bits_nz(dat_actv_nz[61]),
    .io_dat_actv_62_bits_nz(dat_actv_nz[62]),
    .io_dat_actv_63_bits_nz(dat_actv_nz[63]),
    .io_dat_actv_0_valid(dat_actv_pvld[0]),
    .io_dat_actv_1_valid(dat_actv_pvld[1]),
    .io_dat_actv_2_valid(dat_actv_pvld[2]),
    .io_dat_actv_3_valid(dat_actv_pvld[3]),
    .io_dat_actv_4_valid(dat_actv_pvld[4]),
    .io_dat_actv_5_valid(dat_actv_pvld[5]),
    .io_dat_actv_6_valid(dat_actv_pvld[6]),
    .io_dat_actv_7_valid(dat_actv_pvld[7]),
    .io_dat_actv_8_valid(dat_actv_pvld[8]),
    .io_dat_actv_9_valid(dat_actv_pvld[9]),
    .io_dat_actv_10_valid(dat_actv_pvld[10]),
    .io_dat_actv_11_valid(dat_actv_pvld[11]),
    .io_dat_actv_12_valid(dat_actv_pvld[12]),
    .io_dat_actv_13_valid(dat_actv_pvld[13]),
    .io_dat_actv_14_valid(dat_actv_pvld[14]),
    .io_dat_actv_15_valid(dat_actv_pvld[15]),
    .io_dat_actv_16_valid(dat_actv_pvld[16]),
    .io_dat_actv_17_valid(dat_actv_pvld[17]),
    .io_dat_actv_18_valid(dat_actv_pvld[18]),
    .io_dat_actv_19_valid(dat_actv_pvld[19]),
    .io_dat_actv_20_valid(dat_actv_pvld[20]),
    .io_dat_actv_21_valid(dat_actv_pvld[21]),
    .io_dat_actv_22_valid(dat_actv_pvld[22]),
    .io_dat_actv_23_valid(dat_actv_pvld[23]),
    .io_dat_actv_24_valid(dat_actv_pvld[24]),
    .io_dat_actv_25_valid(dat_actv_pvld[25]),
    .io_dat_actv_26_valid(dat_actv_pvld[26]),
    .io_dat_actv_27_valid(dat_actv_pvld[27]),
    .io_dat_actv_28_valid(dat_actv_pvld[28]),
    .io_dat_actv_29_valid(dat_actv_pvld[29]),
    .io_dat_actv_30_valid(dat_actv_pvld[30]),
    .io_dat_actv_31_valid(dat_actv_pvld[31]),
    .io_dat_actv_32_valid(dat_actv_pvld[32]),
    .io_dat_actv_33_valid(dat_actv_pvld[33]),
    .io_dat_actv_34_valid(dat_actv_pvld[34]),
    .io_dat_actv_35_valid(dat_actv_pvld[35]),
    .io_dat_actv_36_valid(dat_actv_pvld[36]),
    .io_dat_actv_37_valid(dat_actv_pvld[37]),
    .io_dat_actv_38_valid(dat_actv_pvld[38]),
    .io_dat_actv_39_valid(dat_actv_pvld[39]),
    .io_dat_actv_40_valid(dat_actv_pvld[40]),
    .io_dat_actv_41_valid(dat_actv_pvld[41]),
    .io_dat_actv_42_valid(dat_actv_pvld[42]),
    .io_dat_actv_43_valid(dat_actv_pvld[43]),
    .io_dat_actv_44_valid(dat_actv_pvld[44]),
    .io_dat_actv_45_valid(dat_actv_pvld[45]),
    .io_dat_actv_46_valid(dat_actv_pvld[46]),
    .io_dat_actv_47_valid(dat_actv_pvld[47]),
    .io_dat_actv_48_valid(dat_actv_pvld[48]),
    .io_dat_actv_49_valid(dat_actv_pvld[49]),
    .io_dat_actv_50_valid(dat_actv_pvld[50]),
    .io_dat_actv_51_valid(dat_actv_pvld[51]),
    .io_dat_actv_52_valid(dat_actv_pvld[52]),
    .io_dat_actv_53_valid(dat_actv_pvld[53]),
    .io_dat_actv_54_valid(dat_actv_pvld[54]),
    .io_dat_actv_55_valid(dat_actv_pvld[55]),
    .io_dat_actv_56_valid(dat_actv_pvld[56]),
    .io_dat_actv_57_valid(dat_actv_pvld[57]),
    .io_dat_actv_58_valid(dat_actv_pvld[58]),
    .io_dat_actv_59_valid(dat_actv_pvld[59]),
    .io_dat_actv_60_valid(dat_actv_pvld[60]),
    .io_dat_actv_61_valid(dat_actv_pvld[61]),
    .io_dat_actv_62_valid(dat_actv_pvld[62]),
    .io_dat_actv_63_valid(dat_actv_pvld[63]),
    .io_wt_actv_0_bits_data(wt_actv_data[7:0]),
    .io_wt_actv_1_bits_data(wt_actv_data[15:8]),
    .io_wt_actv_2_bits_data(wt_actv_data[23:16]),
    .io_wt_actv_3_bits_data(wt_actv_data[31:24]),
    .io_wt_actv_4_bits_data(wt_actv_data[39:32]),
    .io_wt_actv_5_bits_data(wt_actv_data[47:40]),
    .io_wt_actv_6_bits_data(wt_actv_data[55:48]),
    .io_wt_actv_7_bits_data(wt_actv_data[63:56]),
    .io_wt_actv_8_bits_data(wt_actv_data[71:64]),
    .io_wt_actv_9_bits_data(wt_actv_data[79:72]),
    .io_wt_actv_10_bits_data(wt_actv_data[87:80]),
    .io_wt_actv_11_bits_data(wt_actv_data[95:88]),
    .io_wt_actv_12_bits_data(wt_actv_data[103:96]),
    .io_wt_actv_13_bits_data(wt_actv_data[111:104]),
    .io_wt_actv_14_bits_data(wt_actv_data[119:112]),
    .io_wt_actv_15_bits_data(wt_actv_data[127:120]),
    .io_wt_actv_16_bits_data(wt_actv_data[135:128]),
    .io_wt_actv_17_bits_data(wt_actv_data[143:136]),
    .io_wt_actv_18_bits_data(wt_actv_data[151:144]),
    .io_wt_actv_19_bits_data(wt_actv_data[159:152]),
    .io_wt_actv_20_bits_data(wt_actv_data[167:160]),
    .io_wt_actv_21_bits_data(wt_actv_data[175:168]),
    .io_wt_actv_22_bits_data(wt_actv_data[183:176]),
    .io_wt_actv_23_bits_data(wt_actv_data[191:184]),
    .io_wt_actv_24_bits_data(wt_actv_data[199:192]),
    .io_wt_actv_25_bits_data(wt_actv_data[207:200]),
    .io_wt_actv_26_bits_data(wt_actv_data[215:208]),
    .io_wt_actv_27_bits_data(wt_actv_data[223:216]),
    .io_wt_actv_28_bits_data(wt_actv_data[231:224]),
    .io_wt_actv_29_bits_data(wt_actv_data[239:232]),
    .io_wt_actv_30_bits_data(wt_actv_data[247:240]),
    .io_wt_actv_31_bits_data(wt_actv_data[255:248]),
    .io_wt_actv_32_bits_data(wt_actv_data[263:256]),
    .io_wt_actv_33_bits_data(wt_actv_data[271:264]),
    .io_wt_actv_34_bits_data(wt_actv_data[279:272]),
    .io_wt_actv_35_bits_data(wt_actv_data[287:280]),
    .io_wt_actv_36_bits_data(wt_actv_data[295:288]),
    .io_wt_actv_37_bits_data(wt_actv_data[303:296]),
    .io_wt_actv_38_bits_data(wt_actv_data[311:304]),
    .io_wt_actv_39_bits_data(wt_actv_data[319:312]),
    .io_wt_actv_40_bits_data(wt_actv_data[327:320]),
    .io_wt_actv_41_bits_data(wt_actv_data[335:328]),
    .io_wt_actv_42_bits_data(wt_actv_data[343:336]),
    .io_wt_actv_43_bits_data(wt_actv_data[351:344]),
    .io_wt_actv_44_bits_data(wt_actv_data[359:352]),
    .io_wt_actv_45_bits_data(wt_actv_data[367:360]),
    .io_wt_actv_46_bits_data(wt_actv_data[375:368]),
    .io_wt_actv_47_bits_data(wt_actv_data[383:376]),
    .io_wt_actv_48_bits_data(wt_actv_data[391:384]),
    .io_wt_actv_49_bits_data(wt_actv_data[399:392]),
    .io_wt_actv_50_bits_data(wt_actv_data[407:400]),
    .io_wt_actv_51_bits_data(wt_actv_data[415:408]),
    .io_wt_actv_52_bits_data(wt_actv_data[423:416]),
    .io_wt_actv_53_bits_data(wt_actv_data[431:424]),
    .io_wt_actv_54_bits_data(wt_actv_data[439:432]),
    .io_wt_actv_55_bits_data(wt_actv_data[447:440]),
    .io_wt_actv_56_bits_data(wt_actv_data[455:448]),
    .io_wt_actv_57_bits_data(wt_actv_data[463:456]),
    .io_wt_actv_58_bits_data(wt_actv_data[471:464]),
    .io_wt_actv_59_bits_data(wt_actv_data[479:472]),
    .io_wt_actv_60_bits_data(wt_actv_data[487:480]),
    .io_wt_actv_61_bits_data(wt_actv_data[495:488]),
    .io_wt_actv_62_bits_data(wt_actv_data[503:496]),
    .io_wt_actv_63_bits_data(wt_actv_data[511:504]),
    .io_wt_actv_0_bits_nz(wt_actv_nz[0]),
    .io_wt_actv_1_bits_nz(wt_actv_nz[1]),
    .io_wt_actv_2_bits_nz(wt_actv_nz[2]),
    .io_wt_actv_3_bits_nz(wt_actv_nz[3]),
    .io_wt_actv_4_bits_nz(wt_actv_nz[4]),
    .io_wt_actv_5_bits_nz(wt_actv_nz[5]),
    .io_wt_actv_6_bits_nz(wt_actv_nz[6]),
    .io_wt_actv_7_bits_nz(wt_actv_nz[7]),
    .io_wt_actv_8_bits_nz(wt_actv_nz[8]),
    .io_wt_actv_9_bits_nz(wt_actv_nz[9]),
    .io_wt_actv_10_bits_nz(wt_actv_nz[10]),
    .io_wt_actv_11_bits_nz(wt_actv_nz[11]),
    .io_wt_actv_12_bits_nz(wt_actv_nz[12]),
    .io_wt_actv_13_bits_nz(wt_actv_nz[13]),
    .io_wt_actv_14_bits_nz(wt_actv_nz[14]),
    .io_wt_actv_15_bits_nz(wt_actv_nz[15]),
    .io_wt_actv_16_bits_nz(wt_actv_nz[16]),
    .io_wt_actv_17_bits_nz(wt_actv_nz[17]),
    .io_wt_actv_18_bits_nz(wt_actv_nz[18]),
    .io_wt_actv_19_bits_nz(wt_actv_nz[19]),
    .io_wt_actv_20_bits_nz(wt_actv_nz[20]),
    .io_wt_actv_21_bits_nz(wt_actv_nz[21]),
    .io_wt_actv_22_bits_nz(wt_actv_nz[22]),
    .io_wt_actv_23_bits_nz(wt_actv_nz[23]),
    .io_wt_actv_24_bits_nz(wt_actv_nz[24]),
    .io_wt_actv_25_bits_nz(wt_actv_nz[25]),
    .io_wt_actv_26_bits_nz(wt_actv_nz[26]),
    .io_wt_actv_27_bits_nz(wt_actv_nz[27]),
    .io_wt_actv_28_bits_nz(wt_actv_nz[28]),
    .io_wt_actv_29_bits_nz(wt_actv_nz[29]),
    .io_wt_actv_30_bits_nz(wt_actv_nz[30]),
    .io_wt_actv_31_bits_nz(wt_actv_nz[31]),
    .io_wt_actv_32_bits_nz(wt_actv_nz[32]),
    .io_wt_actv_33_bits_nz(wt_actv_nz[33]),
    .io_wt_actv_34_bits_nz(wt_actv_nz[34]),
    .io_wt_actv_35_bits_nz(wt_actv_nz[35]),
    .io_wt_actv_36_bits_nz(wt_actv_nz[36]),
    .io_wt_actv_37_bits_nz(wt_actv_nz[37]),
    .io_wt_actv_38_bits_nz(wt_actv_nz[38]),
    .io_wt_actv_39_bits_nz(wt_actv_nz[39]),
    .io_wt_actv_40_bits_nz(wt_actv_nz[40]),
    .io_wt_actv_41_bits_nz(wt_actv_nz[41]),
    .io_wt_actv_42_bits_nz(wt_actv_nz[42]),
    .io_wt_actv_43_bits_nz(wt_actv_nz[43]),
    .io_wt_actv_44_bits_nz(wt_actv_nz[44]),
    .io_wt_actv_45_bits_nz(wt_actv_nz[45]),
    .io_wt_actv_46_bits_nz(wt_actv_nz[46]),
    .io_wt_actv_47_bits_nz(wt_actv_nz[47]),
    .io_wt_actv_48_bits_nz(wt_actv_nz[48]),
    .io_wt_actv_49_bits_nz(wt_actv_nz[49]),
    .io_wt_actv_50_bits_nz(wt_actv_nz[50]),
    .io_wt_actv_51_bits_nz(wt_actv_nz[51]),
    .io_wt_actv_52_bits_nz(wt_actv_nz[52]),
    .io_wt_actv_53_bits_nz(wt_actv_nz[53]),
    .io_wt_actv_54_bits_nz(wt_actv_nz[54]),
    .io_wt_actv_55_bits_nz(wt_actv_nz[55]),
    .io_wt_actv_56_bits_nz(wt_actv_nz[56]),
    .io_wt_actv_57_bits_nz(wt_actv_nz[57]),
    .io_wt_actv_58_bits_nz(wt_actv_nz[58]),
    .io_wt_actv_59_bits_nz(wt_actv_nz[59]),
    .io_wt_actv_60_bits_nz(wt_actv_nz[60]),
    .io_wt_actv_61_bits_nz(wt_actv_nz[61]),
    .io_wt_actv_62_bits_nz(wt_actv_nz[62]),
    .io_wt_actv_63_bits_nz(wt_actv_nz[63]),
    .io_wt_actv_0_valid(wt_actv_pvld[0]),
    .io_wt_actv_1_valid(wt_actv_pvld[1]),
    .io_wt_actv_2_valid(wt_actv_pvld[2]),
    .io_wt_actv_3_valid(wt_actv_pvld[3]),
    .io_wt_actv_4_valid(wt_actv_pvld[4]),
    .io_wt_actv_5_valid(wt_actv_pvld[5]),
    .io_wt_actv_6_valid(wt_actv_pvld[6]),
    .io_wt_actv_7_valid(wt_actv_pvld[7]),
    .io_wt_actv_8_valid(wt_actv_pvld[8]),
    .io_wt_actv_9_valid(wt_actv_pvld[9]),
    .io_wt_actv_10_valid(wt_actv_pvld[10]),
    .io_wt_actv_11_valid(wt_actv_pvld[11]),
    .io_wt_actv_12_valid(wt_actv_pvld[12]),
    .io_wt_actv_13_valid(wt_actv_pvld[13]),
    .io_wt_actv_14_valid(wt_actv_pvld[14]),
    .io_wt_actv_15_valid(wt_actv_pvld[15]),
    .io_wt_actv_16_valid(wt_actv_pvld[16]),
    .io_wt_actv_17_valid(wt_actv_pvld[17]),
    .io_wt_actv_18_valid(wt_actv_pvld[18]),
    .io_wt_actv_19_valid(wt_actv_pvld[19]),
    .io_wt_actv_20_valid(wt_actv_pvld[20]),
    .io_wt_actv_21_valid(wt_actv_pvld[21]),
    .io_wt_actv_22_valid(wt_actv_pvld[22]),
    .io_wt_actv_23_valid(wt_actv_pvld[23]),
    .io_wt_actv_24_valid(wt_actv_pvld[24]),
    .io_wt_actv_25_valid(wt_actv_pvld[25]),
    .io_wt_actv_26_valid(wt_actv_pvld[26]),
    .io_wt_actv_27_valid(wt_actv_pvld[27]),
    .io_wt_actv_28_valid(wt_actv_pvld[28]),
    .io_wt_actv_29_valid(wt_actv_pvld[29]),
    .io_wt_actv_30_valid(wt_actv_pvld[30]),
    .io_wt_actv_31_valid(wt_actv_pvld[31]),
    .io_wt_actv_32_valid(wt_actv_pvld[32]),
    .io_wt_actv_33_valid(wt_actv_pvld[33]),
    .io_wt_actv_34_valid(wt_actv_pvld[34]),
    .io_wt_actv_35_valid(wt_actv_pvld[35]),
    .io_wt_actv_36_valid(wt_actv_pvld[36]),
    .io_wt_actv_37_valid(wt_actv_pvld[37]),
    .io_wt_actv_38_valid(wt_actv_pvld[38]),
    .io_wt_actv_39_valid(wt_actv_pvld[39]),
    .io_wt_actv_40_valid(wt_actv_pvld[40]),
    .io_wt_actv_41_valid(wt_actv_pvld[41]),
    .io_wt_actv_42_valid(wt_actv_pvld[42]),
    .io_wt_actv_43_valid(wt_actv_pvld[43]),
    .io_wt_actv_44_valid(wt_actv_pvld[44]),
    .io_wt_actv_45_valid(wt_actv_pvld[45]),
    .io_wt_actv_46_valid(wt_actv_pvld[46]),
    .io_wt_actv_47_valid(wt_actv_pvld[47]),
    .io_wt_actv_48_valid(wt_actv_pvld[48]),
    .io_wt_actv_49_valid(wt_actv_pvld[49]),
    .io_wt_actv_50_valid(wt_actv_pvld[50]),
    .io_wt_actv_51_valid(wt_actv_pvld[51]),
    .io_wt_actv_52_valid(wt_actv_pvld[52]),
    .io_wt_actv_53_valid(wt_actv_pvld[53]),
    .io_wt_actv_54_valid(wt_actv_pvld[54]),
    .io_wt_actv_55_valid(wt_actv_pvld[55]),
    .io_wt_actv_56_valid(wt_actv_pvld[56]),
    .io_wt_actv_57_valid(wt_actv_pvld[57]),
    .io_wt_actv_58_valid(wt_actv_pvld[58]),
    .io_wt_actv_59_valid(wt_actv_pvld[59]),
    .io_wt_actv_60_valid(wt_actv_pvld[60]),
    .io_wt_actv_61_valid(wt_actv_pvld[61]),
    .io_wt_actv_62_valid(wt_actv_pvld[62]),
    .io_wt_actv_63_valid(wt_actv_pvld[63])
);
endmodule