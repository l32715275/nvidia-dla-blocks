module nv_ram_rws( // @[:@3.2]
  input          io_clk, // @[:@6.4]
  input          io_re, // @[:@6.4]
  input          io_we, // @[:@6.4]
  input  [8:0]   io_ra, // @[:@6.4]
  input  [8:0]   io_wa, // @[:@6.4]
  input  [255:0] io_di, // @[:@6.4]
  output [255:0] io_dout // @[:@6.4]
);
  reg [255:0] _T_22_0; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_0;
  reg [255:0] _T_22_1; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_1;
  reg [255:0] _T_22_2; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_2;
  reg [255:0] _T_22_3; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_3;
  reg [255:0] _T_22_4; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_4;
  reg [255:0] _T_22_5; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_5;
  reg [255:0] _T_22_6; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_6;
  reg [255:0] _T_22_7; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_7;
  reg [255:0] _T_22_8; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_8;
  reg [255:0] _T_22_9; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_9;
  reg [255:0] _T_22_10; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_10;
  reg [255:0] _T_22_11; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_11;
  reg [255:0] _T_22_12; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_12;
  reg [255:0] _T_22_13; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_13;
  reg [255:0] _T_22_14; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_14;
  reg [255:0] _T_22_15; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_15;
  reg [255:0] _T_22_16; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_16;
  reg [255:0] _T_22_17; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_17;
  reg [255:0] _T_22_18; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_18;
  reg [255:0] _T_22_19; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_19;
  reg [255:0] _T_22_20; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_20;
  reg [255:0] _T_22_21; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_21;
  reg [255:0] _T_22_22; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_22;
  reg [255:0] _T_22_23; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_23;
  reg [255:0] _T_22_24; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_24;
  reg [255:0] _T_22_25; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_25;
  reg [255:0] _T_22_26; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_26;
  reg [255:0] _T_22_27; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_27;
  reg [255:0] _T_22_28; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_28;
  reg [255:0] _T_22_29; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_29;
  reg [255:0] _T_22_30; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_30;
  reg [255:0] _T_22_31; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_31;
  reg [255:0] _T_22_32; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_32;
  reg [255:0] _T_22_33; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_33;
  reg [255:0] _T_22_34; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_34;
  reg [255:0] _T_22_35; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_35;
  reg [255:0] _T_22_36; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_36;
  reg [255:0] _T_22_37; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_37;
  reg [255:0] _T_22_38; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_38;
  reg [255:0] _T_22_39; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_39;
  reg [255:0] _T_22_40; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_40;
  reg [255:0] _T_22_41; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_41;
  reg [255:0] _T_22_42; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_42;
  reg [255:0] _T_22_43; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_43;
  reg [255:0] _T_22_44; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_44;
  reg [255:0] _T_22_45; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_45;
  reg [255:0] _T_22_46; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_46;
  reg [255:0] _T_22_47; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_47;
  reg [255:0] _T_22_48; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_48;
  reg [255:0] _T_22_49; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_49;
  reg [255:0] _T_22_50; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_50;
  reg [255:0] _T_22_51; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_51;
  reg [255:0] _T_22_52; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_52;
  reg [255:0] _T_22_53; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_53;
  reg [255:0] _T_22_54; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_54;
  reg [255:0] _T_22_55; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_55;
  reg [255:0] _T_22_56; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_56;
  reg [255:0] _T_22_57; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_57;
  reg [255:0] _T_22_58; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_58;
  reg [255:0] _T_22_59; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_59;
  reg [255:0] _T_22_60; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_60;
  reg [255:0] _T_22_61; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_61;
  reg [255:0] _T_22_62; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_62;
  reg [255:0] _T_22_63; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_63;
  reg [255:0] _T_22_64; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_64;
  reg [255:0] _T_22_65; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_65;
  reg [255:0] _T_22_66; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_66;
  reg [255:0] _T_22_67; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_67;
  reg [255:0] _T_22_68; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_68;
  reg [255:0] _T_22_69; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_69;
  reg [255:0] _T_22_70; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_70;
  reg [255:0] _T_22_71; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_71;
  reg [255:0] _T_22_72; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_72;
  reg [255:0] _T_22_73; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_73;
  reg [255:0] _T_22_74; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_74;
  reg [255:0] _T_22_75; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_75;
  reg [255:0] _T_22_76; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_76;
  reg [255:0] _T_22_77; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_77;
  reg [255:0] _T_22_78; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_78;
  reg [255:0] _T_22_79; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_79;
  reg [255:0] _T_22_80; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_80;
  reg [255:0] _T_22_81; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_81;
  reg [255:0] _T_22_82; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_82;
  reg [255:0] _T_22_83; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_83;
  reg [255:0] _T_22_84; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_84;
  reg [255:0] _T_22_85; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_85;
  reg [255:0] _T_22_86; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_86;
  reg [255:0] _T_22_87; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_87;
  reg [255:0] _T_22_88; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_88;
  reg [255:0] _T_22_89; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_89;
  reg [255:0] _T_22_90; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_90;
  reg [255:0] _T_22_91; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_91;
  reg [255:0] _T_22_92; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_92;
  reg [255:0] _T_22_93; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_93;
  reg [255:0] _T_22_94; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_94;
  reg [255:0] _T_22_95; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_95;
  reg [255:0] _T_22_96; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_96;
  reg [255:0] _T_22_97; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_97;
  reg [255:0] _T_22_98; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_98;
  reg [255:0] _T_22_99; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_99;
  reg [255:0] _T_22_100; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_100;
  reg [255:0] _T_22_101; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_101;
  reg [255:0] _T_22_102; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_102;
  reg [255:0] _T_22_103; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_103;
  reg [255:0] _T_22_104; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_104;
  reg [255:0] _T_22_105; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_105;
  reg [255:0] _T_22_106; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_106;
  reg [255:0] _T_22_107; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_107;
  reg [255:0] _T_22_108; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_108;
  reg [255:0] _T_22_109; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_109;
  reg [255:0] _T_22_110; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_110;
  reg [255:0] _T_22_111; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_111;
  reg [255:0] _T_22_112; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_112;
  reg [255:0] _T_22_113; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_113;
  reg [255:0] _T_22_114; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_114;
  reg [255:0] _T_22_115; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_115;
  reg [255:0] _T_22_116; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_116;
  reg [255:0] _T_22_117; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_117;
  reg [255:0] _T_22_118; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_118;
  reg [255:0] _T_22_119; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_119;
  reg [255:0] _T_22_120; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_120;
  reg [255:0] _T_22_121; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_121;
  reg [255:0] _T_22_122; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_122;
  reg [255:0] _T_22_123; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_123;
  reg [255:0] _T_22_124; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_124;
  reg [255:0] _T_22_125; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_125;
  reg [255:0] _T_22_126; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_126;
  reg [255:0] _T_22_127; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_127;
  reg [255:0] _T_22_128; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_128;
  reg [255:0] _T_22_129; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_129;
  reg [255:0] _T_22_130; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_130;
  reg [255:0] _T_22_131; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_131;
  reg [255:0] _T_22_132; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_132;
  reg [255:0] _T_22_133; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_133;
  reg [255:0] _T_22_134; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_134;
  reg [255:0] _T_22_135; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_135;
  reg [255:0] _T_22_136; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_136;
  reg [255:0] _T_22_137; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_137;
  reg [255:0] _T_22_138; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_138;
  reg [255:0] _T_22_139; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_139;
  reg [255:0] _T_22_140; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_140;
  reg [255:0] _T_22_141; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_141;
  reg [255:0] _T_22_142; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_142;
  reg [255:0] _T_22_143; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_143;
  reg [255:0] _T_22_144; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_144;
  reg [255:0] _T_22_145; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_145;
  reg [255:0] _T_22_146; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_146;
  reg [255:0] _T_22_147; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_147;
  reg [255:0] _T_22_148; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_148;
  reg [255:0] _T_22_149; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_149;
  reg [255:0] _T_22_150; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_150;
  reg [255:0] _T_22_151; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_151;
  reg [255:0] _T_22_152; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_152;
  reg [255:0] _T_22_153; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_153;
  reg [255:0] _T_22_154; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_154;
  reg [255:0] _T_22_155; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_155;
  reg [255:0] _T_22_156; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_156;
  reg [255:0] _T_22_157; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_157;
  reg [255:0] _T_22_158; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_158;
  reg [255:0] _T_22_159; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_159;
  reg [255:0] _T_22_160; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_160;
  reg [255:0] _T_22_161; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_161;
  reg [255:0] _T_22_162; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_162;
  reg [255:0] _T_22_163; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_163;
  reg [255:0] _T_22_164; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_164;
  reg [255:0] _T_22_165; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_165;
  reg [255:0] _T_22_166; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_166;
  reg [255:0] _T_22_167; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_167;
  reg [255:0] _T_22_168; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_168;
  reg [255:0] _T_22_169; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_169;
  reg [255:0] _T_22_170; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_170;
  reg [255:0] _T_22_171; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_171;
  reg [255:0] _T_22_172; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_172;
  reg [255:0] _T_22_173; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_173;
  reg [255:0] _T_22_174; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_174;
  reg [255:0] _T_22_175; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_175;
  reg [255:0] _T_22_176; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_176;
  reg [255:0] _T_22_177; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_177;
  reg [255:0] _T_22_178; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_178;
  reg [255:0] _T_22_179; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_179;
  reg [255:0] _T_22_180; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_180;
  reg [255:0] _T_22_181; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_181;
  reg [255:0] _T_22_182; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_182;
  reg [255:0] _T_22_183; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_183;
  reg [255:0] _T_22_184; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_184;
  reg [255:0] _T_22_185; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_185;
  reg [255:0] _T_22_186; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_186;
  reg [255:0] _T_22_187; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_187;
  reg [255:0] _T_22_188; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_188;
  reg [255:0] _T_22_189; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_189;
  reg [255:0] _T_22_190; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_190;
  reg [255:0] _T_22_191; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_191;
  reg [255:0] _T_22_192; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_192;
  reg [255:0] _T_22_193; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_193;
  reg [255:0] _T_22_194; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_194;
  reg [255:0] _T_22_195; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_195;
  reg [255:0] _T_22_196; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_196;
  reg [255:0] _T_22_197; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_197;
  reg [255:0] _T_22_198; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_198;
  reg [255:0] _T_22_199; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_199;
  reg [255:0] _T_22_200; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_200;
  reg [255:0] _T_22_201; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_201;
  reg [255:0] _T_22_202; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_202;
  reg [255:0] _T_22_203; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_203;
  reg [255:0] _T_22_204; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_204;
  reg [255:0] _T_22_205; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_205;
  reg [255:0] _T_22_206; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_206;
  reg [255:0] _T_22_207; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_207;
  reg [255:0] _T_22_208; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_208;
  reg [255:0] _T_22_209; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_209;
  reg [255:0] _T_22_210; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_210;
  reg [255:0] _T_22_211; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_211;
  reg [255:0] _T_22_212; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_212;
  reg [255:0] _T_22_213; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_213;
  reg [255:0] _T_22_214; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_214;
  reg [255:0] _T_22_215; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_215;
  reg [255:0] _T_22_216; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_216;
  reg [255:0] _T_22_217; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_217;
  reg [255:0] _T_22_218; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_218;
  reg [255:0] _T_22_219; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_219;
  reg [255:0] _T_22_220; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_220;
  reg [255:0] _T_22_221; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_221;
  reg [255:0] _T_22_222; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_222;
  reg [255:0] _T_22_223; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_223;
  reg [255:0] _T_22_224; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_224;
  reg [255:0] _T_22_225; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_225;
  reg [255:0] _T_22_226; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_226;
  reg [255:0] _T_22_227; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_227;
  reg [255:0] _T_22_228; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_228;
  reg [255:0] _T_22_229; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_229;
  reg [255:0] _T_22_230; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_230;
  reg [255:0] _T_22_231; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_231;
  reg [255:0] _T_22_232; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_232;
  reg [255:0] _T_22_233; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_233;
  reg [255:0] _T_22_234; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_234;
  reg [255:0] _T_22_235; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_235;
  reg [255:0] _T_22_236; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_236;
  reg [255:0] _T_22_237; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_237;
  reg [255:0] _T_22_238; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_238;
  reg [255:0] _T_22_239; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_239;
  reg [255:0] _T_22_240; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_240;
  reg [255:0] _T_22_241; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_241;
  reg [255:0] _T_22_242; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_242;
  reg [255:0] _T_22_243; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_243;
  reg [255:0] _T_22_244; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_244;
  reg [255:0] _T_22_245; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_245;
  reg [255:0] _T_22_246; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_246;
  reg [255:0] _T_22_247; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_247;
  reg [255:0] _T_22_248; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_248;
  reg [255:0] _T_22_249; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_249;
  reg [255:0] _T_22_250; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_250;
  reg [255:0] _T_22_251; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_251;
  reg [255:0] _T_22_252; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_252;
  reg [255:0] _T_22_253; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_253;
  reg [255:0] _T_22_254; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_254;
  reg [255:0] _T_22_255; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_255;
  reg [255:0] _T_22_256; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_256;
  reg [255:0] _T_22_257; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_257;
  reg [255:0] _T_22_258; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_258;
  reg [255:0] _T_22_259; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_259;
  reg [255:0] _T_22_260; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_260;
  reg [255:0] _T_22_261; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_261;
  reg [255:0] _T_22_262; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_262;
  reg [255:0] _T_22_263; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_263;
  reg [255:0] _T_22_264; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_264;
  reg [255:0] _T_22_265; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_265;
  reg [255:0] _T_22_266; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_266;
  reg [255:0] _T_22_267; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_267;
  reg [255:0] _T_22_268; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_268;
  reg [255:0] _T_22_269; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_269;
  reg [255:0] _T_22_270; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_270;
  reg [255:0] _T_22_271; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_271;
  reg [255:0] _T_22_272; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_272;
  reg [255:0] _T_22_273; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_273;
  reg [255:0] _T_22_274; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_274;
  reg [255:0] _T_22_275; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_275;
  reg [255:0] _T_22_276; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_276;
  reg [255:0] _T_22_277; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_277;
  reg [255:0] _T_22_278; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_278;
  reg [255:0] _T_22_279; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_279;
  reg [255:0] _T_22_280; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_280;
  reg [255:0] _T_22_281; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_281;
  reg [255:0] _T_22_282; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_282;
  reg [255:0] _T_22_283; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_283;
  reg [255:0] _T_22_284; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_284;
  reg [255:0] _T_22_285; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_285;
  reg [255:0] _T_22_286; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_286;
  reg [255:0] _T_22_287; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_287;
  reg [255:0] _T_22_288; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_288;
  reg [255:0] _T_22_289; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_289;
  reg [255:0] _T_22_290; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_290;
  reg [255:0] _T_22_291; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_291;
  reg [255:0] _T_22_292; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_292;
  reg [255:0] _T_22_293; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_293;
  reg [255:0] _T_22_294; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_294;
  reg [255:0] _T_22_295; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_295;
  reg [255:0] _T_22_296; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_296;
  reg [255:0] _T_22_297; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_297;
  reg [255:0] _T_22_298; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_298;
  reg [255:0] _T_22_299; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_299;
  reg [255:0] _T_22_300; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_300;
  reg [255:0] _T_22_301; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_301;
  reg [255:0] _T_22_302; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_302;
  reg [255:0] _T_22_303; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_303;
  reg [255:0] _T_22_304; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_304;
  reg [255:0] _T_22_305; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_305;
  reg [255:0] _T_22_306; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_306;
  reg [255:0] _T_22_307; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_307;
  reg [255:0] _T_22_308; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_308;
  reg [255:0] _T_22_309; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_309;
  reg [255:0] _T_22_310; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_310;
  reg [255:0] _T_22_311; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_311;
  reg [255:0] _T_22_312; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_312;
  reg [255:0] _T_22_313; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_313;
  reg [255:0] _T_22_314; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_314;
  reg [255:0] _T_22_315; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_315;
  reg [255:0] _T_22_316; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_316;
  reg [255:0] _T_22_317; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_317;
  reg [255:0] _T_22_318; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_318;
  reg [255:0] _T_22_319; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_319;
  reg [255:0] _T_22_320; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_320;
  reg [255:0] _T_22_321; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_321;
  reg [255:0] _T_22_322; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_322;
  reg [255:0] _T_22_323; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_323;
  reg [255:0] _T_22_324; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_324;
  reg [255:0] _T_22_325; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_325;
  reg [255:0] _T_22_326; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_326;
  reg [255:0] _T_22_327; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_327;
  reg [255:0] _T_22_328; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_328;
  reg [255:0] _T_22_329; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_329;
  reg [255:0] _T_22_330; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_330;
  reg [255:0] _T_22_331; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_331;
  reg [255:0] _T_22_332; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_332;
  reg [255:0] _T_22_333; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_333;
  reg [255:0] _T_22_334; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_334;
  reg [255:0] _T_22_335; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_335;
  reg [255:0] _T_22_336; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_336;
  reg [255:0] _T_22_337; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_337;
  reg [255:0] _T_22_338; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_338;
  reg [255:0] _T_22_339; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_339;
  reg [255:0] _T_22_340; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_340;
  reg [255:0] _T_22_341; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_341;
  reg [255:0] _T_22_342; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_342;
  reg [255:0] _T_22_343; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_343;
  reg [255:0] _T_22_344; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_344;
  reg [255:0] _T_22_345; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_345;
  reg [255:0] _T_22_346; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_346;
  reg [255:0] _T_22_347; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_347;
  reg [255:0] _T_22_348; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_348;
  reg [255:0] _T_22_349; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_349;
  reg [255:0] _T_22_350; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_350;
  reg [255:0] _T_22_351; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_351;
  reg [255:0] _T_22_352; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_352;
  reg [255:0] _T_22_353; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_353;
  reg [255:0] _T_22_354; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_354;
  reg [255:0] _T_22_355; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_355;
  reg [255:0] _T_22_356; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_356;
  reg [255:0] _T_22_357; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_357;
  reg [255:0] _T_22_358; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_358;
  reg [255:0] _T_22_359; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_359;
  reg [255:0] _T_22_360; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_360;
  reg [255:0] _T_22_361; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_361;
  reg [255:0] _T_22_362; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_362;
  reg [255:0] _T_22_363; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_363;
  reg [255:0] _T_22_364; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_364;
  reg [255:0] _T_22_365; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_365;
  reg [255:0] _T_22_366; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_366;
  reg [255:0] _T_22_367; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_367;
  reg [255:0] _T_22_368; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_368;
  reg [255:0] _T_22_369; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_369;
  reg [255:0] _T_22_370; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_370;
  reg [255:0] _T_22_371; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_371;
  reg [255:0] _T_22_372; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_372;
  reg [255:0] _T_22_373; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_373;
  reg [255:0] _T_22_374; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_374;
  reg [255:0] _T_22_375; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_375;
  reg [255:0] _T_22_376; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_376;
  reg [255:0] _T_22_377; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_377;
  reg [255:0] _T_22_378; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_378;
  reg [255:0] _T_22_379; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_379;
  reg [255:0] _T_22_380; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_380;
  reg [255:0] _T_22_381; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_381;
  reg [255:0] _T_22_382; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_382;
  reg [255:0] _T_22_383; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_383;
  reg [255:0] _T_22_384; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_384;
  reg [255:0] _T_22_385; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_385;
  reg [255:0] _T_22_386; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_386;
  reg [255:0] _T_22_387; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_387;
  reg [255:0] _T_22_388; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_388;
  reg [255:0] _T_22_389; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_389;
  reg [255:0] _T_22_390; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_390;
  reg [255:0] _T_22_391; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_391;
  reg [255:0] _T_22_392; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_392;
  reg [255:0] _T_22_393; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_393;
  reg [255:0] _T_22_394; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_394;
  reg [255:0] _T_22_395; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_395;
  reg [255:0] _T_22_396; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_396;
  reg [255:0] _T_22_397; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_397;
  reg [255:0] _T_22_398; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_398;
  reg [255:0] _T_22_399; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_399;
  reg [255:0] _T_22_400; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_400;
  reg [255:0] _T_22_401; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_401;
  reg [255:0] _T_22_402; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_402;
  reg [255:0] _T_22_403; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_403;
  reg [255:0] _T_22_404; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_404;
  reg [255:0] _T_22_405; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_405;
  reg [255:0] _T_22_406; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_406;
  reg [255:0] _T_22_407; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_407;
  reg [255:0] _T_22_408; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_408;
  reg [255:0] _T_22_409; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_409;
  reg [255:0] _T_22_410; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_410;
  reg [255:0] _T_22_411; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_411;
  reg [255:0] _T_22_412; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_412;
  reg [255:0] _T_22_413; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_413;
  reg [255:0] _T_22_414; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_414;
  reg [255:0] _T_22_415; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_415;
  reg [255:0] _T_22_416; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_416;
  reg [255:0] _T_22_417; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_417;
  reg [255:0] _T_22_418; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_418;
  reg [255:0] _T_22_419; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_419;
  reg [255:0] _T_22_420; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_420;
  reg [255:0] _T_22_421; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_421;
  reg [255:0] _T_22_422; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_422;
  reg [255:0] _T_22_423; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_423;
  reg [255:0] _T_22_424; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_424;
  reg [255:0] _T_22_425; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_425;
  reg [255:0] _T_22_426; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_426;
  reg [255:0] _T_22_427; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_427;
  reg [255:0] _T_22_428; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_428;
  reg [255:0] _T_22_429; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_429;
  reg [255:0] _T_22_430; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_430;
  reg [255:0] _T_22_431; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_431;
  reg [255:0] _T_22_432; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_432;
  reg [255:0] _T_22_433; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_433;
  reg [255:0] _T_22_434; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_434;
  reg [255:0] _T_22_435; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_435;
  reg [255:0] _T_22_436; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_436;
  reg [255:0] _T_22_437; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_437;
  reg [255:0] _T_22_438; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_438;
  reg [255:0] _T_22_439; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_439;
  reg [255:0] _T_22_440; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_440;
  reg [255:0] _T_22_441; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_441;
  reg [255:0] _T_22_442; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_442;
  reg [255:0] _T_22_443; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_443;
  reg [255:0] _T_22_444; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_444;
  reg [255:0] _T_22_445; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_445;
  reg [255:0] _T_22_446; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_446;
  reg [255:0] _T_22_447; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_447;
  reg [255:0] _T_22_448; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_448;
  reg [255:0] _T_22_449; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_449;
  reg [255:0] _T_22_450; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_450;
  reg [255:0] _T_22_451; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_451;
  reg [255:0] _T_22_452; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_452;
  reg [255:0] _T_22_453; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_453;
  reg [255:0] _T_22_454; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_454;
  reg [255:0] _T_22_455; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_455;
  reg [255:0] _T_22_456; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_456;
  reg [255:0] _T_22_457; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_457;
  reg [255:0] _T_22_458; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_458;
  reg [255:0] _T_22_459; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_459;
  reg [255:0] _T_22_460; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_460;
  reg [255:0] _T_22_461; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_461;
  reg [255:0] _T_22_462; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_462;
  reg [255:0] _T_22_463; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_463;
  reg [255:0] _T_22_464; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_464;
  reg [255:0] _T_22_465; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_465;
  reg [255:0] _T_22_466; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_466;
  reg [255:0] _T_22_467; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_467;
  reg [255:0] _T_22_468; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_468;
  reg [255:0] _T_22_469; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_469;
  reg [255:0] _T_22_470; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_470;
  reg [255:0] _T_22_471; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_471;
  reg [255:0] _T_22_472; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_472;
  reg [255:0] _T_22_473; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_473;
  reg [255:0] _T_22_474; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_474;
  reg [255:0] _T_22_475; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_475;
  reg [255:0] _T_22_476; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_476;
  reg [255:0] _T_22_477; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_477;
  reg [255:0] _T_22_478; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_478;
  reg [255:0] _T_22_479; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_479;
  reg [255:0] _T_22_480; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_480;
  reg [255:0] _T_22_481; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_481;
  reg [255:0] _T_22_482; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_482;
  reg [255:0] _T_22_483; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_483;
  reg [255:0] _T_22_484; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_484;
  reg [255:0] _T_22_485; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_485;
  reg [255:0] _T_22_486; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_486;
  reg [255:0] _T_22_487; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_487;
  reg [255:0] _T_22_488; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_488;
  reg [255:0] _T_22_489; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_489;
  reg [255:0] _T_22_490; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_490;
  reg [255:0] _T_22_491; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_491;
  reg [255:0] _T_22_492; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_492;
  reg [255:0] _T_22_493; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_493;
  reg [255:0] _T_22_494; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_494;
  reg [255:0] _T_22_495; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_495;
  reg [255:0] _T_22_496; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_496;
  reg [255:0] _T_22_497; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_497;
  reg [255:0] _T_22_498; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_498;
  reg [255:0] _T_22_499; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_499;
  reg [255:0] _T_22_500; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_500;
  reg [255:0] _T_22_501; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_501;
  reg [255:0] _T_22_502; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_502;
  reg [255:0] _T_22_503; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_503;
  reg [255:0] _T_22_504; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_504;
  reg [255:0] _T_22_505; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_505;
  reg [255:0] _T_22_506; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_506;
  reg [255:0] _T_22_507; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_507;
  reg [255:0] _T_22_508; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_508;
  reg [255:0] _T_22_509; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_509;
  reg [255:0] _T_22_510; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_510;
  reg [255:0] _T_22_511; // @[nv_ram_rws.scala 27:18:@8.4]
  reg [255:0] _RAND_511;
  reg [8:0] _T_538; // @[nv_ram_rws.scala 28:19:@9.4]
  reg [31:0] _RAND_512;
  wire [255:0] _GEN_0; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_1; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_2; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_3; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_4; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_5; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_6; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_7; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_8; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_9; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_10; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_11; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_12; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_13; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_14; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_15; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_16; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_17; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_18; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_19; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_20; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_21; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_22; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_23; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_24; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_25; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_26; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_27; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_28; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_29; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_30; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_31; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_32; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_33; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_34; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_35; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_36; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_37; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_38; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_39; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_40; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_41; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_42; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_43; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_44; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_45; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_46; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_47; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_48; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_49; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_50; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_51; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_52; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_53; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_54; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_55; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_56; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_57; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_58; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_59; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_60; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_61; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_62; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_63; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_64; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_65; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_66; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_67; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_68; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_69; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_70; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_71; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_72; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_73; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_74; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_75; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_76; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_77; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_78; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_79; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_80; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_81; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_82; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_83; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_84; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_85; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_86; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_87; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_88; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_89; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_90; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_91; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_92; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_93; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_94; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_95; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_96; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_97; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_98; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_99; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_100; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_101; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_102; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_103; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_104; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_105; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_106; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_107; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_108; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_109; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_110; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_111; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_112; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_113; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_114; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_115; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_116; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_117; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_118; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_119; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_120; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_121; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_122; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_123; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_124; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_125; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_126; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_127; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_128; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_129; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_130; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_131; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_132; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_133; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_134; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_135; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_136; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_137; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_138; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_139; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_140; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_141; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_142; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_143; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_144; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_145; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_146; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_147; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_148; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_149; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_150; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_151; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_152; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_153; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_154; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_155; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_156; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_157; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_158; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_159; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_160; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_161; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_162; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_163; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_164; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_165; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_166; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_167; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_168; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_169; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_170; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_171; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_172; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_173; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_174; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_175; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_176; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_177; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_178; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_179; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_180; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_181; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_182; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_183; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_184; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_185; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_186; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_187; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_188; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_189; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_190; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_191; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_192; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_193; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_194; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_195; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_196; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_197; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_198; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_199; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_200; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_201; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_202; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_203; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_204; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_205; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_206; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_207; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_208; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_209; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_210; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_211; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_212; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_213; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_214; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_215; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_216; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_217; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_218; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_219; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_220; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_221; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_222; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_223; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_224; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_225; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_226; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_227; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_228; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_229; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_230; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_231; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_232; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_233; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_234; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_235; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_236; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_237; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_238; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_239; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_240; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_241; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_242; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_243; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_244; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_245; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_246; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_247; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_248; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_249; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_250; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_251; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_252; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_253; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_254; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_255; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_256; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_257; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_258; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_259; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_260; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_261; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_262; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_263; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_264; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_265; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_266; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_267; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_268; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_269; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_270; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_271; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_272; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_273; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_274; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_275; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_276; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_277; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_278; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_279; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_280; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_281; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_282; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_283; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_284; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_285; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_286; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_287; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_288; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_289; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_290; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_291; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_292; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_293; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_294; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_295; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_296; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_297; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_298; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_299; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_300; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_301; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_302; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_303; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_304; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_305; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_306; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_307; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_308; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_309; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_310; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_311; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_312; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_313; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_314; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_315; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_316; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_317; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_318; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_319; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_320; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_321; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_322; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_323; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_324; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_325; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_326; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_327; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_328; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_329; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_330; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_331; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_332; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_333; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_334; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_335; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_336; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_337; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_338; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_339; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_340; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_341; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_342; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_343; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_344; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_345; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_346; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_347; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_348; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_349; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_350; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_351; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_352; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_353; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_354; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_355; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_356; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_357; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_358; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_359; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_360; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_361; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_362; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_363; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_364; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_365; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_366; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_367; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_368; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_369; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_370; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_371; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_372; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_373; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_374; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_375; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_376; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_377; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_378; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_379; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_380; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_381; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_382; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_383; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_384; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_385; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_386; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_387; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_388; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_389; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_390; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_391; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_392; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_393; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_394; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_395; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_396; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_397; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_398; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_399; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_400; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_401; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_402; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_403; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_404; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_405; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_406; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_407; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_408; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_409; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_410; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_411; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_412; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_413; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_414; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_415; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_416; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_417; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_418; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_419; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_420; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_421; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_422; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_423; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_424; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_425; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_426; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_427; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_428; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_429; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_430; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_431; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_432; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_433; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_434; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_435; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_436; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_437; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_438; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_439; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_440; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_441; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_442; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_443; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_444; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_445; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_446; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_447; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_448; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_449; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_450; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_451; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_452; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_453; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_454; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_455; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_456; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_457; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_458; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_459; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_460; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_461; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_462; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_463; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_464; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_465; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_466; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_467; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_468; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_469; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_470; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_471; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_472; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_473; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_474; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_475; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_476; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_477; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_478; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_479; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_480; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_481; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_482; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_483; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_484; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_485; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_486; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_487; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_488; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_489; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_490; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_491; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_492; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_493; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_494; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_495; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_496; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_497; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_498; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_499; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_500; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_501; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_502; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_503; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_504; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_505; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_506; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_507; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_508; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_509; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_510; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_511; // @[nv_ram_rws.scala 31:20:@11.6]
  wire [255:0] _GEN_1026; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1027; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1028; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1029; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1030; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1031; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1032; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1033; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1034; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1035; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1036; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1037; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1038; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1039; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1040; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1041; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1042; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1043; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1044; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1045; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1046; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1047; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1048; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1049; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1050; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1051; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1052; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1053; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1054; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1055; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1056; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1057; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1058; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1059; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1060; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1061; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1062; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1063; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1064; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1065; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1066; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1067; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1068; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1069; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1070; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1071; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1072; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1073; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1074; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1075; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1076; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1077; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1078; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1079; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1080; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1081; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1082; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1083; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1084; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1085; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1086; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1087; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1088; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1089; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1090; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1091; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1092; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1093; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1094; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1095; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1096; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1097; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1098; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1099; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1100; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1101; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1102; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1103; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1104; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1105; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1106; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1107; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1108; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1109; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1110; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1111; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1112; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1113; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1114; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1115; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1116; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1117; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1118; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1119; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1120; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1121; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1122; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1123; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1124; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1125; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1126; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1127; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1128; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1129; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1130; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1131; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1132; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1133; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1134; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1135; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1136; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1137; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1138; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1139; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1140; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1141; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1142; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1143; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1144; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1145; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1146; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1147; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1148; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1149; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1150; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1151; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1152; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1153; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1154; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1155; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1156; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1157; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1158; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1159; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1160; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1161; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1162; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1163; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1164; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1165; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1166; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1167; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1168; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1169; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1170; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1171; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1172; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1173; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1174; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1175; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1176; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1177; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1178; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1179; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1180; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1181; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1182; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1183; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1184; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1185; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1186; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1187; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1188; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1189; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1190; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1191; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1192; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1193; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1194; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1195; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1196; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1197; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1198; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1199; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1200; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1201; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1202; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1203; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1204; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1205; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1206; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1207; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1208; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1209; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1210; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1211; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1212; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1213; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1214; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1215; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1216; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1217; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1218; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1219; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1220; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1221; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1222; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1223; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1224; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1225; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1226; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1227; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1228; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1229; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1230; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1231; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1232; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1233; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1234; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1235; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1236; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1237; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1238; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1239; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1240; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1241; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1242; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1243; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1244; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1245; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1246; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1247; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1248; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1249; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1250; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1251; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1252; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1253; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1254; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1255; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1256; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1257; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1258; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1259; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1260; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1261; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1262; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1263; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1264; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1265; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1266; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1267; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1268; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1269; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1270; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1271; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1272; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1273; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1274; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1275; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1276; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1277; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1278; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1279; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1280; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1281; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1282; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1283; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1284; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1285; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1286; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1287; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1288; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1289; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1290; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1291; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1292; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1293; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1294; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1295; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1296; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1297; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1298; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1299; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1300; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1301; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1302; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1303; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1304; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1305; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1306; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1307; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1308; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1309; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1310; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1311; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1312; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1313; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1314; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1315; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1316; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1317; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1318; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1319; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1320; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1321; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1322; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1323; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1324; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1325; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1326; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1327; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1328; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1329; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1330; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1331; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1332; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1333; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1334; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1335; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1336; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1337; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1338; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1339; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1340; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1341; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1342; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1343; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1344; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1345; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1346; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1347; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1348; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1349; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1350; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1351; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1352; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1353; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1354; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1355; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1356; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1357; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1358; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1359; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1360; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1361; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1362; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1363; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1364; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1365; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1366; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1367; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1368; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1369; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1370; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1371; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1372; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1373; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1374; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1375; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1376; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1377; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1378; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1379; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1380; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1381; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1382; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1383; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1384; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1385; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1386; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1387; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1388; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1389; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1390; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1391; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1392; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1393; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1394; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1395; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1396; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1397; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1398; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1399; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1400; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1401; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1402; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1403; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1404; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1405; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1406; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1407; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1408; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1409; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1410; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1411; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1412; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1413; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1414; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1415; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1416; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1417; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1418; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1419; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1420; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1421; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1422; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1423; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1424; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1425; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1426; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1427; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1428; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1429; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1430; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1431; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1432; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1433; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1434; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1435; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1436; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1437; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1438; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1439; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1440; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1441; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1442; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1443; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1444; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1445; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1446; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1447; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1448; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1449; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1450; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1451; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1452; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1453; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1454; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1455; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1456; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1457; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1458; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1459; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1460; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1461; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1462; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1463; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1464; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1465; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1466; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1467; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1468; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1469; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1470; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1471; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1472; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1473; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1474; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1475; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1476; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1477; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1478; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1479; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1480; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1481; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1482; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1483; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1484; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1485; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1486; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1487; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1488; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1489; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1490; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1491; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1492; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1493; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1494; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1495; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1496; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1497; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1498; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1499; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1500; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1501; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1502; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1503; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1504; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1505; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1506; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1507; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1508; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1509; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1510; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1511; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1512; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1513; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1514; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1515; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1516; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1517; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1518; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1519; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1520; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1521; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1522; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1523; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1524; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1525; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1526; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1527; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1528; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1529; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1530; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1531; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1532; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1533; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1534; // @[nv_ram_rws.scala 36:13:@16.4]
  wire [255:0] _GEN_1535; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_0 = 9'h0 == io_wa ? io_di : _T_22_0; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_1 = 9'h1 == io_wa ? io_di : _T_22_1; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_2 = 9'h2 == io_wa ? io_di : _T_22_2; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_3 = 9'h3 == io_wa ? io_di : _T_22_3; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_4 = 9'h4 == io_wa ? io_di : _T_22_4; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_5 = 9'h5 == io_wa ? io_di : _T_22_5; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_6 = 9'h6 == io_wa ? io_di : _T_22_6; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_7 = 9'h7 == io_wa ? io_di : _T_22_7; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_8 = 9'h8 == io_wa ? io_di : _T_22_8; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_9 = 9'h9 == io_wa ? io_di : _T_22_9; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_10 = 9'ha == io_wa ? io_di : _T_22_10; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_11 = 9'hb == io_wa ? io_di : _T_22_11; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_12 = 9'hc == io_wa ? io_di : _T_22_12; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_13 = 9'hd == io_wa ? io_di : _T_22_13; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_14 = 9'he == io_wa ? io_di : _T_22_14; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_15 = 9'hf == io_wa ? io_di : _T_22_15; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_16 = 9'h10 == io_wa ? io_di : _T_22_16; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_17 = 9'h11 == io_wa ? io_di : _T_22_17; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_18 = 9'h12 == io_wa ? io_di : _T_22_18; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_19 = 9'h13 == io_wa ? io_di : _T_22_19; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_20 = 9'h14 == io_wa ? io_di : _T_22_20; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_21 = 9'h15 == io_wa ? io_di : _T_22_21; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_22 = 9'h16 == io_wa ? io_di : _T_22_22; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_23 = 9'h17 == io_wa ? io_di : _T_22_23; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_24 = 9'h18 == io_wa ? io_di : _T_22_24; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_25 = 9'h19 == io_wa ? io_di : _T_22_25; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_26 = 9'h1a == io_wa ? io_di : _T_22_26; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_27 = 9'h1b == io_wa ? io_di : _T_22_27; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_28 = 9'h1c == io_wa ? io_di : _T_22_28; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_29 = 9'h1d == io_wa ? io_di : _T_22_29; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_30 = 9'h1e == io_wa ? io_di : _T_22_30; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_31 = 9'h1f == io_wa ? io_di : _T_22_31; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_32 = 9'h20 == io_wa ? io_di : _T_22_32; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_33 = 9'h21 == io_wa ? io_di : _T_22_33; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_34 = 9'h22 == io_wa ? io_di : _T_22_34; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_35 = 9'h23 == io_wa ? io_di : _T_22_35; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_36 = 9'h24 == io_wa ? io_di : _T_22_36; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_37 = 9'h25 == io_wa ? io_di : _T_22_37; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_38 = 9'h26 == io_wa ? io_di : _T_22_38; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_39 = 9'h27 == io_wa ? io_di : _T_22_39; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_40 = 9'h28 == io_wa ? io_di : _T_22_40; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_41 = 9'h29 == io_wa ? io_di : _T_22_41; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_42 = 9'h2a == io_wa ? io_di : _T_22_42; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_43 = 9'h2b == io_wa ? io_di : _T_22_43; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_44 = 9'h2c == io_wa ? io_di : _T_22_44; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_45 = 9'h2d == io_wa ? io_di : _T_22_45; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_46 = 9'h2e == io_wa ? io_di : _T_22_46; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_47 = 9'h2f == io_wa ? io_di : _T_22_47; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_48 = 9'h30 == io_wa ? io_di : _T_22_48; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_49 = 9'h31 == io_wa ? io_di : _T_22_49; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_50 = 9'h32 == io_wa ? io_di : _T_22_50; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_51 = 9'h33 == io_wa ? io_di : _T_22_51; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_52 = 9'h34 == io_wa ? io_di : _T_22_52; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_53 = 9'h35 == io_wa ? io_di : _T_22_53; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_54 = 9'h36 == io_wa ? io_di : _T_22_54; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_55 = 9'h37 == io_wa ? io_di : _T_22_55; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_56 = 9'h38 == io_wa ? io_di : _T_22_56; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_57 = 9'h39 == io_wa ? io_di : _T_22_57; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_58 = 9'h3a == io_wa ? io_di : _T_22_58; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_59 = 9'h3b == io_wa ? io_di : _T_22_59; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_60 = 9'h3c == io_wa ? io_di : _T_22_60; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_61 = 9'h3d == io_wa ? io_di : _T_22_61; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_62 = 9'h3e == io_wa ? io_di : _T_22_62; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_63 = 9'h3f == io_wa ? io_di : _T_22_63; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_64 = 9'h40 == io_wa ? io_di : _T_22_64; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_65 = 9'h41 == io_wa ? io_di : _T_22_65; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_66 = 9'h42 == io_wa ? io_di : _T_22_66; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_67 = 9'h43 == io_wa ? io_di : _T_22_67; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_68 = 9'h44 == io_wa ? io_di : _T_22_68; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_69 = 9'h45 == io_wa ? io_di : _T_22_69; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_70 = 9'h46 == io_wa ? io_di : _T_22_70; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_71 = 9'h47 == io_wa ? io_di : _T_22_71; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_72 = 9'h48 == io_wa ? io_di : _T_22_72; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_73 = 9'h49 == io_wa ? io_di : _T_22_73; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_74 = 9'h4a == io_wa ? io_di : _T_22_74; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_75 = 9'h4b == io_wa ? io_di : _T_22_75; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_76 = 9'h4c == io_wa ? io_di : _T_22_76; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_77 = 9'h4d == io_wa ? io_di : _T_22_77; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_78 = 9'h4e == io_wa ? io_di : _T_22_78; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_79 = 9'h4f == io_wa ? io_di : _T_22_79; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_80 = 9'h50 == io_wa ? io_di : _T_22_80; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_81 = 9'h51 == io_wa ? io_di : _T_22_81; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_82 = 9'h52 == io_wa ? io_di : _T_22_82; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_83 = 9'h53 == io_wa ? io_di : _T_22_83; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_84 = 9'h54 == io_wa ? io_di : _T_22_84; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_85 = 9'h55 == io_wa ? io_di : _T_22_85; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_86 = 9'h56 == io_wa ? io_di : _T_22_86; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_87 = 9'h57 == io_wa ? io_di : _T_22_87; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_88 = 9'h58 == io_wa ? io_di : _T_22_88; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_89 = 9'h59 == io_wa ? io_di : _T_22_89; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_90 = 9'h5a == io_wa ? io_di : _T_22_90; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_91 = 9'h5b == io_wa ? io_di : _T_22_91; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_92 = 9'h5c == io_wa ? io_di : _T_22_92; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_93 = 9'h5d == io_wa ? io_di : _T_22_93; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_94 = 9'h5e == io_wa ? io_di : _T_22_94; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_95 = 9'h5f == io_wa ? io_di : _T_22_95; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_96 = 9'h60 == io_wa ? io_di : _T_22_96; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_97 = 9'h61 == io_wa ? io_di : _T_22_97; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_98 = 9'h62 == io_wa ? io_di : _T_22_98; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_99 = 9'h63 == io_wa ? io_di : _T_22_99; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_100 = 9'h64 == io_wa ? io_di : _T_22_100; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_101 = 9'h65 == io_wa ? io_di : _T_22_101; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_102 = 9'h66 == io_wa ? io_di : _T_22_102; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_103 = 9'h67 == io_wa ? io_di : _T_22_103; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_104 = 9'h68 == io_wa ? io_di : _T_22_104; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_105 = 9'h69 == io_wa ? io_di : _T_22_105; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_106 = 9'h6a == io_wa ? io_di : _T_22_106; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_107 = 9'h6b == io_wa ? io_di : _T_22_107; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_108 = 9'h6c == io_wa ? io_di : _T_22_108; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_109 = 9'h6d == io_wa ? io_di : _T_22_109; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_110 = 9'h6e == io_wa ? io_di : _T_22_110; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_111 = 9'h6f == io_wa ? io_di : _T_22_111; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_112 = 9'h70 == io_wa ? io_di : _T_22_112; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_113 = 9'h71 == io_wa ? io_di : _T_22_113; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_114 = 9'h72 == io_wa ? io_di : _T_22_114; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_115 = 9'h73 == io_wa ? io_di : _T_22_115; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_116 = 9'h74 == io_wa ? io_di : _T_22_116; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_117 = 9'h75 == io_wa ? io_di : _T_22_117; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_118 = 9'h76 == io_wa ? io_di : _T_22_118; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_119 = 9'h77 == io_wa ? io_di : _T_22_119; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_120 = 9'h78 == io_wa ? io_di : _T_22_120; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_121 = 9'h79 == io_wa ? io_di : _T_22_121; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_122 = 9'h7a == io_wa ? io_di : _T_22_122; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_123 = 9'h7b == io_wa ? io_di : _T_22_123; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_124 = 9'h7c == io_wa ? io_di : _T_22_124; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_125 = 9'h7d == io_wa ? io_di : _T_22_125; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_126 = 9'h7e == io_wa ? io_di : _T_22_126; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_127 = 9'h7f == io_wa ? io_di : _T_22_127; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_128 = 9'h80 == io_wa ? io_di : _T_22_128; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_129 = 9'h81 == io_wa ? io_di : _T_22_129; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_130 = 9'h82 == io_wa ? io_di : _T_22_130; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_131 = 9'h83 == io_wa ? io_di : _T_22_131; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_132 = 9'h84 == io_wa ? io_di : _T_22_132; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_133 = 9'h85 == io_wa ? io_di : _T_22_133; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_134 = 9'h86 == io_wa ? io_di : _T_22_134; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_135 = 9'h87 == io_wa ? io_di : _T_22_135; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_136 = 9'h88 == io_wa ? io_di : _T_22_136; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_137 = 9'h89 == io_wa ? io_di : _T_22_137; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_138 = 9'h8a == io_wa ? io_di : _T_22_138; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_139 = 9'h8b == io_wa ? io_di : _T_22_139; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_140 = 9'h8c == io_wa ? io_di : _T_22_140; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_141 = 9'h8d == io_wa ? io_di : _T_22_141; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_142 = 9'h8e == io_wa ? io_di : _T_22_142; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_143 = 9'h8f == io_wa ? io_di : _T_22_143; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_144 = 9'h90 == io_wa ? io_di : _T_22_144; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_145 = 9'h91 == io_wa ? io_di : _T_22_145; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_146 = 9'h92 == io_wa ? io_di : _T_22_146; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_147 = 9'h93 == io_wa ? io_di : _T_22_147; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_148 = 9'h94 == io_wa ? io_di : _T_22_148; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_149 = 9'h95 == io_wa ? io_di : _T_22_149; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_150 = 9'h96 == io_wa ? io_di : _T_22_150; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_151 = 9'h97 == io_wa ? io_di : _T_22_151; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_152 = 9'h98 == io_wa ? io_di : _T_22_152; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_153 = 9'h99 == io_wa ? io_di : _T_22_153; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_154 = 9'h9a == io_wa ? io_di : _T_22_154; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_155 = 9'h9b == io_wa ? io_di : _T_22_155; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_156 = 9'h9c == io_wa ? io_di : _T_22_156; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_157 = 9'h9d == io_wa ? io_di : _T_22_157; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_158 = 9'h9e == io_wa ? io_di : _T_22_158; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_159 = 9'h9f == io_wa ? io_di : _T_22_159; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_160 = 9'ha0 == io_wa ? io_di : _T_22_160; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_161 = 9'ha1 == io_wa ? io_di : _T_22_161; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_162 = 9'ha2 == io_wa ? io_di : _T_22_162; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_163 = 9'ha3 == io_wa ? io_di : _T_22_163; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_164 = 9'ha4 == io_wa ? io_di : _T_22_164; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_165 = 9'ha5 == io_wa ? io_di : _T_22_165; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_166 = 9'ha6 == io_wa ? io_di : _T_22_166; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_167 = 9'ha7 == io_wa ? io_di : _T_22_167; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_168 = 9'ha8 == io_wa ? io_di : _T_22_168; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_169 = 9'ha9 == io_wa ? io_di : _T_22_169; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_170 = 9'haa == io_wa ? io_di : _T_22_170; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_171 = 9'hab == io_wa ? io_di : _T_22_171; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_172 = 9'hac == io_wa ? io_di : _T_22_172; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_173 = 9'had == io_wa ? io_di : _T_22_173; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_174 = 9'hae == io_wa ? io_di : _T_22_174; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_175 = 9'haf == io_wa ? io_di : _T_22_175; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_176 = 9'hb0 == io_wa ? io_di : _T_22_176; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_177 = 9'hb1 == io_wa ? io_di : _T_22_177; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_178 = 9'hb2 == io_wa ? io_di : _T_22_178; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_179 = 9'hb3 == io_wa ? io_di : _T_22_179; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_180 = 9'hb4 == io_wa ? io_di : _T_22_180; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_181 = 9'hb5 == io_wa ? io_di : _T_22_181; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_182 = 9'hb6 == io_wa ? io_di : _T_22_182; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_183 = 9'hb7 == io_wa ? io_di : _T_22_183; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_184 = 9'hb8 == io_wa ? io_di : _T_22_184; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_185 = 9'hb9 == io_wa ? io_di : _T_22_185; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_186 = 9'hba == io_wa ? io_di : _T_22_186; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_187 = 9'hbb == io_wa ? io_di : _T_22_187; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_188 = 9'hbc == io_wa ? io_di : _T_22_188; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_189 = 9'hbd == io_wa ? io_di : _T_22_189; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_190 = 9'hbe == io_wa ? io_di : _T_22_190; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_191 = 9'hbf == io_wa ? io_di : _T_22_191; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_192 = 9'hc0 == io_wa ? io_di : _T_22_192; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_193 = 9'hc1 == io_wa ? io_di : _T_22_193; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_194 = 9'hc2 == io_wa ? io_di : _T_22_194; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_195 = 9'hc3 == io_wa ? io_di : _T_22_195; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_196 = 9'hc4 == io_wa ? io_di : _T_22_196; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_197 = 9'hc5 == io_wa ? io_di : _T_22_197; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_198 = 9'hc6 == io_wa ? io_di : _T_22_198; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_199 = 9'hc7 == io_wa ? io_di : _T_22_199; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_200 = 9'hc8 == io_wa ? io_di : _T_22_200; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_201 = 9'hc9 == io_wa ? io_di : _T_22_201; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_202 = 9'hca == io_wa ? io_di : _T_22_202; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_203 = 9'hcb == io_wa ? io_di : _T_22_203; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_204 = 9'hcc == io_wa ? io_di : _T_22_204; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_205 = 9'hcd == io_wa ? io_di : _T_22_205; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_206 = 9'hce == io_wa ? io_di : _T_22_206; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_207 = 9'hcf == io_wa ? io_di : _T_22_207; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_208 = 9'hd0 == io_wa ? io_di : _T_22_208; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_209 = 9'hd1 == io_wa ? io_di : _T_22_209; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_210 = 9'hd2 == io_wa ? io_di : _T_22_210; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_211 = 9'hd3 == io_wa ? io_di : _T_22_211; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_212 = 9'hd4 == io_wa ? io_di : _T_22_212; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_213 = 9'hd5 == io_wa ? io_di : _T_22_213; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_214 = 9'hd6 == io_wa ? io_di : _T_22_214; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_215 = 9'hd7 == io_wa ? io_di : _T_22_215; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_216 = 9'hd8 == io_wa ? io_di : _T_22_216; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_217 = 9'hd9 == io_wa ? io_di : _T_22_217; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_218 = 9'hda == io_wa ? io_di : _T_22_218; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_219 = 9'hdb == io_wa ? io_di : _T_22_219; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_220 = 9'hdc == io_wa ? io_di : _T_22_220; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_221 = 9'hdd == io_wa ? io_di : _T_22_221; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_222 = 9'hde == io_wa ? io_di : _T_22_222; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_223 = 9'hdf == io_wa ? io_di : _T_22_223; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_224 = 9'he0 == io_wa ? io_di : _T_22_224; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_225 = 9'he1 == io_wa ? io_di : _T_22_225; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_226 = 9'he2 == io_wa ? io_di : _T_22_226; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_227 = 9'he3 == io_wa ? io_di : _T_22_227; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_228 = 9'he4 == io_wa ? io_di : _T_22_228; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_229 = 9'he5 == io_wa ? io_di : _T_22_229; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_230 = 9'he6 == io_wa ? io_di : _T_22_230; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_231 = 9'he7 == io_wa ? io_di : _T_22_231; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_232 = 9'he8 == io_wa ? io_di : _T_22_232; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_233 = 9'he9 == io_wa ? io_di : _T_22_233; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_234 = 9'hea == io_wa ? io_di : _T_22_234; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_235 = 9'heb == io_wa ? io_di : _T_22_235; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_236 = 9'hec == io_wa ? io_di : _T_22_236; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_237 = 9'hed == io_wa ? io_di : _T_22_237; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_238 = 9'hee == io_wa ? io_di : _T_22_238; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_239 = 9'hef == io_wa ? io_di : _T_22_239; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_240 = 9'hf0 == io_wa ? io_di : _T_22_240; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_241 = 9'hf1 == io_wa ? io_di : _T_22_241; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_242 = 9'hf2 == io_wa ? io_di : _T_22_242; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_243 = 9'hf3 == io_wa ? io_di : _T_22_243; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_244 = 9'hf4 == io_wa ? io_di : _T_22_244; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_245 = 9'hf5 == io_wa ? io_di : _T_22_245; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_246 = 9'hf6 == io_wa ? io_di : _T_22_246; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_247 = 9'hf7 == io_wa ? io_di : _T_22_247; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_248 = 9'hf8 == io_wa ? io_di : _T_22_248; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_249 = 9'hf9 == io_wa ? io_di : _T_22_249; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_250 = 9'hfa == io_wa ? io_di : _T_22_250; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_251 = 9'hfb == io_wa ? io_di : _T_22_251; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_252 = 9'hfc == io_wa ? io_di : _T_22_252; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_253 = 9'hfd == io_wa ? io_di : _T_22_253; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_254 = 9'hfe == io_wa ? io_di : _T_22_254; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_255 = 9'hff == io_wa ? io_di : _T_22_255; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_256 = 9'h100 == io_wa ? io_di : _T_22_256; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_257 = 9'h101 == io_wa ? io_di : _T_22_257; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_258 = 9'h102 == io_wa ? io_di : _T_22_258; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_259 = 9'h103 == io_wa ? io_di : _T_22_259; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_260 = 9'h104 == io_wa ? io_di : _T_22_260; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_261 = 9'h105 == io_wa ? io_di : _T_22_261; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_262 = 9'h106 == io_wa ? io_di : _T_22_262; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_263 = 9'h107 == io_wa ? io_di : _T_22_263; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_264 = 9'h108 == io_wa ? io_di : _T_22_264; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_265 = 9'h109 == io_wa ? io_di : _T_22_265; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_266 = 9'h10a == io_wa ? io_di : _T_22_266; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_267 = 9'h10b == io_wa ? io_di : _T_22_267; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_268 = 9'h10c == io_wa ? io_di : _T_22_268; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_269 = 9'h10d == io_wa ? io_di : _T_22_269; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_270 = 9'h10e == io_wa ? io_di : _T_22_270; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_271 = 9'h10f == io_wa ? io_di : _T_22_271; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_272 = 9'h110 == io_wa ? io_di : _T_22_272; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_273 = 9'h111 == io_wa ? io_di : _T_22_273; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_274 = 9'h112 == io_wa ? io_di : _T_22_274; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_275 = 9'h113 == io_wa ? io_di : _T_22_275; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_276 = 9'h114 == io_wa ? io_di : _T_22_276; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_277 = 9'h115 == io_wa ? io_di : _T_22_277; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_278 = 9'h116 == io_wa ? io_di : _T_22_278; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_279 = 9'h117 == io_wa ? io_di : _T_22_279; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_280 = 9'h118 == io_wa ? io_di : _T_22_280; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_281 = 9'h119 == io_wa ? io_di : _T_22_281; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_282 = 9'h11a == io_wa ? io_di : _T_22_282; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_283 = 9'h11b == io_wa ? io_di : _T_22_283; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_284 = 9'h11c == io_wa ? io_di : _T_22_284; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_285 = 9'h11d == io_wa ? io_di : _T_22_285; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_286 = 9'h11e == io_wa ? io_di : _T_22_286; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_287 = 9'h11f == io_wa ? io_di : _T_22_287; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_288 = 9'h120 == io_wa ? io_di : _T_22_288; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_289 = 9'h121 == io_wa ? io_di : _T_22_289; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_290 = 9'h122 == io_wa ? io_di : _T_22_290; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_291 = 9'h123 == io_wa ? io_di : _T_22_291; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_292 = 9'h124 == io_wa ? io_di : _T_22_292; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_293 = 9'h125 == io_wa ? io_di : _T_22_293; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_294 = 9'h126 == io_wa ? io_di : _T_22_294; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_295 = 9'h127 == io_wa ? io_di : _T_22_295; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_296 = 9'h128 == io_wa ? io_di : _T_22_296; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_297 = 9'h129 == io_wa ? io_di : _T_22_297; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_298 = 9'h12a == io_wa ? io_di : _T_22_298; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_299 = 9'h12b == io_wa ? io_di : _T_22_299; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_300 = 9'h12c == io_wa ? io_di : _T_22_300; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_301 = 9'h12d == io_wa ? io_di : _T_22_301; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_302 = 9'h12e == io_wa ? io_di : _T_22_302; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_303 = 9'h12f == io_wa ? io_di : _T_22_303; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_304 = 9'h130 == io_wa ? io_di : _T_22_304; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_305 = 9'h131 == io_wa ? io_di : _T_22_305; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_306 = 9'h132 == io_wa ? io_di : _T_22_306; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_307 = 9'h133 == io_wa ? io_di : _T_22_307; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_308 = 9'h134 == io_wa ? io_di : _T_22_308; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_309 = 9'h135 == io_wa ? io_di : _T_22_309; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_310 = 9'h136 == io_wa ? io_di : _T_22_310; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_311 = 9'h137 == io_wa ? io_di : _T_22_311; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_312 = 9'h138 == io_wa ? io_di : _T_22_312; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_313 = 9'h139 == io_wa ? io_di : _T_22_313; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_314 = 9'h13a == io_wa ? io_di : _T_22_314; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_315 = 9'h13b == io_wa ? io_di : _T_22_315; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_316 = 9'h13c == io_wa ? io_di : _T_22_316; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_317 = 9'h13d == io_wa ? io_di : _T_22_317; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_318 = 9'h13e == io_wa ? io_di : _T_22_318; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_319 = 9'h13f == io_wa ? io_di : _T_22_319; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_320 = 9'h140 == io_wa ? io_di : _T_22_320; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_321 = 9'h141 == io_wa ? io_di : _T_22_321; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_322 = 9'h142 == io_wa ? io_di : _T_22_322; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_323 = 9'h143 == io_wa ? io_di : _T_22_323; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_324 = 9'h144 == io_wa ? io_di : _T_22_324; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_325 = 9'h145 == io_wa ? io_di : _T_22_325; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_326 = 9'h146 == io_wa ? io_di : _T_22_326; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_327 = 9'h147 == io_wa ? io_di : _T_22_327; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_328 = 9'h148 == io_wa ? io_di : _T_22_328; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_329 = 9'h149 == io_wa ? io_di : _T_22_329; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_330 = 9'h14a == io_wa ? io_di : _T_22_330; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_331 = 9'h14b == io_wa ? io_di : _T_22_331; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_332 = 9'h14c == io_wa ? io_di : _T_22_332; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_333 = 9'h14d == io_wa ? io_di : _T_22_333; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_334 = 9'h14e == io_wa ? io_di : _T_22_334; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_335 = 9'h14f == io_wa ? io_di : _T_22_335; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_336 = 9'h150 == io_wa ? io_di : _T_22_336; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_337 = 9'h151 == io_wa ? io_di : _T_22_337; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_338 = 9'h152 == io_wa ? io_di : _T_22_338; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_339 = 9'h153 == io_wa ? io_di : _T_22_339; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_340 = 9'h154 == io_wa ? io_di : _T_22_340; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_341 = 9'h155 == io_wa ? io_di : _T_22_341; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_342 = 9'h156 == io_wa ? io_di : _T_22_342; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_343 = 9'h157 == io_wa ? io_di : _T_22_343; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_344 = 9'h158 == io_wa ? io_di : _T_22_344; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_345 = 9'h159 == io_wa ? io_di : _T_22_345; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_346 = 9'h15a == io_wa ? io_di : _T_22_346; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_347 = 9'h15b == io_wa ? io_di : _T_22_347; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_348 = 9'h15c == io_wa ? io_di : _T_22_348; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_349 = 9'h15d == io_wa ? io_di : _T_22_349; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_350 = 9'h15e == io_wa ? io_di : _T_22_350; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_351 = 9'h15f == io_wa ? io_di : _T_22_351; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_352 = 9'h160 == io_wa ? io_di : _T_22_352; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_353 = 9'h161 == io_wa ? io_di : _T_22_353; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_354 = 9'h162 == io_wa ? io_di : _T_22_354; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_355 = 9'h163 == io_wa ? io_di : _T_22_355; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_356 = 9'h164 == io_wa ? io_di : _T_22_356; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_357 = 9'h165 == io_wa ? io_di : _T_22_357; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_358 = 9'h166 == io_wa ? io_di : _T_22_358; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_359 = 9'h167 == io_wa ? io_di : _T_22_359; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_360 = 9'h168 == io_wa ? io_di : _T_22_360; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_361 = 9'h169 == io_wa ? io_di : _T_22_361; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_362 = 9'h16a == io_wa ? io_di : _T_22_362; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_363 = 9'h16b == io_wa ? io_di : _T_22_363; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_364 = 9'h16c == io_wa ? io_di : _T_22_364; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_365 = 9'h16d == io_wa ? io_di : _T_22_365; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_366 = 9'h16e == io_wa ? io_di : _T_22_366; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_367 = 9'h16f == io_wa ? io_di : _T_22_367; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_368 = 9'h170 == io_wa ? io_di : _T_22_368; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_369 = 9'h171 == io_wa ? io_di : _T_22_369; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_370 = 9'h172 == io_wa ? io_di : _T_22_370; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_371 = 9'h173 == io_wa ? io_di : _T_22_371; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_372 = 9'h174 == io_wa ? io_di : _T_22_372; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_373 = 9'h175 == io_wa ? io_di : _T_22_373; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_374 = 9'h176 == io_wa ? io_di : _T_22_374; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_375 = 9'h177 == io_wa ? io_di : _T_22_375; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_376 = 9'h178 == io_wa ? io_di : _T_22_376; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_377 = 9'h179 == io_wa ? io_di : _T_22_377; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_378 = 9'h17a == io_wa ? io_di : _T_22_378; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_379 = 9'h17b == io_wa ? io_di : _T_22_379; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_380 = 9'h17c == io_wa ? io_di : _T_22_380; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_381 = 9'h17d == io_wa ? io_di : _T_22_381; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_382 = 9'h17e == io_wa ? io_di : _T_22_382; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_383 = 9'h17f == io_wa ? io_di : _T_22_383; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_384 = 9'h180 == io_wa ? io_di : _T_22_384; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_385 = 9'h181 == io_wa ? io_di : _T_22_385; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_386 = 9'h182 == io_wa ? io_di : _T_22_386; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_387 = 9'h183 == io_wa ? io_di : _T_22_387; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_388 = 9'h184 == io_wa ? io_di : _T_22_388; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_389 = 9'h185 == io_wa ? io_di : _T_22_389; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_390 = 9'h186 == io_wa ? io_di : _T_22_390; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_391 = 9'h187 == io_wa ? io_di : _T_22_391; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_392 = 9'h188 == io_wa ? io_di : _T_22_392; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_393 = 9'h189 == io_wa ? io_di : _T_22_393; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_394 = 9'h18a == io_wa ? io_di : _T_22_394; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_395 = 9'h18b == io_wa ? io_di : _T_22_395; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_396 = 9'h18c == io_wa ? io_di : _T_22_396; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_397 = 9'h18d == io_wa ? io_di : _T_22_397; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_398 = 9'h18e == io_wa ? io_di : _T_22_398; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_399 = 9'h18f == io_wa ? io_di : _T_22_399; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_400 = 9'h190 == io_wa ? io_di : _T_22_400; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_401 = 9'h191 == io_wa ? io_di : _T_22_401; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_402 = 9'h192 == io_wa ? io_di : _T_22_402; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_403 = 9'h193 == io_wa ? io_di : _T_22_403; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_404 = 9'h194 == io_wa ? io_di : _T_22_404; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_405 = 9'h195 == io_wa ? io_di : _T_22_405; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_406 = 9'h196 == io_wa ? io_di : _T_22_406; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_407 = 9'h197 == io_wa ? io_di : _T_22_407; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_408 = 9'h198 == io_wa ? io_di : _T_22_408; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_409 = 9'h199 == io_wa ? io_di : _T_22_409; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_410 = 9'h19a == io_wa ? io_di : _T_22_410; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_411 = 9'h19b == io_wa ? io_di : _T_22_411; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_412 = 9'h19c == io_wa ? io_di : _T_22_412; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_413 = 9'h19d == io_wa ? io_di : _T_22_413; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_414 = 9'h19e == io_wa ? io_di : _T_22_414; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_415 = 9'h19f == io_wa ? io_di : _T_22_415; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_416 = 9'h1a0 == io_wa ? io_di : _T_22_416; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_417 = 9'h1a1 == io_wa ? io_di : _T_22_417; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_418 = 9'h1a2 == io_wa ? io_di : _T_22_418; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_419 = 9'h1a3 == io_wa ? io_di : _T_22_419; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_420 = 9'h1a4 == io_wa ? io_di : _T_22_420; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_421 = 9'h1a5 == io_wa ? io_di : _T_22_421; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_422 = 9'h1a6 == io_wa ? io_di : _T_22_422; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_423 = 9'h1a7 == io_wa ? io_di : _T_22_423; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_424 = 9'h1a8 == io_wa ? io_di : _T_22_424; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_425 = 9'h1a9 == io_wa ? io_di : _T_22_425; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_426 = 9'h1aa == io_wa ? io_di : _T_22_426; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_427 = 9'h1ab == io_wa ? io_di : _T_22_427; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_428 = 9'h1ac == io_wa ? io_di : _T_22_428; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_429 = 9'h1ad == io_wa ? io_di : _T_22_429; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_430 = 9'h1ae == io_wa ? io_di : _T_22_430; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_431 = 9'h1af == io_wa ? io_di : _T_22_431; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_432 = 9'h1b0 == io_wa ? io_di : _T_22_432; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_433 = 9'h1b1 == io_wa ? io_di : _T_22_433; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_434 = 9'h1b2 == io_wa ? io_di : _T_22_434; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_435 = 9'h1b3 == io_wa ? io_di : _T_22_435; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_436 = 9'h1b4 == io_wa ? io_di : _T_22_436; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_437 = 9'h1b5 == io_wa ? io_di : _T_22_437; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_438 = 9'h1b6 == io_wa ? io_di : _T_22_438; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_439 = 9'h1b7 == io_wa ? io_di : _T_22_439; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_440 = 9'h1b8 == io_wa ? io_di : _T_22_440; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_441 = 9'h1b9 == io_wa ? io_di : _T_22_441; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_442 = 9'h1ba == io_wa ? io_di : _T_22_442; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_443 = 9'h1bb == io_wa ? io_di : _T_22_443; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_444 = 9'h1bc == io_wa ? io_di : _T_22_444; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_445 = 9'h1bd == io_wa ? io_di : _T_22_445; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_446 = 9'h1be == io_wa ? io_di : _T_22_446; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_447 = 9'h1bf == io_wa ? io_di : _T_22_447; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_448 = 9'h1c0 == io_wa ? io_di : _T_22_448; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_449 = 9'h1c1 == io_wa ? io_di : _T_22_449; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_450 = 9'h1c2 == io_wa ? io_di : _T_22_450; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_451 = 9'h1c3 == io_wa ? io_di : _T_22_451; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_452 = 9'h1c4 == io_wa ? io_di : _T_22_452; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_453 = 9'h1c5 == io_wa ? io_di : _T_22_453; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_454 = 9'h1c6 == io_wa ? io_di : _T_22_454; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_455 = 9'h1c7 == io_wa ? io_di : _T_22_455; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_456 = 9'h1c8 == io_wa ? io_di : _T_22_456; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_457 = 9'h1c9 == io_wa ? io_di : _T_22_457; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_458 = 9'h1ca == io_wa ? io_di : _T_22_458; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_459 = 9'h1cb == io_wa ? io_di : _T_22_459; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_460 = 9'h1cc == io_wa ? io_di : _T_22_460; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_461 = 9'h1cd == io_wa ? io_di : _T_22_461; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_462 = 9'h1ce == io_wa ? io_di : _T_22_462; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_463 = 9'h1cf == io_wa ? io_di : _T_22_463; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_464 = 9'h1d0 == io_wa ? io_di : _T_22_464; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_465 = 9'h1d1 == io_wa ? io_di : _T_22_465; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_466 = 9'h1d2 == io_wa ? io_di : _T_22_466; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_467 = 9'h1d3 == io_wa ? io_di : _T_22_467; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_468 = 9'h1d4 == io_wa ? io_di : _T_22_468; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_469 = 9'h1d5 == io_wa ? io_di : _T_22_469; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_470 = 9'h1d6 == io_wa ? io_di : _T_22_470; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_471 = 9'h1d7 == io_wa ? io_di : _T_22_471; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_472 = 9'h1d8 == io_wa ? io_di : _T_22_472; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_473 = 9'h1d9 == io_wa ? io_di : _T_22_473; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_474 = 9'h1da == io_wa ? io_di : _T_22_474; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_475 = 9'h1db == io_wa ? io_di : _T_22_475; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_476 = 9'h1dc == io_wa ? io_di : _T_22_476; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_477 = 9'h1dd == io_wa ? io_di : _T_22_477; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_478 = 9'h1de == io_wa ? io_di : _T_22_478; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_479 = 9'h1df == io_wa ? io_di : _T_22_479; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_480 = 9'h1e0 == io_wa ? io_di : _T_22_480; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_481 = 9'h1e1 == io_wa ? io_di : _T_22_481; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_482 = 9'h1e2 == io_wa ? io_di : _T_22_482; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_483 = 9'h1e3 == io_wa ? io_di : _T_22_483; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_484 = 9'h1e4 == io_wa ? io_di : _T_22_484; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_485 = 9'h1e5 == io_wa ? io_di : _T_22_485; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_486 = 9'h1e6 == io_wa ? io_di : _T_22_486; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_487 = 9'h1e7 == io_wa ? io_di : _T_22_487; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_488 = 9'h1e8 == io_wa ? io_di : _T_22_488; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_489 = 9'h1e9 == io_wa ? io_di : _T_22_489; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_490 = 9'h1ea == io_wa ? io_di : _T_22_490; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_491 = 9'h1eb == io_wa ? io_di : _T_22_491; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_492 = 9'h1ec == io_wa ? io_di : _T_22_492; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_493 = 9'h1ed == io_wa ? io_di : _T_22_493; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_494 = 9'h1ee == io_wa ? io_di : _T_22_494; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_495 = 9'h1ef == io_wa ? io_di : _T_22_495; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_496 = 9'h1f0 == io_wa ? io_di : _T_22_496; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_497 = 9'h1f1 == io_wa ? io_di : _T_22_497; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_498 = 9'h1f2 == io_wa ? io_di : _T_22_498; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_499 = 9'h1f3 == io_wa ? io_di : _T_22_499; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_500 = 9'h1f4 == io_wa ? io_di : _T_22_500; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_501 = 9'h1f5 == io_wa ? io_di : _T_22_501; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_502 = 9'h1f6 == io_wa ? io_di : _T_22_502; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_503 = 9'h1f7 == io_wa ? io_di : _T_22_503; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_504 = 9'h1f8 == io_wa ? io_di : _T_22_504; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_505 = 9'h1f9 == io_wa ? io_di : _T_22_505; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_506 = 9'h1fa == io_wa ? io_di : _T_22_506; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_507 = 9'h1fb == io_wa ? io_di : _T_22_507; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_508 = 9'h1fc == io_wa ? io_di : _T_22_508; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_509 = 9'h1fd == io_wa ? io_di : _T_22_509; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_510 = 9'h1fe == io_wa ? io_di : _T_22_510; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_511 = 9'h1ff == io_wa ? io_di : _T_22_511; // @[nv_ram_rws.scala 31:20:@11.6]
  assign _GEN_1026 = 9'h1 == _T_538 ? _T_22_1 : _T_22_0; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1027 = 9'h2 == _T_538 ? _T_22_2 : _GEN_1026; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1028 = 9'h3 == _T_538 ? _T_22_3 : _GEN_1027; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1029 = 9'h4 == _T_538 ? _T_22_4 : _GEN_1028; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1030 = 9'h5 == _T_538 ? _T_22_5 : _GEN_1029; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1031 = 9'h6 == _T_538 ? _T_22_6 : _GEN_1030; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1032 = 9'h7 == _T_538 ? _T_22_7 : _GEN_1031; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1033 = 9'h8 == _T_538 ? _T_22_8 : _GEN_1032; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1034 = 9'h9 == _T_538 ? _T_22_9 : _GEN_1033; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1035 = 9'ha == _T_538 ? _T_22_10 : _GEN_1034; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1036 = 9'hb == _T_538 ? _T_22_11 : _GEN_1035; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1037 = 9'hc == _T_538 ? _T_22_12 : _GEN_1036; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1038 = 9'hd == _T_538 ? _T_22_13 : _GEN_1037; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1039 = 9'he == _T_538 ? _T_22_14 : _GEN_1038; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1040 = 9'hf == _T_538 ? _T_22_15 : _GEN_1039; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1041 = 9'h10 == _T_538 ? _T_22_16 : _GEN_1040; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1042 = 9'h11 == _T_538 ? _T_22_17 : _GEN_1041; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1043 = 9'h12 == _T_538 ? _T_22_18 : _GEN_1042; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1044 = 9'h13 == _T_538 ? _T_22_19 : _GEN_1043; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1045 = 9'h14 == _T_538 ? _T_22_20 : _GEN_1044; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1046 = 9'h15 == _T_538 ? _T_22_21 : _GEN_1045; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1047 = 9'h16 == _T_538 ? _T_22_22 : _GEN_1046; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1048 = 9'h17 == _T_538 ? _T_22_23 : _GEN_1047; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1049 = 9'h18 == _T_538 ? _T_22_24 : _GEN_1048; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1050 = 9'h19 == _T_538 ? _T_22_25 : _GEN_1049; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1051 = 9'h1a == _T_538 ? _T_22_26 : _GEN_1050; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1052 = 9'h1b == _T_538 ? _T_22_27 : _GEN_1051; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1053 = 9'h1c == _T_538 ? _T_22_28 : _GEN_1052; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1054 = 9'h1d == _T_538 ? _T_22_29 : _GEN_1053; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1055 = 9'h1e == _T_538 ? _T_22_30 : _GEN_1054; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1056 = 9'h1f == _T_538 ? _T_22_31 : _GEN_1055; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1057 = 9'h20 == _T_538 ? _T_22_32 : _GEN_1056; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1058 = 9'h21 == _T_538 ? _T_22_33 : _GEN_1057; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1059 = 9'h22 == _T_538 ? _T_22_34 : _GEN_1058; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1060 = 9'h23 == _T_538 ? _T_22_35 : _GEN_1059; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1061 = 9'h24 == _T_538 ? _T_22_36 : _GEN_1060; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1062 = 9'h25 == _T_538 ? _T_22_37 : _GEN_1061; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1063 = 9'h26 == _T_538 ? _T_22_38 : _GEN_1062; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1064 = 9'h27 == _T_538 ? _T_22_39 : _GEN_1063; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1065 = 9'h28 == _T_538 ? _T_22_40 : _GEN_1064; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1066 = 9'h29 == _T_538 ? _T_22_41 : _GEN_1065; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1067 = 9'h2a == _T_538 ? _T_22_42 : _GEN_1066; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1068 = 9'h2b == _T_538 ? _T_22_43 : _GEN_1067; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1069 = 9'h2c == _T_538 ? _T_22_44 : _GEN_1068; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1070 = 9'h2d == _T_538 ? _T_22_45 : _GEN_1069; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1071 = 9'h2e == _T_538 ? _T_22_46 : _GEN_1070; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1072 = 9'h2f == _T_538 ? _T_22_47 : _GEN_1071; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1073 = 9'h30 == _T_538 ? _T_22_48 : _GEN_1072; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1074 = 9'h31 == _T_538 ? _T_22_49 : _GEN_1073; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1075 = 9'h32 == _T_538 ? _T_22_50 : _GEN_1074; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1076 = 9'h33 == _T_538 ? _T_22_51 : _GEN_1075; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1077 = 9'h34 == _T_538 ? _T_22_52 : _GEN_1076; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1078 = 9'h35 == _T_538 ? _T_22_53 : _GEN_1077; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1079 = 9'h36 == _T_538 ? _T_22_54 : _GEN_1078; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1080 = 9'h37 == _T_538 ? _T_22_55 : _GEN_1079; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1081 = 9'h38 == _T_538 ? _T_22_56 : _GEN_1080; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1082 = 9'h39 == _T_538 ? _T_22_57 : _GEN_1081; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1083 = 9'h3a == _T_538 ? _T_22_58 : _GEN_1082; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1084 = 9'h3b == _T_538 ? _T_22_59 : _GEN_1083; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1085 = 9'h3c == _T_538 ? _T_22_60 : _GEN_1084; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1086 = 9'h3d == _T_538 ? _T_22_61 : _GEN_1085; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1087 = 9'h3e == _T_538 ? _T_22_62 : _GEN_1086; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1088 = 9'h3f == _T_538 ? _T_22_63 : _GEN_1087; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1089 = 9'h40 == _T_538 ? _T_22_64 : _GEN_1088; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1090 = 9'h41 == _T_538 ? _T_22_65 : _GEN_1089; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1091 = 9'h42 == _T_538 ? _T_22_66 : _GEN_1090; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1092 = 9'h43 == _T_538 ? _T_22_67 : _GEN_1091; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1093 = 9'h44 == _T_538 ? _T_22_68 : _GEN_1092; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1094 = 9'h45 == _T_538 ? _T_22_69 : _GEN_1093; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1095 = 9'h46 == _T_538 ? _T_22_70 : _GEN_1094; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1096 = 9'h47 == _T_538 ? _T_22_71 : _GEN_1095; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1097 = 9'h48 == _T_538 ? _T_22_72 : _GEN_1096; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1098 = 9'h49 == _T_538 ? _T_22_73 : _GEN_1097; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1099 = 9'h4a == _T_538 ? _T_22_74 : _GEN_1098; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1100 = 9'h4b == _T_538 ? _T_22_75 : _GEN_1099; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1101 = 9'h4c == _T_538 ? _T_22_76 : _GEN_1100; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1102 = 9'h4d == _T_538 ? _T_22_77 : _GEN_1101; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1103 = 9'h4e == _T_538 ? _T_22_78 : _GEN_1102; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1104 = 9'h4f == _T_538 ? _T_22_79 : _GEN_1103; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1105 = 9'h50 == _T_538 ? _T_22_80 : _GEN_1104; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1106 = 9'h51 == _T_538 ? _T_22_81 : _GEN_1105; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1107 = 9'h52 == _T_538 ? _T_22_82 : _GEN_1106; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1108 = 9'h53 == _T_538 ? _T_22_83 : _GEN_1107; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1109 = 9'h54 == _T_538 ? _T_22_84 : _GEN_1108; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1110 = 9'h55 == _T_538 ? _T_22_85 : _GEN_1109; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1111 = 9'h56 == _T_538 ? _T_22_86 : _GEN_1110; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1112 = 9'h57 == _T_538 ? _T_22_87 : _GEN_1111; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1113 = 9'h58 == _T_538 ? _T_22_88 : _GEN_1112; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1114 = 9'h59 == _T_538 ? _T_22_89 : _GEN_1113; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1115 = 9'h5a == _T_538 ? _T_22_90 : _GEN_1114; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1116 = 9'h5b == _T_538 ? _T_22_91 : _GEN_1115; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1117 = 9'h5c == _T_538 ? _T_22_92 : _GEN_1116; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1118 = 9'h5d == _T_538 ? _T_22_93 : _GEN_1117; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1119 = 9'h5e == _T_538 ? _T_22_94 : _GEN_1118; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1120 = 9'h5f == _T_538 ? _T_22_95 : _GEN_1119; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1121 = 9'h60 == _T_538 ? _T_22_96 : _GEN_1120; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1122 = 9'h61 == _T_538 ? _T_22_97 : _GEN_1121; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1123 = 9'h62 == _T_538 ? _T_22_98 : _GEN_1122; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1124 = 9'h63 == _T_538 ? _T_22_99 : _GEN_1123; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1125 = 9'h64 == _T_538 ? _T_22_100 : _GEN_1124; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1126 = 9'h65 == _T_538 ? _T_22_101 : _GEN_1125; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1127 = 9'h66 == _T_538 ? _T_22_102 : _GEN_1126; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1128 = 9'h67 == _T_538 ? _T_22_103 : _GEN_1127; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1129 = 9'h68 == _T_538 ? _T_22_104 : _GEN_1128; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1130 = 9'h69 == _T_538 ? _T_22_105 : _GEN_1129; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1131 = 9'h6a == _T_538 ? _T_22_106 : _GEN_1130; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1132 = 9'h6b == _T_538 ? _T_22_107 : _GEN_1131; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1133 = 9'h6c == _T_538 ? _T_22_108 : _GEN_1132; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1134 = 9'h6d == _T_538 ? _T_22_109 : _GEN_1133; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1135 = 9'h6e == _T_538 ? _T_22_110 : _GEN_1134; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1136 = 9'h6f == _T_538 ? _T_22_111 : _GEN_1135; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1137 = 9'h70 == _T_538 ? _T_22_112 : _GEN_1136; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1138 = 9'h71 == _T_538 ? _T_22_113 : _GEN_1137; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1139 = 9'h72 == _T_538 ? _T_22_114 : _GEN_1138; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1140 = 9'h73 == _T_538 ? _T_22_115 : _GEN_1139; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1141 = 9'h74 == _T_538 ? _T_22_116 : _GEN_1140; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1142 = 9'h75 == _T_538 ? _T_22_117 : _GEN_1141; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1143 = 9'h76 == _T_538 ? _T_22_118 : _GEN_1142; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1144 = 9'h77 == _T_538 ? _T_22_119 : _GEN_1143; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1145 = 9'h78 == _T_538 ? _T_22_120 : _GEN_1144; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1146 = 9'h79 == _T_538 ? _T_22_121 : _GEN_1145; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1147 = 9'h7a == _T_538 ? _T_22_122 : _GEN_1146; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1148 = 9'h7b == _T_538 ? _T_22_123 : _GEN_1147; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1149 = 9'h7c == _T_538 ? _T_22_124 : _GEN_1148; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1150 = 9'h7d == _T_538 ? _T_22_125 : _GEN_1149; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1151 = 9'h7e == _T_538 ? _T_22_126 : _GEN_1150; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1152 = 9'h7f == _T_538 ? _T_22_127 : _GEN_1151; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1153 = 9'h80 == _T_538 ? _T_22_128 : _GEN_1152; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1154 = 9'h81 == _T_538 ? _T_22_129 : _GEN_1153; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1155 = 9'h82 == _T_538 ? _T_22_130 : _GEN_1154; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1156 = 9'h83 == _T_538 ? _T_22_131 : _GEN_1155; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1157 = 9'h84 == _T_538 ? _T_22_132 : _GEN_1156; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1158 = 9'h85 == _T_538 ? _T_22_133 : _GEN_1157; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1159 = 9'h86 == _T_538 ? _T_22_134 : _GEN_1158; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1160 = 9'h87 == _T_538 ? _T_22_135 : _GEN_1159; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1161 = 9'h88 == _T_538 ? _T_22_136 : _GEN_1160; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1162 = 9'h89 == _T_538 ? _T_22_137 : _GEN_1161; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1163 = 9'h8a == _T_538 ? _T_22_138 : _GEN_1162; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1164 = 9'h8b == _T_538 ? _T_22_139 : _GEN_1163; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1165 = 9'h8c == _T_538 ? _T_22_140 : _GEN_1164; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1166 = 9'h8d == _T_538 ? _T_22_141 : _GEN_1165; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1167 = 9'h8e == _T_538 ? _T_22_142 : _GEN_1166; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1168 = 9'h8f == _T_538 ? _T_22_143 : _GEN_1167; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1169 = 9'h90 == _T_538 ? _T_22_144 : _GEN_1168; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1170 = 9'h91 == _T_538 ? _T_22_145 : _GEN_1169; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1171 = 9'h92 == _T_538 ? _T_22_146 : _GEN_1170; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1172 = 9'h93 == _T_538 ? _T_22_147 : _GEN_1171; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1173 = 9'h94 == _T_538 ? _T_22_148 : _GEN_1172; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1174 = 9'h95 == _T_538 ? _T_22_149 : _GEN_1173; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1175 = 9'h96 == _T_538 ? _T_22_150 : _GEN_1174; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1176 = 9'h97 == _T_538 ? _T_22_151 : _GEN_1175; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1177 = 9'h98 == _T_538 ? _T_22_152 : _GEN_1176; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1178 = 9'h99 == _T_538 ? _T_22_153 : _GEN_1177; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1179 = 9'h9a == _T_538 ? _T_22_154 : _GEN_1178; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1180 = 9'h9b == _T_538 ? _T_22_155 : _GEN_1179; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1181 = 9'h9c == _T_538 ? _T_22_156 : _GEN_1180; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1182 = 9'h9d == _T_538 ? _T_22_157 : _GEN_1181; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1183 = 9'h9e == _T_538 ? _T_22_158 : _GEN_1182; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1184 = 9'h9f == _T_538 ? _T_22_159 : _GEN_1183; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1185 = 9'ha0 == _T_538 ? _T_22_160 : _GEN_1184; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1186 = 9'ha1 == _T_538 ? _T_22_161 : _GEN_1185; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1187 = 9'ha2 == _T_538 ? _T_22_162 : _GEN_1186; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1188 = 9'ha3 == _T_538 ? _T_22_163 : _GEN_1187; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1189 = 9'ha4 == _T_538 ? _T_22_164 : _GEN_1188; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1190 = 9'ha5 == _T_538 ? _T_22_165 : _GEN_1189; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1191 = 9'ha6 == _T_538 ? _T_22_166 : _GEN_1190; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1192 = 9'ha7 == _T_538 ? _T_22_167 : _GEN_1191; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1193 = 9'ha8 == _T_538 ? _T_22_168 : _GEN_1192; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1194 = 9'ha9 == _T_538 ? _T_22_169 : _GEN_1193; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1195 = 9'haa == _T_538 ? _T_22_170 : _GEN_1194; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1196 = 9'hab == _T_538 ? _T_22_171 : _GEN_1195; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1197 = 9'hac == _T_538 ? _T_22_172 : _GEN_1196; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1198 = 9'had == _T_538 ? _T_22_173 : _GEN_1197; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1199 = 9'hae == _T_538 ? _T_22_174 : _GEN_1198; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1200 = 9'haf == _T_538 ? _T_22_175 : _GEN_1199; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1201 = 9'hb0 == _T_538 ? _T_22_176 : _GEN_1200; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1202 = 9'hb1 == _T_538 ? _T_22_177 : _GEN_1201; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1203 = 9'hb2 == _T_538 ? _T_22_178 : _GEN_1202; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1204 = 9'hb3 == _T_538 ? _T_22_179 : _GEN_1203; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1205 = 9'hb4 == _T_538 ? _T_22_180 : _GEN_1204; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1206 = 9'hb5 == _T_538 ? _T_22_181 : _GEN_1205; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1207 = 9'hb6 == _T_538 ? _T_22_182 : _GEN_1206; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1208 = 9'hb7 == _T_538 ? _T_22_183 : _GEN_1207; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1209 = 9'hb8 == _T_538 ? _T_22_184 : _GEN_1208; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1210 = 9'hb9 == _T_538 ? _T_22_185 : _GEN_1209; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1211 = 9'hba == _T_538 ? _T_22_186 : _GEN_1210; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1212 = 9'hbb == _T_538 ? _T_22_187 : _GEN_1211; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1213 = 9'hbc == _T_538 ? _T_22_188 : _GEN_1212; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1214 = 9'hbd == _T_538 ? _T_22_189 : _GEN_1213; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1215 = 9'hbe == _T_538 ? _T_22_190 : _GEN_1214; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1216 = 9'hbf == _T_538 ? _T_22_191 : _GEN_1215; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1217 = 9'hc0 == _T_538 ? _T_22_192 : _GEN_1216; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1218 = 9'hc1 == _T_538 ? _T_22_193 : _GEN_1217; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1219 = 9'hc2 == _T_538 ? _T_22_194 : _GEN_1218; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1220 = 9'hc3 == _T_538 ? _T_22_195 : _GEN_1219; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1221 = 9'hc4 == _T_538 ? _T_22_196 : _GEN_1220; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1222 = 9'hc5 == _T_538 ? _T_22_197 : _GEN_1221; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1223 = 9'hc6 == _T_538 ? _T_22_198 : _GEN_1222; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1224 = 9'hc7 == _T_538 ? _T_22_199 : _GEN_1223; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1225 = 9'hc8 == _T_538 ? _T_22_200 : _GEN_1224; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1226 = 9'hc9 == _T_538 ? _T_22_201 : _GEN_1225; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1227 = 9'hca == _T_538 ? _T_22_202 : _GEN_1226; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1228 = 9'hcb == _T_538 ? _T_22_203 : _GEN_1227; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1229 = 9'hcc == _T_538 ? _T_22_204 : _GEN_1228; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1230 = 9'hcd == _T_538 ? _T_22_205 : _GEN_1229; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1231 = 9'hce == _T_538 ? _T_22_206 : _GEN_1230; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1232 = 9'hcf == _T_538 ? _T_22_207 : _GEN_1231; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1233 = 9'hd0 == _T_538 ? _T_22_208 : _GEN_1232; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1234 = 9'hd1 == _T_538 ? _T_22_209 : _GEN_1233; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1235 = 9'hd2 == _T_538 ? _T_22_210 : _GEN_1234; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1236 = 9'hd3 == _T_538 ? _T_22_211 : _GEN_1235; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1237 = 9'hd4 == _T_538 ? _T_22_212 : _GEN_1236; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1238 = 9'hd5 == _T_538 ? _T_22_213 : _GEN_1237; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1239 = 9'hd6 == _T_538 ? _T_22_214 : _GEN_1238; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1240 = 9'hd7 == _T_538 ? _T_22_215 : _GEN_1239; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1241 = 9'hd8 == _T_538 ? _T_22_216 : _GEN_1240; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1242 = 9'hd9 == _T_538 ? _T_22_217 : _GEN_1241; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1243 = 9'hda == _T_538 ? _T_22_218 : _GEN_1242; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1244 = 9'hdb == _T_538 ? _T_22_219 : _GEN_1243; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1245 = 9'hdc == _T_538 ? _T_22_220 : _GEN_1244; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1246 = 9'hdd == _T_538 ? _T_22_221 : _GEN_1245; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1247 = 9'hde == _T_538 ? _T_22_222 : _GEN_1246; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1248 = 9'hdf == _T_538 ? _T_22_223 : _GEN_1247; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1249 = 9'he0 == _T_538 ? _T_22_224 : _GEN_1248; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1250 = 9'he1 == _T_538 ? _T_22_225 : _GEN_1249; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1251 = 9'he2 == _T_538 ? _T_22_226 : _GEN_1250; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1252 = 9'he3 == _T_538 ? _T_22_227 : _GEN_1251; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1253 = 9'he4 == _T_538 ? _T_22_228 : _GEN_1252; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1254 = 9'he5 == _T_538 ? _T_22_229 : _GEN_1253; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1255 = 9'he6 == _T_538 ? _T_22_230 : _GEN_1254; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1256 = 9'he7 == _T_538 ? _T_22_231 : _GEN_1255; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1257 = 9'he8 == _T_538 ? _T_22_232 : _GEN_1256; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1258 = 9'he9 == _T_538 ? _T_22_233 : _GEN_1257; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1259 = 9'hea == _T_538 ? _T_22_234 : _GEN_1258; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1260 = 9'heb == _T_538 ? _T_22_235 : _GEN_1259; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1261 = 9'hec == _T_538 ? _T_22_236 : _GEN_1260; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1262 = 9'hed == _T_538 ? _T_22_237 : _GEN_1261; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1263 = 9'hee == _T_538 ? _T_22_238 : _GEN_1262; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1264 = 9'hef == _T_538 ? _T_22_239 : _GEN_1263; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1265 = 9'hf0 == _T_538 ? _T_22_240 : _GEN_1264; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1266 = 9'hf1 == _T_538 ? _T_22_241 : _GEN_1265; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1267 = 9'hf2 == _T_538 ? _T_22_242 : _GEN_1266; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1268 = 9'hf3 == _T_538 ? _T_22_243 : _GEN_1267; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1269 = 9'hf4 == _T_538 ? _T_22_244 : _GEN_1268; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1270 = 9'hf5 == _T_538 ? _T_22_245 : _GEN_1269; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1271 = 9'hf6 == _T_538 ? _T_22_246 : _GEN_1270; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1272 = 9'hf7 == _T_538 ? _T_22_247 : _GEN_1271; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1273 = 9'hf8 == _T_538 ? _T_22_248 : _GEN_1272; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1274 = 9'hf9 == _T_538 ? _T_22_249 : _GEN_1273; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1275 = 9'hfa == _T_538 ? _T_22_250 : _GEN_1274; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1276 = 9'hfb == _T_538 ? _T_22_251 : _GEN_1275; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1277 = 9'hfc == _T_538 ? _T_22_252 : _GEN_1276; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1278 = 9'hfd == _T_538 ? _T_22_253 : _GEN_1277; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1279 = 9'hfe == _T_538 ? _T_22_254 : _GEN_1278; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1280 = 9'hff == _T_538 ? _T_22_255 : _GEN_1279; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1281 = 9'h100 == _T_538 ? _T_22_256 : _GEN_1280; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1282 = 9'h101 == _T_538 ? _T_22_257 : _GEN_1281; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1283 = 9'h102 == _T_538 ? _T_22_258 : _GEN_1282; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1284 = 9'h103 == _T_538 ? _T_22_259 : _GEN_1283; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1285 = 9'h104 == _T_538 ? _T_22_260 : _GEN_1284; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1286 = 9'h105 == _T_538 ? _T_22_261 : _GEN_1285; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1287 = 9'h106 == _T_538 ? _T_22_262 : _GEN_1286; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1288 = 9'h107 == _T_538 ? _T_22_263 : _GEN_1287; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1289 = 9'h108 == _T_538 ? _T_22_264 : _GEN_1288; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1290 = 9'h109 == _T_538 ? _T_22_265 : _GEN_1289; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1291 = 9'h10a == _T_538 ? _T_22_266 : _GEN_1290; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1292 = 9'h10b == _T_538 ? _T_22_267 : _GEN_1291; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1293 = 9'h10c == _T_538 ? _T_22_268 : _GEN_1292; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1294 = 9'h10d == _T_538 ? _T_22_269 : _GEN_1293; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1295 = 9'h10e == _T_538 ? _T_22_270 : _GEN_1294; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1296 = 9'h10f == _T_538 ? _T_22_271 : _GEN_1295; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1297 = 9'h110 == _T_538 ? _T_22_272 : _GEN_1296; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1298 = 9'h111 == _T_538 ? _T_22_273 : _GEN_1297; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1299 = 9'h112 == _T_538 ? _T_22_274 : _GEN_1298; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1300 = 9'h113 == _T_538 ? _T_22_275 : _GEN_1299; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1301 = 9'h114 == _T_538 ? _T_22_276 : _GEN_1300; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1302 = 9'h115 == _T_538 ? _T_22_277 : _GEN_1301; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1303 = 9'h116 == _T_538 ? _T_22_278 : _GEN_1302; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1304 = 9'h117 == _T_538 ? _T_22_279 : _GEN_1303; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1305 = 9'h118 == _T_538 ? _T_22_280 : _GEN_1304; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1306 = 9'h119 == _T_538 ? _T_22_281 : _GEN_1305; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1307 = 9'h11a == _T_538 ? _T_22_282 : _GEN_1306; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1308 = 9'h11b == _T_538 ? _T_22_283 : _GEN_1307; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1309 = 9'h11c == _T_538 ? _T_22_284 : _GEN_1308; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1310 = 9'h11d == _T_538 ? _T_22_285 : _GEN_1309; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1311 = 9'h11e == _T_538 ? _T_22_286 : _GEN_1310; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1312 = 9'h11f == _T_538 ? _T_22_287 : _GEN_1311; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1313 = 9'h120 == _T_538 ? _T_22_288 : _GEN_1312; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1314 = 9'h121 == _T_538 ? _T_22_289 : _GEN_1313; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1315 = 9'h122 == _T_538 ? _T_22_290 : _GEN_1314; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1316 = 9'h123 == _T_538 ? _T_22_291 : _GEN_1315; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1317 = 9'h124 == _T_538 ? _T_22_292 : _GEN_1316; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1318 = 9'h125 == _T_538 ? _T_22_293 : _GEN_1317; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1319 = 9'h126 == _T_538 ? _T_22_294 : _GEN_1318; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1320 = 9'h127 == _T_538 ? _T_22_295 : _GEN_1319; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1321 = 9'h128 == _T_538 ? _T_22_296 : _GEN_1320; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1322 = 9'h129 == _T_538 ? _T_22_297 : _GEN_1321; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1323 = 9'h12a == _T_538 ? _T_22_298 : _GEN_1322; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1324 = 9'h12b == _T_538 ? _T_22_299 : _GEN_1323; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1325 = 9'h12c == _T_538 ? _T_22_300 : _GEN_1324; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1326 = 9'h12d == _T_538 ? _T_22_301 : _GEN_1325; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1327 = 9'h12e == _T_538 ? _T_22_302 : _GEN_1326; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1328 = 9'h12f == _T_538 ? _T_22_303 : _GEN_1327; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1329 = 9'h130 == _T_538 ? _T_22_304 : _GEN_1328; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1330 = 9'h131 == _T_538 ? _T_22_305 : _GEN_1329; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1331 = 9'h132 == _T_538 ? _T_22_306 : _GEN_1330; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1332 = 9'h133 == _T_538 ? _T_22_307 : _GEN_1331; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1333 = 9'h134 == _T_538 ? _T_22_308 : _GEN_1332; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1334 = 9'h135 == _T_538 ? _T_22_309 : _GEN_1333; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1335 = 9'h136 == _T_538 ? _T_22_310 : _GEN_1334; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1336 = 9'h137 == _T_538 ? _T_22_311 : _GEN_1335; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1337 = 9'h138 == _T_538 ? _T_22_312 : _GEN_1336; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1338 = 9'h139 == _T_538 ? _T_22_313 : _GEN_1337; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1339 = 9'h13a == _T_538 ? _T_22_314 : _GEN_1338; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1340 = 9'h13b == _T_538 ? _T_22_315 : _GEN_1339; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1341 = 9'h13c == _T_538 ? _T_22_316 : _GEN_1340; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1342 = 9'h13d == _T_538 ? _T_22_317 : _GEN_1341; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1343 = 9'h13e == _T_538 ? _T_22_318 : _GEN_1342; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1344 = 9'h13f == _T_538 ? _T_22_319 : _GEN_1343; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1345 = 9'h140 == _T_538 ? _T_22_320 : _GEN_1344; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1346 = 9'h141 == _T_538 ? _T_22_321 : _GEN_1345; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1347 = 9'h142 == _T_538 ? _T_22_322 : _GEN_1346; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1348 = 9'h143 == _T_538 ? _T_22_323 : _GEN_1347; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1349 = 9'h144 == _T_538 ? _T_22_324 : _GEN_1348; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1350 = 9'h145 == _T_538 ? _T_22_325 : _GEN_1349; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1351 = 9'h146 == _T_538 ? _T_22_326 : _GEN_1350; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1352 = 9'h147 == _T_538 ? _T_22_327 : _GEN_1351; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1353 = 9'h148 == _T_538 ? _T_22_328 : _GEN_1352; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1354 = 9'h149 == _T_538 ? _T_22_329 : _GEN_1353; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1355 = 9'h14a == _T_538 ? _T_22_330 : _GEN_1354; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1356 = 9'h14b == _T_538 ? _T_22_331 : _GEN_1355; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1357 = 9'h14c == _T_538 ? _T_22_332 : _GEN_1356; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1358 = 9'h14d == _T_538 ? _T_22_333 : _GEN_1357; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1359 = 9'h14e == _T_538 ? _T_22_334 : _GEN_1358; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1360 = 9'h14f == _T_538 ? _T_22_335 : _GEN_1359; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1361 = 9'h150 == _T_538 ? _T_22_336 : _GEN_1360; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1362 = 9'h151 == _T_538 ? _T_22_337 : _GEN_1361; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1363 = 9'h152 == _T_538 ? _T_22_338 : _GEN_1362; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1364 = 9'h153 == _T_538 ? _T_22_339 : _GEN_1363; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1365 = 9'h154 == _T_538 ? _T_22_340 : _GEN_1364; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1366 = 9'h155 == _T_538 ? _T_22_341 : _GEN_1365; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1367 = 9'h156 == _T_538 ? _T_22_342 : _GEN_1366; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1368 = 9'h157 == _T_538 ? _T_22_343 : _GEN_1367; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1369 = 9'h158 == _T_538 ? _T_22_344 : _GEN_1368; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1370 = 9'h159 == _T_538 ? _T_22_345 : _GEN_1369; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1371 = 9'h15a == _T_538 ? _T_22_346 : _GEN_1370; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1372 = 9'h15b == _T_538 ? _T_22_347 : _GEN_1371; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1373 = 9'h15c == _T_538 ? _T_22_348 : _GEN_1372; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1374 = 9'h15d == _T_538 ? _T_22_349 : _GEN_1373; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1375 = 9'h15e == _T_538 ? _T_22_350 : _GEN_1374; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1376 = 9'h15f == _T_538 ? _T_22_351 : _GEN_1375; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1377 = 9'h160 == _T_538 ? _T_22_352 : _GEN_1376; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1378 = 9'h161 == _T_538 ? _T_22_353 : _GEN_1377; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1379 = 9'h162 == _T_538 ? _T_22_354 : _GEN_1378; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1380 = 9'h163 == _T_538 ? _T_22_355 : _GEN_1379; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1381 = 9'h164 == _T_538 ? _T_22_356 : _GEN_1380; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1382 = 9'h165 == _T_538 ? _T_22_357 : _GEN_1381; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1383 = 9'h166 == _T_538 ? _T_22_358 : _GEN_1382; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1384 = 9'h167 == _T_538 ? _T_22_359 : _GEN_1383; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1385 = 9'h168 == _T_538 ? _T_22_360 : _GEN_1384; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1386 = 9'h169 == _T_538 ? _T_22_361 : _GEN_1385; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1387 = 9'h16a == _T_538 ? _T_22_362 : _GEN_1386; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1388 = 9'h16b == _T_538 ? _T_22_363 : _GEN_1387; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1389 = 9'h16c == _T_538 ? _T_22_364 : _GEN_1388; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1390 = 9'h16d == _T_538 ? _T_22_365 : _GEN_1389; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1391 = 9'h16e == _T_538 ? _T_22_366 : _GEN_1390; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1392 = 9'h16f == _T_538 ? _T_22_367 : _GEN_1391; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1393 = 9'h170 == _T_538 ? _T_22_368 : _GEN_1392; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1394 = 9'h171 == _T_538 ? _T_22_369 : _GEN_1393; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1395 = 9'h172 == _T_538 ? _T_22_370 : _GEN_1394; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1396 = 9'h173 == _T_538 ? _T_22_371 : _GEN_1395; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1397 = 9'h174 == _T_538 ? _T_22_372 : _GEN_1396; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1398 = 9'h175 == _T_538 ? _T_22_373 : _GEN_1397; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1399 = 9'h176 == _T_538 ? _T_22_374 : _GEN_1398; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1400 = 9'h177 == _T_538 ? _T_22_375 : _GEN_1399; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1401 = 9'h178 == _T_538 ? _T_22_376 : _GEN_1400; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1402 = 9'h179 == _T_538 ? _T_22_377 : _GEN_1401; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1403 = 9'h17a == _T_538 ? _T_22_378 : _GEN_1402; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1404 = 9'h17b == _T_538 ? _T_22_379 : _GEN_1403; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1405 = 9'h17c == _T_538 ? _T_22_380 : _GEN_1404; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1406 = 9'h17d == _T_538 ? _T_22_381 : _GEN_1405; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1407 = 9'h17e == _T_538 ? _T_22_382 : _GEN_1406; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1408 = 9'h17f == _T_538 ? _T_22_383 : _GEN_1407; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1409 = 9'h180 == _T_538 ? _T_22_384 : _GEN_1408; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1410 = 9'h181 == _T_538 ? _T_22_385 : _GEN_1409; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1411 = 9'h182 == _T_538 ? _T_22_386 : _GEN_1410; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1412 = 9'h183 == _T_538 ? _T_22_387 : _GEN_1411; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1413 = 9'h184 == _T_538 ? _T_22_388 : _GEN_1412; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1414 = 9'h185 == _T_538 ? _T_22_389 : _GEN_1413; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1415 = 9'h186 == _T_538 ? _T_22_390 : _GEN_1414; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1416 = 9'h187 == _T_538 ? _T_22_391 : _GEN_1415; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1417 = 9'h188 == _T_538 ? _T_22_392 : _GEN_1416; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1418 = 9'h189 == _T_538 ? _T_22_393 : _GEN_1417; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1419 = 9'h18a == _T_538 ? _T_22_394 : _GEN_1418; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1420 = 9'h18b == _T_538 ? _T_22_395 : _GEN_1419; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1421 = 9'h18c == _T_538 ? _T_22_396 : _GEN_1420; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1422 = 9'h18d == _T_538 ? _T_22_397 : _GEN_1421; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1423 = 9'h18e == _T_538 ? _T_22_398 : _GEN_1422; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1424 = 9'h18f == _T_538 ? _T_22_399 : _GEN_1423; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1425 = 9'h190 == _T_538 ? _T_22_400 : _GEN_1424; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1426 = 9'h191 == _T_538 ? _T_22_401 : _GEN_1425; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1427 = 9'h192 == _T_538 ? _T_22_402 : _GEN_1426; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1428 = 9'h193 == _T_538 ? _T_22_403 : _GEN_1427; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1429 = 9'h194 == _T_538 ? _T_22_404 : _GEN_1428; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1430 = 9'h195 == _T_538 ? _T_22_405 : _GEN_1429; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1431 = 9'h196 == _T_538 ? _T_22_406 : _GEN_1430; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1432 = 9'h197 == _T_538 ? _T_22_407 : _GEN_1431; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1433 = 9'h198 == _T_538 ? _T_22_408 : _GEN_1432; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1434 = 9'h199 == _T_538 ? _T_22_409 : _GEN_1433; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1435 = 9'h19a == _T_538 ? _T_22_410 : _GEN_1434; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1436 = 9'h19b == _T_538 ? _T_22_411 : _GEN_1435; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1437 = 9'h19c == _T_538 ? _T_22_412 : _GEN_1436; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1438 = 9'h19d == _T_538 ? _T_22_413 : _GEN_1437; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1439 = 9'h19e == _T_538 ? _T_22_414 : _GEN_1438; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1440 = 9'h19f == _T_538 ? _T_22_415 : _GEN_1439; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1441 = 9'h1a0 == _T_538 ? _T_22_416 : _GEN_1440; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1442 = 9'h1a1 == _T_538 ? _T_22_417 : _GEN_1441; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1443 = 9'h1a2 == _T_538 ? _T_22_418 : _GEN_1442; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1444 = 9'h1a3 == _T_538 ? _T_22_419 : _GEN_1443; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1445 = 9'h1a4 == _T_538 ? _T_22_420 : _GEN_1444; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1446 = 9'h1a5 == _T_538 ? _T_22_421 : _GEN_1445; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1447 = 9'h1a6 == _T_538 ? _T_22_422 : _GEN_1446; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1448 = 9'h1a7 == _T_538 ? _T_22_423 : _GEN_1447; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1449 = 9'h1a8 == _T_538 ? _T_22_424 : _GEN_1448; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1450 = 9'h1a9 == _T_538 ? _T_22_425 : _GEN_1449; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1451 = 9'h1aa == _T_538 ? _T_22_426 : _GEN_1450; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1452 = 9'h1ab == _T_538 ? _T_22_427 : _GEN_1451; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1453 = 9'h1ac == _T_538 ? _T_22_428 : _GEN_1452; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1454 = 9'h1ad == _T_538 ? _T_22_429 : _GEN_1453; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1455 = 9'h1ae == _T_538 ? _T_22_430 : _GEN_1454; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1456 = 9'h1af == _T_538 ? _T_22_431 : _GEN_1455; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1457 = 9'h1b0 == _T_538 ? _T_22_432 : _GEN_1456; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1458 = 9'h1b1 == _T_538 ? _T_22_433 : _GEN_1457; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1459 = 9'h1b2 == _T_538 ? _T_22_434 : _GEN_1458; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1460 = 9'h1b3 == _T_538 ? _T_22_435 : _GEN_1459; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1461 = 9'h1b4 == _T_538 ? _T_22_436 : _GEN_1460; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1462 = 9'h1b5 == _T_538 ? _T_22_437 : _GEN_1461; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1463 = 9'h1b6 == _T_538 ? _T_22_438 : _GEN_1462; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1464 = 9'h1b7 == _T_538 ? _T_22_439 : _GEN_1463; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1465 = 9'h1b8 == _T_538 ? _T_22_440 : _GEN_1464; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1466 = 9'h1b9 == _T_538 ? _T_22_441 : _GEN_1465; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1467 = 9'h1ba == _T_538 ? _T_22_442 : _GEN_1466; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1468 = 9'h1bb == _T_538 ? _T_22_443 : _GEN_1467; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1469 = 9'h1bc == _T_538 ? _T_22_444 : _GEN_1468; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1470 = 9'h1bd == _T_538 ? _T_22_445 : _GEN_1469; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1471 = 9'h1be == _T_538 ? _T_22_446 : _GEN_1470; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1472 = 9'h1bf == _T_538 ? _T_22_447 : _GEN_1471; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1473 = 9'h1c0 == _T_538 ? _T_22_448 : _GEN_1472; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1474 = 9'h1c1 == _T_538 ? _T_22_449 : _GEN_1473; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1475 = 9'h1c2 == _T_538 ? _T_22_450 : _GEN_1474; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1476 = 9'h1c3 == _T_538 ? _T_22_451 : _GEN_1475; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1477 = 9'h1c4 == _T_538 ? _T_22_452 : _GEN_1476; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1478 = 9'h1c5 == _T_538 ? _T_22_453 : _GEN_1477; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1479 = 9'h1c6 == _T_538 ? _T_22_454 : _GEN_1478; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1480 = 9'h1c7 == _T_538 ? _T_22_455 : _GEN_1479; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1481 = 9'h1c8 == _T_538 ? _T_22_456 : _GEN_1480; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1482 = 9'h1c9 == _T_538 ? _T_22_457 : _GEN_1481; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1483 = 9'h1ca == _T_538 ? _T_22_458 : _GEN_1482; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1484 = 9'h1cb == _T_538 ? _T_22_459 : _GEN_1483; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1485 = 9'h1cc == _T_538 ? _T_22_460 : _GEN_1484; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1486 = 9'h1cd == _T_538 ? _T_22_461 : _GEN_1485; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1487 = 9'h1ce == _T_538 ? _T_22_462 : _GEN_1486; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1488 = 9'h1cf == _T_538 ? _T_22_463 : _GEN_1487; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1489 = 9'h1d0 == _T_538 ? _T_22_464 : _GEN_1488; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1490 = 9'h1d1 == _T_538 ? _T_22_465 : _GEN_1489; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1491 = 9'h1d2 == _T_538 ? _T_22_466 : _GEN_1490; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1492 = 9'h1d3 == _T_538 ? _T_22_467 : _GEN_1491; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1493 = 9'h1d4 == _T_538 ? _T_22_468 : _GEN_1492; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1494 = 9'h1d5 == _T_538 ? _T_22_469 : _GEN_1493; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1495 = 9'h1d6 == _T_538 ? _T_22_470 : _GEN_1494; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1496 = 9'h1d7 == _T_538 ? _T_22_471 : _GEN_1495; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1497 = 9'h1d8 == _T_538 ? _T_22_472 : _GEN_1496; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1498 = 9'h1d9 == _T_538 ? _T_22_473 : _GEN_1497; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1499 = 9'h1da == _T_538 ? _T_22_474 : _GEN_1498; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1500 = 9'h1db == _T_538 ? _T_22_475 : _GEN_1499; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1501 = 9'h1dc == _T_538 ? _T_22_476 : _GEN_1500; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1502 = 9'h1dd == _T_538 ? _T_22_477 : _GEN_1501; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1503 = 9'h1de == _T_538 ? _T_22_478 : _GEN_1502; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1504 = 9'h1df == _T_538 ? _T_22_479 : _GEN_1503; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1505 = 9'h1e0 == _T_538 ? _T_22_480 : _GEN_1504; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1506 = 9'h1e1 == _T_538 ? _T_22_481 : _GEN_1505; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1507 = 9'h1e2 == _T_538 ? _T_22_482 : _GEN_1506; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1508 = 9'h1e3 == _T_538 ? _T_22_483 : _GEN_1507; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1509 = 9'h1e4 == _T_538 ? _T_22_484 : _GEN_1508; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1510 = 9'h1e5 == _T_538 ? _T_22_485 : _GEN_1509; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1511 = 9'h1e6 == _T_538 ? _T_22_486 : _GEN_1510; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1512 = 9'h1e7 == _T_538 ? _T_22_487 : _GEN_1511; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1513 = 9'h1e8 == _T_538 ? _T_22_488 : _GEN_1512; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1514 = 9'h1e9 == _T_538 ? _T_22_489 : _GEN_1513; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1515 = 9'h1ea == _T_538 ? _T_22_490 : _GEN_1514; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1516 = 9'h1eb == _T_538 ? _T_22_491 : _GEN_1515; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1517 = 9'h1ec == _T_538 ? _T_22_492 : _GEN_1516; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1518 = 9'h1ed == _T_538 ? _T_22_493 : _GEN_1517; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1519 = 9'h1ee == _T_538 ? _T_22_494 : _GEN_1518; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1520 = 9'h1ef == _T_538 ? _T_22_495 : _GEN_1519; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1521 = 9'h1f0 == _T_538 ? _T_22_496 : _GEN_1520; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1522 = 9'h1f1 == _T_538 ? _T_22_497 : _GEN_1521; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1523 = 9'h1f2 == _T_538 ? _T_22_498 : _GEN_1522; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1524 = 9'h1f3 == _T_538 ? _T_22_499 : _GEN_1523; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1525 = 9'h1f4 == _T_538 ? _T_22_500 : _GEN_1524; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1526 = 9'h1f5 == _T_538 ? _T_22_501 : _GEN_1525; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1527 = 9'h1f6 == _T_538 ? _T_22_502 : _GEN_1526; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1528 = 9'h1f7 == _T_538 ? _T_22_503 : _GEN_1527; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1529 = 9'h1f8 == _T_538 ? _T_22_504 : _GEN_1528; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1530 = 9'h1f9 == _T_538 ? _T_22_505 : _GEN_1529; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1531 = 9'h1fa == _T_538 ? _T_22_506 : _GEN_1530; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1532 = 9'h1fb == _T_538 ? _T_22_507 : _GEN_1531; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1533 = 9'h1fc == _T_538 ? _T_22_508 : _GEN_1532; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1534 = 9'h1fd == _T_538 ? _T_22_509 : _GEN_1533; // @[nv_ram_rws.scala 36:13:@16.4]
  assign _GEN_1535 = 9'h1fe == _T_538 ? _T_22_510 : _GEN_1534; // @[nv_ram_rws.scala 36:13:@16.4]
  assign io_dout = 9'h1ff == _T_538 ? _T_22_511 : _GEN_1535; // @[nv_ram_rws.scala 36:13:@16.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {8{`RANDOM}};
  _T_22_0 = _RAND_0[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {8{`RANDOM}};
  _T_22_1 = _RAND_1[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {8{`RANDOM}};
  _T_22_2 = _RAND_2[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {8{`RANDOM}};
  _T_22_3 = _RAND_3[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {8{`RANDOM}};
  _T_22_4 = _RAND_4[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {8{`RANDOM}};
  _T_22_5 = _RAND_5[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {8{`RANDOM}};
  _T_22_6 = _RAND_6[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {8{`RANDOM}};
  _T_22_7 = _RAND_7[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {8{`RANDOM}};
  _T_22_8 = _RAND_8[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {8{`RANDOM}};
  _T_22_9 = _RAND_9[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {8{`RANDOM}};
  _T_22_10 = _RAND_10[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {8{`RANDOM}};
  _T_22_11 = _RAND_11[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {8{`RANDOM}};
  _T_22_12 = _RAND_12[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {8{`RANDOM}};
  _T_22_13 = _RAND_13[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {8{`RANDOM}};
  _T_22_14 = _RAND_14[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {8{`RANDOM}};
  _T_22_15 = _RAND_15[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {8{`RANDOM}};
  _T_22_16 = _RAND_16[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {8{`RANDOM}};
  _T_22_17 = _RAND_17[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {8{`RANDOM}};
  _T_22_18 = _RAND_18[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {8{`RANDOM}};
  _T_22_19 = _RAND_19[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {8{`RANDOM}};
  _T_22_20 = _RAND_20[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {8{`RANDOM}};
  _T_22_21 = _RAND_21[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {8{`RANDOM}};
  _T_22_22 = _RAND_22[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {8{`RANDOM}};
  _T_22_23 = _RAND_23[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {8{`RANDOM}};
  _T_22_24 = _RAND_24[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {8{`RANDOM}};
  _T_22_25 = _RAND_25[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {8{`RANDOM}};
  _T_22_26 = _RAND_26[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {8{`RANDOM}};
  _T_22_27 = _RAND_27[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {8{`RANDOM}};
  _T_22_28 = _RAND_28[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {8{`RANDOM}};
  _T_22_29 = _RAND_29[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {8{`RANDOM}};
  _T_22_30 = _RAND_30[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {8{`RANDOM}};
  _T_22_31 = _RAND_31[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {8{`RANDOM}};
  _T_22_32 = _RAND_32[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {8{`RANDOM}};
  _T_22_33 = _RAND_33[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {8{`RANDOM}};
  _T_22_34 = _RAND_34[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {8{`RANDOM}};
  _T_22_35 = _RAND_35[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {8{`RANDOM}};
  _T_22_36 = _RAND_36[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {8{`RANDOM}};
  _T_22_37 = _RAND_37[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {8{`RANDOM}};
  _T_22_38 = _RAND_38[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {8{`RANDOM}};
  _T_22_39 = _RAND_39[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {8{`RANDOM}};
  _T_22_40 = _RAND_40[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {8{`RANDOM}};
  _T_22_41 = _RAND_41[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {8{`RANDOM}};
  _T_22_42 = _RAND_42[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {8{`RANDOM}};
  _T_22_43 = _RAND_43[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {8{`RANDOM}};
  _T_22_44 = _RAND_44[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {8{`RANDOM}};
  _T_22_45 = _RAND_45[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {8{`RANDOM}};
  _T_22_46 = _RAND_46[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {8{`RANDOM}};
  _T_22_47 = _RAND_47[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {8{`RANDOM}};
  _T_22_48 = _RAND_48[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {8{`RANDOM}};
  _T_22_49 = _RAND_49[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {8{`RANDOM}};
  _T_22_50 = _RAND_50[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {8{`RANDOM}};
  _T_22_51 = _RAND_51[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {8{`RANDOM}};
  _T_22_52 = _RAND_52[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {8{`RANDOM}};
  _T_22_53 = _RAND_53[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {8{`RANDOM}};
  _T_22_54 = _RAND_54[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {8{`RANDOM}};
  _T_22_55 = _RAND_55[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {8{`RANDOM}};
  _T_22_56 = _RAND_56[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {8{`RANDOM}};
  _T_22_57 = _RAND_57[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {8{`RANDOM}};
  _T_22_58 = _RAND_58[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {8{`RANDOM}};
  _T_22_59 = _RAND_59[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {8{`RANDOM}};
  _T_22_60 = _RAND_60[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {8{`RANDOM}};
  _T_22_61 = _RAND_61[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {8{`RANDOM}};
  _T_22_62 = _RAND_62[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {8{`RANDOM}};
  _T_22_63 = _RAND_63[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {8{`RANDOM}};
  _T_22_64 = _RAND_64[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {8{`RANDOM}};
  _T_22_65 = _RAND_65[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {8{`RANDOM}};
  _T_22_66 = _RAND_66[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {8{`RANDOM}};
  _T_22_67 = _RAND_67[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {8{`RANDOM}};
  _T_22_68 = _RAND_68[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {8{`RANDOM}};
  _T_22_69 = _RAND_69[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {8{`RANDOM}};
  _T_22_70 = _RAND_70[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {8{`RANDOM}};
  _T_22_71 = _RAND_71[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {8{`RANDOM}};
  _T_22_72 = _RAND_72[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {8{`RANDOM}};
  _T_22_73 = _RAND_73[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {8{`RANDOM}};
  _T_22_74 = _RAND_74[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {8{`RANDOM}};
  _T_22_75 = _RAND_75[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {8{`RANDOM}};
  _T_22_76 = _RAND_76[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {8{`RANDOM}};
  _T_22_77 = _RAND_77[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {8{`RANDOM}};
  _T_22_78 = _RAND_78[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {8{`RANDOM}};
  _T_22_79 = _RAND_79[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {8{`RANDOM}};
  _T_22_80 = _RAND_80[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {8{`RANDOM}};
  _T_22_81 = _RAND_81[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {8{`RANDOM}};
  _T_22_82 = _RAND_82[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {8{`RANDOM}};
  _T_22_83 = _RAND_83[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {8{`RANDOM}};
  _T_22_84 = _RAND_84[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {8{`RANDOM}};
  _T_22_85 = _RAND_85[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {8{`RANDOM}};
  _T_22_86 = _RAND_86[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {8{`RANDOM}};
  _T_22_87 = _RAND_87[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {8{`RANDOM}};
  _T_22_88 = _RAND_88[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {8{`RANDOM}};
  _T_22_89 = _RAND_89[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {8{`RANDOM}};
  _T_22_90 = _RAND_90[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {8{`RANDOM}};
  _T_22_91 = _RAND_91[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {8{`RANDOM}};
  _T_22_92 = _RAND_92[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {8{`RANDOM}};
  _T_22_93 = _RAND_93[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {8{`RANDOM}};
  _T_22_94 = _RAND_94[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {8{`RANDOM}};
  _T_22_95 = _RAND_95[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {8{`RANDOM}};
  _T_22_96 = _RAND_96[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {8{`RANDOM}};
  _T_22_97 = _RAND_97[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {8{`RANDOM}};
  _T_22_98 = _RAND_98[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {8{`RANDOM}};
  _T_22_99 = _RAND_99[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {8{`RANDOM}};
  _T_22_100 = _RAND_100[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {8{`RANDOM}};
  _T_22_101 = _RAND_101[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {8{`RANDOM}};
  _T_22_102 = _RAND_102[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {8{`RANDOM}};
  _T_22_103 = _RAND_103[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {8{`RANDOM}};
  _T_22_104 = _RAND_104[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {8{`RANDOM}};
  _T_22_105 = _RAND_105[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {8{`RANDOM}};
  _T_22_106 = _RAND_106[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {8{`RANDOM}};
  _T_22_107 = _RAND_107[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {8{`RANDOM}};
  _T_22_108 = _RAND_108[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {8{`RANDOM}};
  _T_22_109 = _RAND_109[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {8{`RANDOM}};
  _T_22_110 = _RAND_110[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {8{`RANDOM}};
  _T_22_111 = _RAND_111[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {8{`RANDOM}};
  _T_22_112 = _RAND_112[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {8{`RANDOM}};
  _T_22_113 = _RAND_113[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {8{`RANDOM}};
  _T_22_114 = _RAND_114[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {8{`RANDOM}};
  _T_22_115 = _RAND_115[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {8{`RANDOM}};
  _T_22_116 = _RAND_116[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {8{`RANDOM}};
  _T_22_117 = _RAND_117[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {8{`RANDOM}};
  _T_22_118 = _RAND_118[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {8{`RANDOM}};
  _T_22_119 = _RAND_119[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {8{`RANDOM}};
  _T_22_120 = _RAND_120[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {8{`RANDOM}};
  _T_22_121 = _RAND_121[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {8{`RANDOM}};
  _T_22_122 = _RAND_122[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {8{`RANDOM}};
  _T_22_123 = _RAND_123[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {8{`RANDOM}};
  _T_22_124 = _RAND_124[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {8{`RANDOM}};
  _T_22_125 = _RAND_125[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {8{`RANDOM}};
  _T_22_126 = _RAND_126[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {8{`RANDOM}};
  _T_22_127 = _RAND_127[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {8{`RANDOM}};
  _T_22_128 = _RAND_128[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {8{`RANDOM}};
  _T_22_129 = _RAND_129[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {8{`RANDOM}};
  _T_22_130 = _RAND_130[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {8{`RANDOM}};
  _T_22_131 = _RAND_131[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {8{`RANDOM}};
  _T_22_132 = _RAND_132[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {8{`RANDOM}};
  _T_22_133 = _RAND_133[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {8{`RANDOM}};
  _T_22_134 = _RAND_134[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {8{`RANDOM}};
  _T_22_135 = _RAND_135[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {8{`RANDOM}};
  _T_22_136 = _RAND_136[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {8{`RANDOM}};
  _T_22_137 = _RAND_137[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {8{`RANDOM}};
  _T_22_138 = _RAND_138[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {8{`RANDOM}};
  _T_22_139 = _RAND_139[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {8{`RANDOM}};
  _T_22_140 = _RAND_140[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {8{`RANDOM}};
  _T_22_141 = _RAND_141[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {8{`RANDOM}};
  _T_22_142 = _RAND_142[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {8{`RANDOM}};
  _T_22_143 = _RAND_143[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {8{`RANDOM}};
  _T_22_144 = _RAND_144[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {8{`RANDOM}};
  _T_22_145 = _RAND_145[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {8{`RANDOM}};
  _T_22_146 = _RAND_146[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {8{`RANDOM}};
  _T_22_147 = _RAND_147[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {8{`RANDOM}};
  _T_22_148 = _RAND_148[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {8{`RANDOM}};
  _T_22_149 = _RAND_149[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {8{`RANDOM}};
  _T_22_150 = _RAND_150[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {8{`RANDOM}};
  _T_22_151 = _RAND_151[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {8{`RANDOM}};
  _T_22_152 = _RAND_152[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {8{`RANDOM}};
  _T_22_153 = _RAND_153[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {8{`RANDOM}};
  _T_22_154 = _RAND_154[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {8{`RANDOM}};
  _T_22_155 = _RAND_155[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {8{`RANDOM}};
  _T_22_156 = _RAND_156[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {8{`RANDOM}};
  _T_22_157 = _RAND_157[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {8{`RANDOM}};
  _T_22_158 = _RAND_158[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {8{`RANDOM}};
  _T_22_159 = _RAND_159[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {8{`RANDOM}};
  _T_22_160 = _RAND_160[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {8{`RANDOM}};
  _T_22_161 = _RAND_161[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {8{`RANDOM}};
  _T_22_162 = _RAND_162[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {8{`RANDOM}};
  _T_22_163 = _RAND_163[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {8{`RANDOM}};
  _T_22_164 = _RAND_164[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {8{`RANDOM}};
  _T_22_165 = _RAND_165[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {8{`RANDOM}};
  _T_22_166 = _RAND_166[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {8{`RANDOM}};
  _T_22_167 = _RAND_167[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {8{`RANDOM}};
  _T_22_168 = _RAND_168[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {8{`RANDOM}};
  _T_22_169 = _RAND_169[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {8{`RANDOM}};
  _T_22_170 = _RAND_170[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {8{`RANDOM}};
  _T_22_171 = _RAND_171[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {8{`RANDOM}};
  _T_22_172 = _RAND_172[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {8{`RANDOM}};
  _T_22_173 = _RAND_173[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {8{`RANDOM}};
  _T_22_174 = _RAND_174[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {8{`RANDOM}};
  _T_22_175 = _RAND_175[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {8{`RANDOM}};
  _T_22_176 = _RAND_176[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {8{`RANDOM}};
  _T_22_177 = _RAND_177[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {8{`RANDOM}};
  _T_22_178 = _RAND_178[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {8{`RANDOM}};
  _T_22_179 = _RAND_179[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {8{`RANDOM}};
  _T_22_180 = _RAND_180[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {8{`RANDOM}};
  _T_22_181 = _RAND_181[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {8{`RANDOM}};
  _T_22_182 = _RAND_182[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {8{`RANDOM}};
  _T_22_183 = _RAND_183[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {8{`RANDOM}};
  _T_22_184 = _RAND_184[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {8{`RANDOM}};
  _T_22_185 = _RAND_185[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {8{`RANDOM}};
  _T_22_186 = _RAND_186[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {8{`RANDOM}};
  _T_22_187 = _RAND_187[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {8{`RANDOM}};
  _T_22_188 = _RAND_188[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {8{`RANDOM}};
  _T_22_189 = _RAND_189[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {8{`RANDOM}};
  _T_22_190 = _RAND_190[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {8{`RANDOM}};
  _T_22_191 = _RAND_191[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {8{`RANDOM}};
  _T_22_192 = _RAND_192[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {8{`RANDOM}};
  _T_22_193 = _RAND_193[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {8{`RANDOM}};
  _T_22_194 = _RAND_194[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {8{`RANDOM}};
  _T_22_195 = _RAND_195[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {8{`RANDOM}};
  _T_22_196 = _RAND_196[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {8{`RANDOM}};
  _T_22_197 = _RAND_197[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {8{`RANDOM}};
  _T_22_198 = _RAND_198[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {8{`RANDOM}};
  _T_22_199 = _RAND_199[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {8{`RANDOM}};
  _T_22_200 = _RAND_200[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {8{`RANDOM}};
  _T_22_201 = _RAND_201[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {8{`RANDOM}};
  _T_22_202 = _RAND_202[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {8{`RANDOM}};
  _T_22_203 = _RAND_203[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {8{`RANDOM}};
  _T_22_204 = _RAND_204[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {8{`RANDOM}};
  _T_22_205 = _RAND_205[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {8{`RANDOM}};
  _T_22_206 = _RAND_206[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {8{`RANDOM}};
  _T_22_207 = _RAND_207[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {8{`RANDOM}};
  _T_22_208 = _RAND_208[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {8{`RANDOM}};
  _T_22_209 = _RAND_209[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {8{`RANDOM}};
  _T_22_210 = _RAND_210[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {8{`RANDOM}};
  _T_22_211 = _RAND_211[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {8{`RANDOM}};
  _T_22_212 = _RAND_212[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {8{`RANDOM}};
  _T_22_213 = _RAND_213[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {8{`RANDOM}};
  _T_22_214 = _RAND_214[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {8{`RANDOM}};
  _T_22_215 = _RAND_215[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {8{`RANDOM}};
  _T_22_216 = _RAND_216[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {8{`RANDOM}};
  _T_22_217 = _RAND_217[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {8{`RANDOM}};
  _T_22_218 = _RAND_218[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {8{`RANDOM}};
  _T_22_219 = _RAND_219[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {8{`RANDOM}};
  _T_22_220 = _RAND_220[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {8{`RANDOM}};
  _T_22_221 = _RAND_221[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {8{`RANDOM}};
  _T_22_222 = _RAND_222[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {8{`RANDOM}};
  _T_22_223 = _RAND_223[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {8{`RANDOM}};
  _T_22_224 = _RAND_224[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {8{`RANDOM}};
  _T_22_225 = _RAND_225[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {8{`RANDOM}};
  _T_22_226 = _RAND_226[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {8{`RANDOM}};
  _T_22_227 = _RAND_227[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {8{`RANDOM}};
  _T_22_228 = _RAND_228[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {8{`RANDOM}};
  _T_22_229 = _RAND_229[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {8{`RANDOM}};
  _T_22_230 = _RAND_230[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {8{`RANDOM}};
  _T_22_231 = _RAND_231[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {8{`RANDOM}};
  _T_22_232 = _RAND_232[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {8{`RANDOM}};
  _T_22_233 = _RAND_233[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {8{`RANDOM}};
  _T_22_234 = _RAND_234[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {8{`RANDOM}};
  _T_22_235 = _RAND_235[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {8{`RANDOM}};
  _T_22_236 = _RAND_236[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {8{`RANDOM}};
  _T_22_237 = _RAND_237[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {8{`RANDOM}};
  _T_22_238 = _RAND_238[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {8{`RANDOM}};
  _T_22_239 = _RAND_239[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {8{`RANDOM}};
  _T_22_240 = _RAND_240[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {8{`RANDOM}};
  _T_22_241 = _RAND_241[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {8{`RANDOM}};
  _T_22_242 = _RAND_242[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {8{`RANDOM}};
  _T_22_243 = _RAND_243[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {8{`RANDOM}};
  _T_22_244 = _RAND_244[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {8{`RANDOM}};
  _T_22_245 = _RAND_245[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {8{`RANDOM}};
  _T_22_246 = _RAND_246[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {8{`RANDOM}};
  _T_22_247 = _RAND_247[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {8{`RANDOM}};
  _T_22_248 = _RAND_248[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {8{`RANDOM}};
  _T_22_249 = _RAND_249[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {8{`RANDOM}};
  _T_22_250 = _RAND_250[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {8{`RANDOM}};
  _T_22_251 = _RAND_251[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {8{`RANDOM}};
  _T_22_252 = _RAND_252[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {8{`RANDOM}};
  _T_22_253 = _RAND_253[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {8{`RANDOM}};
  _T_22_254 = _RAND_254[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {8{`RANDOM}};
  _T_22_255 = _RAND_255[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {8{`RANDOM}};
  _T_22_256 = _RAND_256[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {8{`RANDOM}};
  _T_22_257 = _RAND_257[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {8{`RANDOM}};
  _T_22_258 = _RAND_258[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {8{`RANDOM}};
  _T_22_259 = _RAND_259[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {8{`RANDOM}};
  _T_22_260 = _RAND_260[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {8{`RANDOM}};
  _T_22_261 = _RAND_261[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {8{`RANDOM}};
  _T_22_262 = _RAND_262[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {8{`RANDOM}};
  _T_22_263 = _RAND_263[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {8{`RANDOM}};
  _T_22_264 = _RAND_264[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {8{`RANDOM}};
  _T_22_265 = _RAND_265[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {8{`RANDOM}};
  _T_22_266 = _RAND_266[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {8{`RANDOM}};
  _T_22_267 = _RAND_267[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {8{`RANDOM}};
  _T_22_268 = _RAND_268[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {8{`RANDOM}};
  _T_22_269 = _RAND_269[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {8{`RANDOM}};
  _T_22_270 = _RAND_270[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {8{`RANDOM}};
  _T_22_271 = _RAND_271[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {8{`RANDOM}};
  _T_22_272 = _RAND_272[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {8{`RANDOM}};
  _T_22_273 = _RAND_273[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {8{`RANDOM}};
  _T_22_274 = _RAND_274[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {8{`RANDOM}};
  _T_22_275 = _RAND_275[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {8{`RANDOM}};
  _T_22_276 = _RAND_276[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {8{`RANDOM}};
  _T_22_277 = _RAND_277[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {8{`RANDOM}};
  _T_22_278 = _RAND_278[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {8{`RANDOM}};
  _T_22_279 = _RAND_279[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {8{`RANDOM}};
  _T_22_280 = _RAND_280[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {8{`RANDOM}};
  _T_22_281 = _RAND_281[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {8{`RANDOM}};
  _T_22_282 = _RAND_282[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {8{`RANDOM}};
  _T_22_283 = _RAND_283[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {8{`RANDOM}};
  _T_22_284 = _RAND_284[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {8{`RANDOM}};
  _T_22_285 = _RAND_285[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {8{`RANDOM}};
  _T_22_286 = _RAND_286[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {8{`RANDOM}};
  _T_22_287 = _RAND_287[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {8{`RANDOM}};
  _T_22_288 = _RAND_288[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {8{`RANDOM}};
  _T_22_289 = _RAND_289[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {8{`RANDOM}};
  _T_22_290 = _RAND_290[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {8{`RANDOM}};
  _T_22_291 = _RAND_291[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {8{`RANDOM}};
  _T_22_292 = _RAND_292[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {8{`RANDOM}};
  _T_22_293 = _RAND_293[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {8{`RANDOM}};
  _T_22_294 = _RAND_294[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {8{`RANDOM}};
  _T_22_295 = _RAND_295[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {8{`RANDOM}};
  _T_22_296 = _RAND_296[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {8{`RANDOM}};
  _T_22_297 = _RAND_297[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {8{`RANDOM}};
  _T_22_298 = _RAND_298[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {8{`RANDOM}};
  _T_22_299 = _RAND_299[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {8{`RANDOM}};
  _T_22_300 = _RAND_300[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {8{`RANDOM}};
  _T_22_301 = _RAND_301[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {8{`RANDOM}};
  _T_22_302 = _RAND_302[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {8{`RANDOM}};
  _T_22_303 = _RAND_303[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {8{`RANDOM}};
  _T_22_304 = _RAND_304[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {8{`RANDOM}};
  _T_22_305 = _RAND_305[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {8{`RANDOM}};
  _T_22_306 = _RAND_306[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {8{`RANDOM}};
  _T_22_307 = _RAND_307[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {8{`RANDOM}};
  _T_22_308 = _RAND_308[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {8{`RANDOM}};
  _T_22_309 = _RAND_309[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {8{`RANDOM}};
  _T_22_310 = _RAND_310[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {8{`RANDOM}};
  _T_22_311 = _RAND_311[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {8{`RANDOM}};
  _T_22_312 = _RAND_312[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {8{`RANDOM}};
  _T_22_313 = _RAND_313[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {8{`RANDOM}};
  _T_22_314 = _RAND_314[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {8{`RANDOM}};
  _T_22_315 = _RAND_315[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {8{`RANDOM}};
  _T_22_316 = _RAND_316[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {8{`RANDOM}};
  _T_22_317 = _RAND_317[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {8{`RANDOM}};
  _T_22_318 = _RAND_318[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {8{`RANDOM}};
  _T_22_319 = _RAND_319[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {8{`RANDOM}};
  _T_22_320 = _RAND_320[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {8{`RANDOM}};
  _T_22_321 = _RAND_321[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {8{`RANDOM}};
  _T_22_322 = _RAND_322[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {8{`RANDOM}};
  _T_22_323 = _RAND_323[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {8{`RANDOM}};
  _T_22_324 = _RAND_324[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {8{`RANDOM}};
  _T_22_325 = _RAND_325[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {8{`RANDOM}};
  _T_22_326 = _RAND_326[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {8{`RANDOM}};
  _T_22_327 = _RAND_327[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {8{`RANDOM}};
  _T_22_328 = _RAND_328[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {8{`RANDOM}};
  _T_22_329 = _RAND_329[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {8{`RANDOM}};
  _T_22_330 = _RAND_330[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {8{`RANDOM}};
  _T_22_331 = _RAND_331[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {8{`RANDOM}};
  _T_22_332 = _RAND_332[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {8{`RANDOM}};
  _T_22_333 = _RAND_333[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {8{`RANDOM}};
  _T_22_334 = _RAND_334[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {8{`RANDOM}};
  _T_22_335 = _RAND_335[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {8{`RANDOM}};
  _T_22_336 = _RAND_336[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {8{`RANDOM}};
  _T_22_337 = _RAND_337[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {8{`RANDOM}};
  _T_22_338 = _RAND_338[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {8{`RANDOM}};
  _T_22_339 = _RAND_339[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {8{`RANDOM}};
  _T_22_340 = _RAND_340[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {8{`RANDOM}};
  _T_22_341 = _RAND_341[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {8{`RANDOM}};
  _T_22_342 = _RAND_342[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {8{`RANDOM}};
  _T_22_343 = _RAND_343[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {8{`RANDOM}};
  _T_22_344 = _RAND_344[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {8{`RANDOM}};
  _T_22_345 = _RAND_345[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {8{`RANDOM}};
  _T_22_346 = _RAND_346[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {8{`RANDOM}};
  _T_22_347 = _RAND_347[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {8{`RANDOM}};
  _T_22_348 = _RAND_348[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {8{`RANDOM}};
  _T_22_349 = _RAND_349[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {8{`RANDOM}};
  _T_22_350 = _RAND_350[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {8{`RANDOM}};
  _T_22_351 = _RAND_351[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {8{`RANDOM}};
  _T_22_352 = _RAND_352[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {8{`RANDOM}};
  _T_22_353 = _RAND_353[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {8{`RANDOM}};
  _T_22_354 = _RAND_354[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {8{`RANDOM}};
  _T_22_355 = _RAND_355[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {8{`RANDOM}};
  _T_22_356 = _RAND_356[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {8{`RANDOM}};
  _T_22_357 = _RAND_357[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {8{`RANDOM}};
  _T_22_358 = _RAND_358[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {8{`RANDOM}};
  _T_22_359 = _RAND_359[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {8{`RANDOM}};
  _T_22_360 = _RAND_360[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {8{`RANDOM}};
  _T_22_361 = _RAND_361[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {8{`RANDOM}};
  _T_22_362 = _RAND_362[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {8{`RANDOM}};
  _T_22_363 = _RAND_363[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {8{`RANDOM}};
  _T_22_364 = _RAND_364[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {8{`RANDOM}};
  _T_22_365 = _RAND_365[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {8{`RANDOM}};
  _T_22_366 = _RAND_366[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {8{`RANDOM}};
  _T_22_367 = _RAND_367[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {8{`RANDOM}};
  _T_22_368 = _RAND_368[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {8{`RANDOM}};
  _T_22_369 = _RAND_369[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {8{`RANDOM}};
  _T_22_370 = _RAND_370[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {8{`RANDOM}};
  _T_22_371 = _RAND_371[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {8{`RANDOM}};
  _T_22_372 = _RAND_372[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {8{`RANDOM}};
  _T_22_373 = _RAND_373[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {8{`RANDOM}};
  _T_22_374 = _RAND_374[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {8{`RANDOM}};
  _T_22_375 = _RAND_375[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {8{`RANDOM}};
  _T_22_376 = _RAND_376[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {8{`RANDOM}};
  _T_22_377 = _RAND_377[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {8{`RANDOM}};
  _T_22_378 = _RAND_378[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {8{`RANDOM}};
  _T_22_379 = _RAND_379[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {8{`RANDOM}};
  _T_22_380 = _RAND_380[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {8{`RANDOM}};
  _T_22_381 = _RAND_381[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {8{`RANDOM}};
  _T_22_382 = _RAND_382[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {8{`RANDOM}};
  _T_22_383 = _RAND_383[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {8{`RANDOM}};
  _T_22_384 = _RAND_384[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {8{`RANDOM}};
  _T_22_385 = _RAND_385[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {8{`RANDOM}};
  _T_22_386 = _RAND_386[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {8{`RANDOM}};
  _T_22_387 = _RAND_387[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {8{`RANDOM}};
  _T_22_388 = _RAND_388[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {8{`RANDOM}};
  _T_22_389 = _RAND_389[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {8{`RANDOM}};
  _T_22_390 = _RAND_390[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {8{`RANDOM}};
  _T_22_391 = _RAND_391[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {8{`RANDOM}};
  _T_22_392 = _RAND_392[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {8{`RANDOM}};
  _T_22_393 = _RAND_393[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {8{`RANDOM}};
  _T_22_394 = _RAND_394[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {8{`RANDOM}};
  _T_22_395 = _RAND_395[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {8{`RANDOM}};
  _T_22_396 = _RAND_396[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {8{`RANDOM}};
  _T_22_397 = _RAND_397[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {8{`RANDOM}};
  _T_22_398 = _RAND_398[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {8{`RANDOM}};
  _T_22_399 = _RAND_399[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {8{`RANDOM}};
  _T_22_400 = _RAND_400[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {8{`RANDOM}};
  _T_22_401 = _RAND_401[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {8{`RANDOM}};
  _T_22_402 = _RAND_402[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {8{`RANDOM}};
  _T_22_403 = _RAND_403[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {8{`RANDOM}};
  _T_22_404 = _RAND_404[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {8{`RANDOM}};
  _T_22_405 = _RAND_405[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {8{`RANDOM}};
  _T_22_406 = _RAND_406[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {8{`RANDOM}};
  _T_22_407 = _RAND_407[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {8{`RANDOM}};
  _T_22_408 = _RAND_408[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {8{`RANDOM}};
  _T_22_409 = _RAND_409[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {8{`RANDOM}};
  _T_22_410 = _RAND_410[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {8{`RANDOM}};
  _T_22_411 = _RAND_411[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {8{`RANDOM}};
  _T_22_412 = _RAND_412[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {8{`RANDOM}};
  _T_22_413 = _RAND_413[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {8{`RANDOM}};
  _T_22_414 = _RAND_414[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {8{`RANDOM}};
  _T_22_415 = _RAND_415[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {8{`RANDOM}};
  _T_22_416 = _RAND_416[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {8{`RANDOM}};
  _T_22_417 = _RAND_417[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {8{`RANDOM}};
  _T_22_418 = _RAND_418[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {8{`RANDOM}};
  _T_22_419 = _RAND_419[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {8{`RANDOM}};
  _T_22_420 = _RAND_420[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {8{`RANDOM}};
  _T_22_421 = _RAND_421[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {8{`RANDOM}};
  _T_22_422 = _RAND_422[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {8{`RANDOM}};
  _T_22_423 = _RAND_423[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {8{`RANDOM}};
  _T_22_424 = _RAND_424[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {8{`RANDOM}};
  _T_22_425 = _RAND_425[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {8{`RANDOM}};
  _T_22_426 = _RAND_426[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {8{`RANDOM}};
  _T_22_427 = _RAND_427[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {8{`RANDOM}};
  _T_22_428 = _RAND_428[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {8{`RANDOM}};
  _T_22_429 = _RAND_429[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {8{`RANDOM}};
  _T_22_430 = _RAND_430[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {8{`RANDOM}};
  _T_22_431 = _RAND_431[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {8{`RANDOM}};
  _T_22_432 = _RAND_432[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {8{`RANDOM}};
  _T_22_433 = _RAND_433[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {8{`RANDOM}};
  _T_22_434 = _RAND_434[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {8{`RANDOM}};
  _T_22_435 = _RAND_435[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {8{`RANDOM}};
  _T_22_436 = _RAND_436[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {8{`RANDOM}};
  _T_22_437 = _RAND_437[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {8{`RANDOM}};
  _T_22_438 = _RAND_438[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {8{`RANDOM}};
  _T_22_439 = _RAND_439[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {8{`RANDOM}};
  _T_22_440 = _RAND_440[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {8{`RANDOM}};
  _T_22_441 = _RAND_441[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {8{`RANDOM}};
  _T_22_442 = _RAND_442[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {8{`RANDOM}};
  _T_22_443 = _RAND_443[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {8{`RANDOM}};
  _T_22_444 = _RAND_444[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {8{`RANDOM}};
  _T_22_445 = _RAND_445[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {8{`RANDOM}};
  _T_22_446 = _RAND_446[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {8{`RANDOM}};
  _T_22_447 = _RAND_447[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {8{`RANDOM}};
  _T_22_448 = _RAND_448[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {8{`RANDOM}};
  _T_22_449 = _RAND_449[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {8{`RANDOM}};
  _T_22_450 = _RAND_450[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {8{`RANDOM}};
  _T_22_451 = _RAND_451[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {8{`RANDOM}};
  _T_22_452 = _RAND_452[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {8{`RANDOM}};
  _T_22_453 = _RAND_453[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {8{`RANDOM}};
  _T_22_454 = _RAND_454[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {8{`RANDOM}};
  _T_22_455 = _RAND_455[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {8{`RANDOM}};
  _T_22_456 = _RAND_456[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {8{`RANDOM}};
  _T_22_457 = _RAND_457[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {8{`RANDOM}};
  _T_22_458 = _RAND_458[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {8{`RANDOM}};
  _T_22_459 = _RAND_459[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {8{`RANDOM}};
  _T_22_460 = _RAND_460[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {8{`RANDOM}};
  _T_22_461 = _RAND_461[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {8{`RANDOM}};
  _T_22_462 = _RAND_462[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {8{`RANDOM}};
  _T_22_463 = _RAND_463[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {8{`RANDOM}};
  _T_22_464 = _RAND_464[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {8{`RANDOM}};
  _T_22_465 = _RAND_465[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {8{`RANDOM}};
  _T_22_466 = _RAND_466[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {8{`RANDOM}};
  _T_22_467 = _RAND_467[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {8{`RANDOM}};
  _T_22_468 = _RAND_468[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {8{`RANDOM}};
  _T_22_469 = _RAND_469[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {8{`RANDOM}};
  _T_22_470 = _RAND_470[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {8{`RANDOM}};
  _T_22_471 = _RAND_471[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {8{`RANDOM}};
  _T_22_472 = _RAND_472[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {8{`RANDOM}};
  _T_22_473 = _RAND_473[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {8{`RANDOM}};
  _T_22_474 = _RAND_474[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {8{`RANDOM}};
  _T_22_475 = _RAND_475[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {8{`RANDOM}};
  _T_22_476 = _RAND_476[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {8{`RANDOM}};
  _T_22_477 = _RAND_477[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {8{`RANDOM}};
  _T_22_478 = _RAND_478[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {8{`RANDOM}};
  _T_22_479 = _RAND_479[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {8{`RANDOM}};
  _T_22_480 = _RAND_480[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {8{`RANDOM}};
  _T_22_481 = _RAND_481[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {8{`RANDOM}};
  _T_22_482 = _RAND_482[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {8{`RANDOM}};
  _T_22_483 = _RAND_483[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {8{`RANDOM}};
  _T_22_484 = _RAND_484[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {8{`RANDOM}};
  _T_22_485 = _RAND_485[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {8{`RANDOM}};
  _T_22_486 = _RAND_486[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {8{`RANDOM}};
  _T_22_487 = _RAND_487[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {8{`RANDOM}};
  _T_22_488 = _RAND_488[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {8{`RANDOM}};
  _T_22_489 = _RAND_489[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {8{`RANDOM}};
  _T_22_490 = _RAND_490[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {8{`RANDOM}};
  _T_22_491 = _RAND_491[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {8{`RANDOM}};
  _T_22_492 = _RAND_492[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {8{`RANDOM}};
  _T_22_493 = _RAND_493[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {8{`RANDOM}};
  _T_22_494 = _RAND_494[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {8{`RANDOM}};
  _T_22_495 = _RAND_495[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {8{`RANDOM}};
  _T_22_496 = _RAND_496[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {8{`RANDOM}};
  _T_22_497 = _RAND_497[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {8{`RANDOM}};
  _T_22_498 = _RAND_498[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {8{`RANDOM}};
  _T_22_499 = _RAND_499[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {8{`RANDOM}};
  _T_22_500 = _RAND_500[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {8{`RANDOM}};
  _T_22_501 = _RAND_501[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {8{`RANDOM}};
  _T_22_502 = _RAND_502[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {8{`RANDOM}};
  _T_22_503 = _RAND_503[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {8{`RANDOM}};
  _T_22_504 = _RAND_504[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {8{`RANDOM}};
  _T_22_505 = _RAND_505[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {8{`RANDOM}};
  _T_22_506 = _RAND_506[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {8{`RANDOM}};
  _T_22_507 = _RAND_507[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {8{`RANDOM}};
  _T_22_508 = _RAND_508[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {8{`RANDOM}};
  _T_22_509 = _RAND_509[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {8{`RANDOM}};
  _T_22_510 = _RAND_510[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {8{`RANDOM}};
  _T_22_511 = _RAND_511[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_538 = _RAND_512[8:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_clk) begin
    if (io_we) begin
      if (9'h0 == io_wa) begin
        _T_22_0 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1 == io_wa) begin
        _T_22_1 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h2 == io_wa) begin
        _T_22_2 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h3 == io_wa) begin
        _T_22_3 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h4 == io_wa) begin
        _T_22_4 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h5 == io_wa) begin
        _T_22_5 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h6 == io_wa) begin
        _T_22_6 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h7 == io_wa) begin
        _T_22_7 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h8 == io_wa) begin
        _T_22_8 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h9 == io_wa) begin
        _T_22_9 <= io_di;
      end
    end
    if (io_we) begin
      if (9'ha == io_wa) begin
        _T_22_10 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hb == io_wa) begin
        _T_22_11 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hc == io_wa) begin
        _T_22_12 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hd == io_wa) begin
        _T_22_13 <= io_di;
      end
    end
    if (io_we) begin
      if (9'he == io_wa) begin
        _T_22_14 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hf == io_wa) begin
        _T_22_15 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h10 == io_wa) begin
        _T_22_16 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h11 == io_wa) begin
        _T_22_17 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h12 == io_wa) begin
        _T_22_18 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h13 == io_wa) begin
        _T_22_19 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h14 == io_wa) begin
        _T_22_20 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h15 == io_wa) begin
        _T_22_21 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h16 == io_wa) begin
        _T_22_22 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h17 == io_wa) begin
        _T_22_23 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h18 == io_wa) begin
        _T_22_24 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h19 == io_wa) begin
        _T_22_25 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1a == io_wa) begin
        _T_22_26 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1b == io_wa) begin
        _T_22_27 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1c == io_wa) begin
        _T_22_28 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1d == io_wa) begin
        _T_22_29 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1e == io_wa) begin
        _T_22_30 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1f == io_wa) begin
        _T_22_31 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h20 == io_wa) begin
        _T_22_32 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h21 == io_wa) begin
        _T_22_33 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h22 == io_wa) begin
        _T_22_34 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h23 == io_wa) begin
        _T_22_35 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h24 == io_wa) begin
        _T_22_36 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h25 == io_wa) begin
        _T_22_37 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h26 == io_wa) begin
        _T_22_38 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h27 == io_wa) begin
        _T_22_39 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h28 == io_wa) begin
        _T_22_40 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h29 == io_wa) begin
        _T_22_41 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h2a == io_wa) begin
        _T_22_42 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h2b == io_wa) begin
        _T_22_43 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h2c == io_wa) begin
        _T_22_44 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h2d == io_wa) begin
        _T_22_45 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h2e == io_wa) begin
        _T_22_46 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h2f == io_wa) begin
        _T_22_47 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h30 == io_wa) begin
        _T_22_48 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h31 == io_wa) begin
        _T_22_49 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h32 == io_wa) begin
        _T_22_50 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h33 == io_wa) begin
        _T_22_51 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h34 == io_wa) begin
        _T_22_52 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h35 == io_wa) begin
        _T_22_53 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h36 == io_wa) begin
        _T_22_54 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h37 == io_wa) begin
        _T_22_55 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h38 == io_wa) begin
        _T_22_56 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h39 == io_wa) begin
        _T_22_57 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h3a == io_wa) begin
        _T_22_58 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h3b == io_wa) begin
        _T_22_59 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h3c == io_wa) begin
        _T_22_60 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h3d == io_wa) begin
        _T_22_61 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h3e == io_wa) begin
        _T_22_62 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h3f == io_wa) begin
        _T_22_63 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h40 == io_wa) begin
        _T_22_64 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h41 == io_wa) begin
        _T_22_65 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h42 == io_wa) begin
        _T_22_66 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h43 == io_wa) begin
        _T_22_67 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h44 == io_wa) begin
        _T_22_68 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h45 == io_wa) begin
        _T_22_69 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h46 == io_wa) begin
        _T_22_70 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h47 == io_wa) begin
        _T_22_71 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h48 == io_wa) begin
        _T_22_72 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h49 == io_wa) begin
        _T_22_73 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h4a == io_wa) begin
        _T_22_74 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h4b == io_wa) begin
        _T_22_75 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h4c == io_wa) begin
        _T_22_76 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h4d == io_wa) begin
        _T_22_77 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h4e == io_wa) begin
        _T_22_78 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h4f == io_wa) begin
        _T_22_79 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h50 == io_wa) begin
        _T_22_80 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h51 == io_wa) begin
        _T_22_81 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h52 == io_wa) begin
        _T_22_82 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h53 == io_wa) begin
        _T_22_83 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h54 == io_wa) begin
        _T_22_84 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h55 == io_wa) begin
        _T_22_85 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h56 == io_wa) begin
        _T_22_86 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h57 == io_wa) begin
        _T_22_87 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h58 == io_wa) begin
        _T_22_88 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h59 == io_wa) begin
        _T_22_89 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h5a == io_wa) begin
        _T_22_90 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h5b == io_wa) begin
        _T_22_91 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h5c == io_wa) begin
        _T_22_92 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h5d == io_wa) begin
        _T_22_93 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h5e == io_wa) begin
        _T_22_94 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h5f == io_wa) begin
        _T_22_95 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h60 == io_wa) begin
        _T_22_96 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h61 == io_wa) begin
        _T_22_97 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h62 == io_wa) begin
        _T_22_98 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h63 == io_wa) begin
        _T_22_99 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h64 == io_wa) begin
        _T_22_100 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h65 == io_wa) begin
        _T_22_101 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h66 == io_wa) begin
        _T_22_102 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h67 == io_wa) begin
        _T_22_103 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h68 == io_wa) begin
        _T_22_104 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h69 == io_wa) begin
        _T_22_105 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h6a == io_wa) begin
        _T_22_106 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h6b == io_wa) begin
        _T_22_107 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h6c == io_wa) begin
        _T_22_108 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h6d == io_wa) begin
        _T_22_109 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h6e == io_wa) begin
        _T_22_110 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h6f == io_wa) begin
        _T_22_111 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h70 == io_wa) begin
        _T_22_112 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h71 == io_wa) begin
        _T_22_113 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h72 == io_wa) begin
        _T_22_114 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h73 == io_wa) begin
        _T_22_115 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h74 == io_wa) begin
        _T_22_116 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h75 == io_wa) begin
        _T_22_117 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h76 == io_wa) begin
        _T_22_118 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h77 == io_wa) begin
        _T_22_119 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h78 == io_wa) begin
        _T_22_120 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h79 == io_wa) begin
        _T_22_121 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h7a == io_wa) begin
        _T_22_122 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h7b == io_wa) begin
        _T_22_123 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h7c == io_wa) begin
        _T_22_124 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h7d == io_wa) begin
        _T_22_125 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h7e == io_wa) begin
        _T_22_126 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h7f == io_wa) begin
        _T_22_127 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h80 == io_wa) begin
        _T_22_128 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h81 == io_wa) begin
        _T_22_129 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h82 == io_wa) begin
        _T_22_130 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h83 == io_wa) begin
        _T_22_131 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h84 == io_wa) begin
        _T_22_132 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h85 == io_wa) begin
        _T_22_133 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h86 == io_wa) begin
        _T_22_134 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h87 == io_wa) begin
        _T_22_135 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h88 == io_wa) begin
        _T_22_136 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h89 == io_wa) begin
        _T_22_137 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h8a == io_wa) begin
        _T_22_138 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h8b == io_wa) begin
        _T_22_139 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h8c == io_wa) begin
        _T_22_140 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h8d == io_wa) begin
        _T_22_141 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h8e == io_wa) begin
        _T_22_142 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h8f == io_wa) begin
        _T_22_143 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h90 == io_wa) begin
        _T_22_144 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h91 == io_wa) begin
        _T_22_145 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h92 == io_wa) begin
        _T_22_146 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h93 == io_wa) begin
        _T_22_147 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h94 == io_wa) begin
        _T_22_148 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h95 == io_wa) begin
        _T_22_149 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h96 == io_wa) begin
        _T_22_150 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h97 == io_wa) begin
        _T_22_151 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h98 == io_wa) begin
        _T_22_152 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h99 == io_wa) begin
        _T_22_153 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h9a == io_wa) begin
        _T_22_154 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h9b == io_wa) begin
        _T_22_155 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h9c == io_wa) begin
        _T_22_156 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h9d == io_wa) begin
        _T_22_157 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h9e == io_wa) begin
        _T_22_158 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h9f == io_wa) begin
        _T_22_159 <= io_di;
      end
    end
    if (io_we) begin
      if (9'ha0 == io_wa) begin
        _T_22_160 <= io_di;
      end
    end
    if (io_we) begin
      if (9'ha1 == io_wa) begin
        _T_22_161 <= io_di;
      end
    end
    if (io_we) begin
      if (9'ha2 == io_wa) begin
        _T_22_162 <= io_di;
      end
    end
    if (io_we) begin
      if (9'ha3 == io_wa) begin
        _T_22_163 <= io_di;
      end
    end
    if (io_we) begin
      if (9'ha4 == io_wa) begin
        _T_22_164 <= io_di;
      end
    end
    if (io_we) begin
      if (9'ha5 == io_wa) begin
        _T_22_165 <= io_di;
      end
    end
    if (io_we) begin
      if (9'ha6 == io_wa) begin
        _T_22_166 <= io_di;
      end
    end
    if (io_we) begin
      if (9'ha7 == io_wa) begin
        _T_22_167 <= io_di;
      end
    end
    if (io_we) begin
      if (9'ha8 == io_wa) begin
        _T_22_168 <= io_di;
      end
    end
    if (io_we) begin
      if (9'ha9 == io_wa) begin
        _T_22_169 <= io_di;
      end
    end
    if (io_we) begin
      if (9'haa == io_wa) begin
        _T_22_170 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hab == io_wa) begin
        _T_22_171 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hac == io_wa) begin
        _T_22_172 <= io_di;
      end
    end
    if (io_we) begin
      if (9'had == io_wa) begin
        _T_22_173 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hae == io_wa) begin
        _T_22_174 <= io_di;
      end
    end
    if (io_we) begin
      if (9'haf == io_wa) begin
        _T_22_175 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hb0 == io_wa) begin
        _T_22_176 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hb1 == io_wa) begin
        _T_22_177 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hb2 == io_wa) begin
        _T_22_178 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hb3 == io_wa) begin
        _T_22_179 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hb4 == io_wa) begin
        _T_22_180 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hb5 == io_wa) begin
        _T_22_181 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hb6 == io_wa) begin
        _T_22_182 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hb7 == io_wa) begin
        _T_22_183 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hb8 == io_wa) begin
        _T_22_184 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hb9 == io_wa) begin
        _T_22_185 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hba == io_wa) begin
        _T_22_186 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hbb == io_wa) begin
        _T_22_187 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hbc == io_wa) begin
        _T_22_188 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hbd == io_wa) begin
        _T_22_189 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hbe == io_wa) begin
        _T_22_190 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hbf == io_wa) begin
        _T_22_191 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hc0 == io_wa) begin
        _T_22_192 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hc1 == io_wa) begin
        _T_22_193 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hc2 == io_wa) begin
        _T_22_194 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hc3 == io_wa) begin
        _T_22_195 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hc4 == io_wa) begin
        _T_22_196 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hc5 == io_wa) begin
        _T_22_197 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hc6 == io_wa) begin
        _T_22_198 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hc7 == io_wa) begin
        _T_22_199 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hc8 == io_wa) begin
        _T_22_200 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hc9 == io_wa) begin
        _T_22_201 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hca == io_wa) begin
        _T_22_202 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hcb == io_wa) begin
        _T_22_203 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hcc == io_wa) begin
        _T_22_204 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hcd == io_wa) begin
        _T_22_205 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hce == io_wa) begin
        _T_22_206 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hcf == io_wa) begin
        _T_22_207 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hd0 == io_wa) begin
        _T_22_208 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hd1 == io_wa) begin
        _T_22_209 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hd2 == io_wa) begin
        _T_22_210 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hd3 == io_wa) begin
        _T_22_211 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hd4 == io_wa) begin
        _T_22_212 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hd5 == io_wa) begin
        _T_22_213 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hd6 == io_wa) begin
        _T_22_214 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hd7 == io_wa) begin
        _T_22_215 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hd8 == io_wa) begin
        _T_22_216 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hd9 == io_wa) begin
        _T_22_217 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hda == io_wa) begin
        _T_22_218 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hdb == io_wa) begin
        _T_22_219 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hdc == io_wa) begin
        _T_22_220 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hdd == io_wa) begin
        _T_22_221 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hde == io_wa) begin
        _T_22_222 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hdf == io_wa) begin
        _T_22_223 <= io_di;
      end
    end
    if (io_we) begin
      if (9'he0 == io_wa) begin
        _T_22_224 <= io_di;
      end
    end
    if (io_we) begin
      if (9'he1 == io_wa) begin
        _T_22_225 <= io_di;
      end
    end
    if (io_we) begin
      if (9'he2 == io_wa) begin
        _T_22_226 <= io_di;
      end
    end
    if (io_we) begin
      if (9'he3 == io_wa) begin
        _T_22_227 <= io_di;
      end
    end
    if (io_we) begin
      if (9'he4 == io_wa) begin
        _T_22_228 <= io_di;
      end
    end
    if (io_we) begin
      if (9'he5 == io_wa) begin
        _T_22_229 <= io_di;
      end
    end
    if (io_we) begin
      if (9'he6 == io_wa) begin
        _T_22_230 <= io_di;
      end
    end
    if (io_we) begin
      if (9'he7 == io_wa) begin
        _T_22_231 <= io_di;
      end
    end
    if (io_we) begin
      if (9'he8 == io_wa) begin
        _T_22_232 <= io_di;
      end
    end
    if (io_we) begin
      if (9'he9 == io_wa) begin
        _T_22_233 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hea == io_wa) begin
        _T_22_234 <= io_di;
      end
    end
    if (io_we) begin
      if (9'heb == io_wa) begin
        _T_22_235 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hec == io_wa) begin
        _T_22_236 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hed == io_wa) begin
        _T_22_237 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hee == io_wa) begin
        _T_22_238 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hef == io_wa) begin
        _T_22_239 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hf0 == io_wa) begin
        _T_22_240 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hf1 == io_wa) begin
        _T_22_241 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hf2 == io_wa) begin
        _T_22_242 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hf3 == io_wa) begin
        _T_22_243 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hf4 == io_wa) begin
        _T_22_244 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hf5 == io_wa) begin
        _T_22_245 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hf6 == io_wa) begin
        _T_22_246 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hf7 == io_wa) begin
        _T_22_247 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hf8 == io_wa) begin
        _T_22_248 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hf9 == io_wa) begin
        _T_22_249 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hfa == io_wa) begin
        _T_22_250 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hfb == io_wa) begin
        _T_22_251 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hfc == io_wa) begin
        _T_22_252 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hfd == io_wa) begin
        _T_22_253 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hfe == io_wa) begin
        _T_22_254 <= io_di;
      end
    end
    if (io_we) begin
      if (9'hff == io_wa) begin
        _T_22_255 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h100 == io_wa) begin
        _T_22_256 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h101 == io_wa) begin
        _T_22_257 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h102 == io_wa) begin
        _T_22_258 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h103 == io_wa) begin
        _T_22_259 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h104 == io_wa) begin
        _T_22_260 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h105 == io_wa) begin
        _T_22_261 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h106 == io_wa) begin
        _T_22_262 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h107 == io_wa) begin
        _T_22_263 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h108 == io_wa) begin
        _T_22_264 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h109 == io_wa) begin
        _T_22_265 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h10a == io_wa) begin
        _T_22_266 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h10b == io_wa) begin
        _T_22_267 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h10c == io_wa) begin
        _T_22_268 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h10d == io_wa) begin
        _T_22_269 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h10e == io_wa) begin
        _T_22_270 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h10f == io_wa) begin
        _T_22_271 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h110 == io_wa) begin
        _T_22_272 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h111 == io_wa) begin
        _T_22_273 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h112 == io_wa) begin
        _T_22_274 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h113 == io_wa) begin
        _T_22_275 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h114 == io_wa) begin
        _T_22_276 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h115 == io_wa) begin
        _T_22_277 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h116 == io_wa) begin
        _T_22_278 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h117 == io_wa) begin
        _T_22_279 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h118 == io_wa) begin
        _T_22_280 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h119 == io_wa) begin
        _T_22_281 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h11a == io_wa) begin
        _T_22_282 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h11b == io_wa) begin
        _T_22_283 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h11c == io_wa) begin
        _T_22_284 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h11d == io_wa) begin
        _T_22_285 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h11e == io_wa) begin
        _T_22_286 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h11f == io_wa) begin
        _T_22_287 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h120 == io_wa) begin
        _T_22_288 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h121 == io_wa) begin
        _T_22_289 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h122 == io_wa) begin
        _T_22_290 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h123 == io_wa) begin
        _T_22_291 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h124 == io_wa) begin
        _T_22_292 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h125 == io_wa) begin
        _T_22_293 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h126 == io_wa) begin
        _T_22_294 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h127 == io_wa) begin
        _T_22_295 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h128 == io_wa) begin
        _T_22_296 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h129 == io_wa) begin
        _T_22_297 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h12a == io_wa) begin
        _T_22_298 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h12b == io_wa) begin
        _T_22_299 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h12c == io_wa) begin
        _T_22_300 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h12d == io_wa) begin
        _T_22_301 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h12e == io_wa) begin
        _T_22_302 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h12f == io_wa) begin
        _T_22_303 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h130 == io_wa) begin
        _T_22_304 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h131 == io_wa) begin
        _T_22_305 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h132 == io_wa) begin
        _T_22_306 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h133 == io_wa) begin
        _T_22_307 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h134 == io_wa) begin
        _T_22_308 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h135 == io_wa) begin
        _T_22_309 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h136 == io_wa) begin
        _T_22_310 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h137 == io_wa) begin
        _T_22_311 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h138 == io_wa) begin
        _T_22_312 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h139 == io_wa) begin
        _T_22_313 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h13a == io_wa) begin
        _T_22_314 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h13b == io_wa) begin
        _T_22_315 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h13c == io_wa) begin
        _T_22_316 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h13d == io_wa) begin
        _T_22_317 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h13e == io_wa) begin
        _T_22_318 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h13f == io_wa) begin
        _T_22_319 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h140 == io_wa) begin
        _T_22_320 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h141 == io_wa) begin
        _T_22_321 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h142 == io_wa) begin
        _T_22_322 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h143 == io_wa) begin
        _T_22_323 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h144 == io_wa) begin
        _T_22_324 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h145 == io_wa) begin
        _T_22_325 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h146 == io_wa) begin
        _T_22_326 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h147 == io_wa) begin
        _T_22_327 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h148 == io_wa) begin
        _T_22_328 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h149 == io_wa) begin
        _T_22_329 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h14a == io_wa) begin
        _T_22_330 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h14b == io_wa) begin
        _T_22_331 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h14c == io_wa) begin
        _T_22_332 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h14d == io_wa) begin
        _T_22_333 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h14e == io_wa) begin
        _T_22_334 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h14f == io_wa) begin
        _T_22_335 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h150 == io_wa) begin
        _T_22_336 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h151 == io_wa) begin
        _T_22_337 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h152 == io_wa) begin
        _T_22_338 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h153 == io_wa) begin
        _T_22_339 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h154 == io_wa) begin
        _T_22_340 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h155 == io_wa) begin
        _T_22_341 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h156 == io_wa) begin
        _T_22_342 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h157 == io_wa) begin
        _T_22_343 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h158 == io_wa) begin
        _T_22_344 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h159 == io_wa) begin
        _T_22_345 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h15a == io_wa) begin
        _T_22_346 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h15b == io_wa) begin
        _T_22_347 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h15c == io_wa) begin
        _T_22_348 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h15d == io_wa) begin
        _T_22_349 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h15e == io_wa) begin
        _T_22_350 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h15f == io_wa) begin
        _T_22_351 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h160 == io_wa) begin
        _T_22_352 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h161 == io_wa) begin
        _T_22_353 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h162 == io_wa) begin
        _T_22_354 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h163 == io_wa) begin
        _T_22_355 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h164 == io_wa) begin
        _T_22_356 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h165 == io_wa) begin
        _T_22_357 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h166 == io_wa) begin
        _T_22_358 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h167 == io_wa) begin
        _T_22_359 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h168 == io_wa) begin
        _T_22_360 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h169 == io_wa) begin
        _T_22_361 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h16a == io_wa) begin
        _T_22_362 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h16b == io_wa) begin
        _T_22_363 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h16c == io_wa) begin
        _T_22_364 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h16d == io_wa) begin
        _T_22_365 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h16e == io_wa) begin
        _T_22_366 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h16f == io_wa) begin
        _T_22_367 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h170 == io_wa) begin
        _T_22_368 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h171 == io_wa) begin
        _T_22_369 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h172 == io_wa) begin
        _T_22_370 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h173 == io_wa) begin
        _T_22_371 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h174 == io_wa) begin
        _T_22_372 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h175 == io_wa) begin
        _T_22_373 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h176 == io_wa) begin
        _T_22_374 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h177 == io_wa) begin
        _T_22_375 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h178 == io_wa) begin
        _T_22_376 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h179 == io_wa) begin
        _T_22_377 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h17a == io_wa) begin
        _T_22_378 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h17b == io_wa) begin
        _T_22_379 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h17c == io_wa) begin
        _T_22_380 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h17d == io_wa) begin
        _T_22_381 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h17e == io_wa) begin
        _T_22_382 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h17f == io_wa) begin
        _T_22_383 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h180 == io_wa) begin
        _T_22_384 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h181 == io_wa) begin
        _T_22_385 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h182 == io_wa) begin
        _T_22_386 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h183 == io_wa) begin
        _T_22_387 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h184 == io_wa) begin
        _T_22_388 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h185 == io_wa) begin
        _T_22_389 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h186 == io_wa) begin
        _T_22_390 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h187 == io_wa) begin
        _T_22_391 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h188 == io_wa) begin
        _T_22_392 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h189 == io_wa) begin
        _T_22_393 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h18a == io_wa) begin
        _T_22_394 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h18b == io_wa) begin
        _T_22_395 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h18c == io_wa) begin
        _T_22_396 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h18d == io_wa) begin
        _T_22_397 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h18e == io_wa) begin
        _T_22_398 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h18f == io_wa) begin
        _T_22_399 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h190 == io_wa) begin
        _T_22_400 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h191 == io_wa) begin
        _T_22_401 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h192 == io_wa) begin
        _T_22_402 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h193 == io_wa) begin
        _T_22_403 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h194 == io_wa) begin
        _T_22_404 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h195 == io_wa) begin
        _T_22_405 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h196 == io_wa) begin
        _T_22_406 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h197 == io_wa) begin
        _T_22_407 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h198 == io_wa) begin
        _T_22_408 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h199 == io_wa) begin
        _T_22_409 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h19a == io_wa) begin
        _T_22_410 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h19b == io_wa) begin
        _T_22_411 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h19c == io_wa) begin
        _T_22_412 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h19d == io_wa) begin
        _T_22_413 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h19e == io_wa) begin
        _T_22_414 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h19f == io_wa) begin
        _T_22_415 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1a0 == io_wa) begin
        _T_22_416 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1a1 == io_wa) begin
        _T_22_417 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1a2 == io_wa) begin
        _T_22_418 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1a3 == io_wa) begin
        _T_22_419 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1a4 == io_wa) begin
        _T_22_420 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1a5 == io_wa) begin
        _T_22_421 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1a6 == io_wa) begin
        _T_22_422 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1a7 == io_wa) begin
        _T_22_423 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1a8 == io_wa) begin
        _T_22_424 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1a9 == io_wa) begin
        _T_22_425 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1aa == io_wa) begin
        _T_22_426 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1ab == io_wa) begin
        _T_22_427 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1ac == io_wa) begin
        _T_22_428 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1ad == io_wa) begin
        _T_22_429 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1ae == io_wa) begin
        _T_22_430 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1af == io_wa) begin
        _T_22_431 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1b0 == io_wa) begin
        _T_22_432 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1b1 == io_wa) begin
        _T_22_433 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1b2 == io_wa) begin
        _T_22_434 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1b3 == io_wa) begin
        _T_22_435 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1b4 == io_wa) begin
        _T_22_436 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1b5 == io_wa) begin
        _T_22_437 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1b6 == io_wa) begin
        _T_22_438 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1b7 == io_wa) begin
        _T_22_439 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1b8 == io_wa) begin
        _T_22_440 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1b9 == io_wa) begin
        _T_22_441 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1ba == io_wa) begin
        _T_22_442 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1bb == io_wa) begin
        _T_22_443 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1bc == io_wa) begin
        _T_22_444 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1bd == io_wa) begin
        _T_22_445 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1be == io_wa) begin
        _T_22_446 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1bf == io_wa) begin
        _T_22_447 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1c0 == io_wa) begin
        _T_22_448 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1c1 == io_wa) begin
        _T_22_449 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1c2 == io_wa) begin
        _T_22_450 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1c3 == io_wa) begin
        _T_22_451 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1c4 == io_wa) begin
        _T_22_452 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1c5 == io_wa) begin
        _T_22_453 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1c6 == io_wa) begin
        _T_22_454 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1c7 == io_wa) begin
        _T_22_455 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1c8 == io_wa) begin
        _T_22_456 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1c9 == io_wa) begin
        _T_22_457 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1ca == io_wa) begin
        _T_22_458 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1cb == io_wa) begin
        _T_22_459 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1cc == io_wa) begin
        _T_22_460 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1cd == io_wa) begin
        _T_22_461 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1ce == io_wa) begin
        _T_22_462 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1cf == io_wa) begin
        _T_22_463 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1d0 == io_wa) begin
        _T_22_464 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1d1 == io_wa) begin
        _T_22_465 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1d2 == io_wa) begin
        _T_22_466 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1d3 == io_wa) begin
        _T_22_467 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1d4 == io_wa) begin
        _T_22_468 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1d5 == io_wa) begin
        _T_22_469 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1d6 == io_wa) begin
        _T_22_470 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1d7 == io_wa) begin
        _T_22_471 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1d8 == io_wa) begin
        _T_22_472 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1d9 == io_wa) begin
        _T_22_473 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1da == io_wa) begin
        _T_22_474 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1db == io_wa) begin
        _T_22_475 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1dc == io_wa) begin
        _T_22_476 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1dd == io_wa) begin
        _T_22_477 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1de == io_wa) begin
        _T_22_478 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1df == io_wa) begin
        _T_22_479 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1e0 == io_wa) begin
        _T_22_480 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1e1 == io_wa) begin
        _T_22_481 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1e2 == io_wa) begin
        _T_22_482 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1e3 == io_wa) begin
        _T_22_483 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1e4 == io_wa) begin
        _T_22_484 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1e5 == io_wa) begin
        _T_22_485 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1e6 == io_wa) begin
        _T_22_486 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1e7 == io_wa) begin
        _T_22_487 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1e8 == io_wa) begin
        _T_22_488 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1e9 == io_wa) begin
        _T_22_489 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1ea == io_wa) begin
        _T_22_490 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1eb == io_wa) begin
        _T_22_491 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1ec == io_wa) begin
        _T_22_492 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1ed == io_wa) begin
        _T_22_493 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1ee == io_wa) begin
        _T_22_494 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1ef == io_wa) begin
        _T_22_495 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1f0 == io_wa) begin
        _T_22_496 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1f1 == io_wa) begin
        _T_22_497 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1f2 == io_wa) begin
        _T_22_498 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1f3 == io_wa) begin
        _T_22_499 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1f4 == io_wa) begin
        _T_22_500 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1f5 == io_wa) begin
        _T_22_501 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1f6 == io_wa) begin
        _T_22_502 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1f7 == io_wa) begin
        _T_22_503 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1f8 == io_wa) begin
        _T_22_504 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1f9 == io_wa) begin
        _T_22_505 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1fa == io_wa) begin
        _T_22_506 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1fb == io_wa) begin
        _T_22_507 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1fc == io_wa) begin
        _T_22_508 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1fd == io_wa) begin
        _T_22_509 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1fe == io_wa) begin
        _T_22_510 <= io_di;
      end
    end
    if (io_we) begin
      if (9'h1ff == io_wa) begin
        _T_22_511 <= io_di;
      end
    end
    if (io_re) begin
      _T_538 <= io_ra;
    end
  end
endmodule
module NV_soDLA_cbuf( // @[:@483.2]
  input          clock, // @[:@484.4]
  input          reset, // @[:@485.4]
  input          io_nvdla_core_clk, // @[:@486.4]
  input          io_nvdla_core_rstn, // @[:@486.4]
  input  [31:0]  io_pwrbus_ram_pd, // @[:@486.4]
  input          io_cdma2buf_wr_en_0, // @[:@486.4]
  input          io_cdma2buf_wr_en_1, // @[:@486.4]
  input  [1:0]   io_cdma2buf_wr_sel_0, // @[:@486.4]
  input  [1:0]   io_cdma2buf_wr_sel_1, // @[:@486.4]
  input  [12:0]  io_cdma2buf_wr_addr_0, // @[:@486.4]
  input  [12:0]  io_cdma2buf_wr_addr_1, // @[:@486.4]
  input  [255:0] io_cdma2buf_wr_data_0, // @[:@486.4]
  input  [255:0] io_cdma2buf_wr_data_1, // @[:@486.4]
  input          io_sc2buf_dat_rd_addr_valid, // @[:@486.4]
  input  [12:0]  io_sc2buf_dat_rd_addr_bits, // @[:@486.4]
  output         io_sc2buf_dat_rd_data_valid, // @[:@486.4]
  output [511:0] io_sc2buf_dat_rd_data_bits, // @[:@486.4]
  input          io_sc2buf_wt_rd_addr_valid, // @[:@486.4]
  input  [12:0]  io_sc2buf_wt_rd_addr_bits, // @[:@486.4]
  output         io_sc2buf_wt_rd_data_valid, // @[:@486.4]
  output [511:0] io_sc2buf_wt_rd_data_bits // @[:@486.4]
);
  wire  nv_ram_rws_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3837.4]
  wire  nv_ram_rws_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3837.4]
  wire  nv_ram_rws_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3837.4]
  wire [8:0] nv_ram_rws_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3837.4]
  wire [8:0] nv_ram_rws_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3837.4]
  wire [255:0] nv_ram_rws_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3837.4]
  wire [255:0] nv_ram_rws_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3837.4]
  wire  nv_ram_rws_1_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3840.4]
  wire  nv_ram_rws_1_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3840.4]
  wire  nv_ram_rws_1_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3840.4]
  wire [8:0] nv_ram_rws_1_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3840.4]
  wire [8:0] nv_ram_rws_1_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3840.4]
  wire [255:0] nv_ram_rws_1_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3840.4]
  wire [255:0] nv_ram_rws_1_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3840.4]
  wire  nv_ram_rws_2_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3843.4]
  wire  nv_ram_rws_2_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3843.4]
  wire  nv_ram_rws_2_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3843.4]
  wire [8:0] nv_ram_rws_2_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3843.4]
  wire [8:0] nv_ram_rws_2_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3843.4]
  wire [255:0] nv_ram_rws_2_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3843.4]
  wire [255:0] nv_ram_rws_2_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3843.4]
  wire  nv_ram_rws_3_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3846.4]
  wire  nv_ram_rws_3_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3846.4]
  wire  nv_ram_rws_3_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3846.4]
  wire [8:0] nv_ram_rws_3_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3846.4]
  wire [8:0] nv_ram_rws_3_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3846.4]
  wire [255:0] nv_ram_rws_3_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3846.4]
  wire [255:0] nv_ram_rws_3_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3846.4]
  wire  nv_ram_rws_4_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3849.4]
  wire  nv_ram_rws_4_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3849.4]
  wire  nv_ram_rws_4_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3849.4]
  wire [8:0] nv_ram_rws_4_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3849.4]
  wire [8:0] nv_ram_rws_4_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3849.4]
  wire [255:0] nv_ram_rws_4_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3849.4]
  wire [255:0] nv_ram_rws_4_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3849.4]
  wire  nv_ram_rws_5_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3852.4]
  wire  nv_ram_rws_5_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3852.4]
  wire  nv_ram_rws_5_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3852.4]
  wire [8:0] nv_ram_rws_5_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3852.4]
  wire [8:0] nv_ram_rws_5_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3852.4]
  wire [255:0] nv_ram_rws_5_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3852.4]
  wire [255:0] nv_ram_rws_5_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3852.4]
  wire  nv_ram_rws_6_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3855.4]
  wire  nv_ram_rws_6_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3855.4]
  wire  nv_ram_rws_6_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3855.4]
  wire [8:0] nv_ram_rws_6_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3855.4]
  wire [8:0] nv_ram_rws_6_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3855.4]
  wire [255:0] nv_ram_rws_6_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3855.4]
  wire [255:0] nv_ram_rws_6_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3855.4]
  wire  nv_ram_rws_7_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3858.4]
  wire  nv_ram_rws_7_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3858.4]
  wire  nv_ram_rws_7_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3858.4]
  wire [8:0] nv_ram_rws_7_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3858.4]
  wire [8:0] nv_ram_rws_7_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3858.4]
  wire [255:0] nv_ram_rws_7_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3858.4]
  wire [255:0] nv_ram_rws_7_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3858.4]
  wire  nv_ram_rws_8_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3861.4]
  wire  nv_ram_rws_8_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3861.4]
  wire  nv_ram_rws_8_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3861.4]
  wire [8:0] nv_ram_rws_8_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3861.4]
  wire [8:0] nv_ram_rws_8_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3861.4]
  wire [255:0] nv_ram_rws_8_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3861.4]
  wire [255:0] nv_ram_rws_8_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3861.4]
  wire  nv_ram_rws_9_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3864.4]
  wire  nv_ram_rws_9_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3864.4]
  wire  nv_ram_rws_9_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3864.4]
  wire [8:0] nv_ram_rws_9_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3864.4]
  wire [8:0] nv_ram_rws_9_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3864.4]
  wire [255:0] nv_ram_rws_9_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3864.4]
  wire [255:0] nv_ram_rws_9_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3864.4]
  wire  nv_ram_rws_10_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3867.4]
  wire  nv_ram_rws_10_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3867.4]
  wire  nv_ram_rws_10_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3867.4]
  wire [8:0] nv_ram_rws_10_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3867.4]
  wire [8:0] nv_ram_rws_10_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3867.4]
  wire [255:0] nv_ram_rws_10_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3867.4]
  wire [255:0] nv_ram_rws_10_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3867.4]
  wire  nv_ram_rws_11_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3870.4]
  wire  nv_ram_rws_11_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3870.4]
  wire  nv_ram_rws_11_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3870.4]
  wire [8:0] nv_ram_rws_11_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3870.4]
  wire [8:0] nv_ram_rws_11_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3870.4]
  wire [255:0] nv_ram_rws_11_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3870.4]
  wire [255:0] nv_ram_rws_11_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3870.4]
  wire  nv_ram_rws_12_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3873.4]
  wire  nv_ram_rws_12_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3873.4]
  wire  nv_ram_rws_12_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3873.4]
  wire [8:0] nv_ram_rws_12_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3873.4]
  wire [8:0] nv_ram_rws_12_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3873.4]
  wire [255:0] nv_ram_rws_12_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3873.4]
  wire [255:0] nv_ram_rws_12_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3873.4]
  wire  nv_ram_rws_13_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3876.4]
  wire  nv_ram_rws_13_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3876.4]
  wire  nv_ram_rws_13_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3876.4]
  wire [8:0] nv_ram_rws_13_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3876.4]
  wire [8:0] nv_ram_rws_13_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3876.4]
  wire [255:0] nv_ram_rws_13_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3876.4]
  wire [255:0] nv_ram_rws_13_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3876.4]
  wire  nv_ram_rws_14_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3879.4]
  wire  nv_ram_rws_14_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3879.4]
  wire  nv_ram_rws_14_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3879.4]
  wire [8:0] nv_ram_rws_14_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3879.4]
  wire [8:0] nv_ram_rws_14_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3879.4]
  wire [255:0] nv_ram_rws_14_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3879.4]
  wire [255:0] nv_ram_rws_14_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3879.4]
  wire  nv_ram_rws_15_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3882.4]
  wire  nv_ram_rws_15_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3882.4]
  wire  nv_ram_rws_15_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3882.4]
  wire [8:0] nv_ram_rws_15_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3882.4]
  wire [8:0] nv_ram_rws_15_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3882.4]
  wire [255:0] nv_ram_rws_15_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3882.4]
  wire [255:0] nv_ram_rws_15_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3882.4]
  wire  nv_ram_rws_16_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3885.4]
  wire  nv_ram_rws_16_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3885.4]
  wire  nv_ram_rws_16_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3885.4]
  wire [8:0] nv_ram_rws_16_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3885.4]
  wire [8:0] nv_ram_rws_16_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3885.4]
  wire [255:0] nv_ram_rws_16_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3885.4]
  wire [255:0] nv_ram_rws_16_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3885.4]
  wire  nv_ram_rws_17_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3888.4]
  wire  nv_ram_rws_17_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3888.4]
  wire  nv_ram_rws_17_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3888.4]
  wire [8:0] nv_ram_rws_17_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3888.4]
  wire [8:0] nv_ram_rws_17_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3888.4]
  wire [255:0] nv_ram_rws_17_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3888.4]
  wire [255:0] nv_ram_rws_17_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3888.4]
  wire  nv_ram_rws_18_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3891.4]
  wire  nv_ram_rws_18_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3891.4]
  wire  nv_ram_rws_18_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3891.4]
  wire [8:0] nv_ram_rws_18_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3891.4]
  wire [8:0] nv_ram_rws_18_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3891.4]
  wire [255:0] nv_ram_rws_18_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3891.4]
  wire [255:0] nv_ram_rws_18_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3891.4]
  wire  nv_ram_rws_19_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3894.4]
  wire  nv_ram_rws_19_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3894.4]
  wire  nv_ram_rws_19_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3894.4]
  wire [8:0] nv_ram_rws_19_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3894.4]
  wire [8:0] nv_ram_rws_19_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3894.4]
  wire [255:0] nv_ram_rws_19_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3894.4]
  wire [255:0] nv_ram_rws_19_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3894.4]
  wire  nv_ram_rws_20_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3897.4]
  wire  nv_ram_rws_20_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3897.4]
  wire  nv_ram_rws_20_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3897.4]
  wire [8:0] nv_ram_rws_20_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3897.4]
  wire [8:0] nv_ram_rws_20_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3897.4]
  wire [255:0] nv_ram_rws_20_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3897.4]
  wire [255:0] nv_ram_rws_20_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3897.4]
  wire  nv_ram_rws_21_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3900.4]
  wire  nv_ram_rws_21_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3900.4]
  wire  nv_ram_rws_21_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3900.4]
  wire [8:0] nv_ram_rws_21_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3900.4]
  wire [8:0] nv_ram_rws_21_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3900.4]
  wire [255:0] nv_ram_rws_21_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3900.4]
  wire [255:0] nv_ram_rws_21_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3900.4]
  wire  nv_ram_rws_22_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3903.4]
  wire  nv_ram_rws_22_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3903.4]
  wire  nv_ram_rws_22_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3903.4]
  wire [8:0] nv_ram_rws_22_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3903.4]
  wire [8:0] nv_ram_rws_22_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3903.4]
  wire [255:0] nv_ram_rws_22_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3903.4]
  wire [255:0] nv_ram_rws_22_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3903.4]
  wire  nv_ram_rws_23_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3906.4]
  wire  nv_ram_rws_23_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3906.4]
  wire  nv_ram_rws_23_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3906.4]
  wire [8:0] nv_ram_rws_23_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3906.4]
  wire [8:0] nv_ram_rws_23_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3906.4]
  wire [255:0] nv_ram_rws_23_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3906.4]
  wire [255:0] nv_ram_rws_23_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3906.4]
  wire  nv_ram_rws_24_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3909.4]
  wire  nv_ram_rws_24_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3909.4]
  wire  nv_ram_rws_24_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3909.4]
  wire [8:0] nv_ram_rws_24_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3909.4]
  wire [8:0] nv_ram_rws_24_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3909.4]
  wire [255:0] nv_ram_rws_24_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3909.4]
  wire [255:0] nv_ram_rws_24_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3909.4]
  wire  nv_ram_rws_25_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3912.4]
  wire  nv_ram_rws_25_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3912.4]
  wire  nv_ram_rws_25_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3912.4]
  wire [8:0] nv_ram_rws_25_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3912.4]
  wire [8:0] nv_ram_rws_25_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3912.4]
  wire [255:0] nv_ram_rws_25_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3912.4]
  wire [255:0] nv_ram_rws_25_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3912.4]
  wire  nv_ram_rws_26_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3915.4]
  wire  nv_ram_rws_26_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3915.4]
  wire  nv_ram_rws_26_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3915.4]
  wire [8:0] nv_ram_rws_26_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3915.4]
  wire [8:0] nv_ram_rws_26_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3915.4]
  wire [255:0] nv_ram_rws_26_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3915.4]
  wire [255:0] nv_ram_rws_26_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3915.4]
  wire  nv_ram_rws_27_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3918.4]
  wire  nv_ram_rws_27_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3918.4]
  wire  nv_ram_rws_27_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3918.4]
  wire [8:0] nv_ram_rws_27_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3918.4]
  wire [8:0] nv_ram_rws_27_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3918.4]
  wire [255:0] nv_ram_rws_27_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3918.4]
  wire [255:0] nv_ram_rws_27_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3918.4]
  wire  nv_ram_rws_28_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3921.4]
  wire  nv_ram_rws_28_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3921.4]
  wire  nv_ram_rws_28_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3921.4]
  wire [8:0] nv_ram_rws_28_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3921.4]
  wire [8:0] nv_ram_rws_28_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3921.4]
  wire [255:0] nv_ram_rws_28_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3921.4]
  wire [255:0] nv_ram_rws_28_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3921.4]
  wire  nv_ram_rws_29_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3924.4]
  wire  nv_ram_rws_29_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3924.4]
  wire  nv_ram_rws_29_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3924.4]
  wire [8:0] nv_ram_rws_29_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3924.4]
  wire [8:0] nv_ram_rws_29_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3924.4]
  wire [255:0] nv_ram_rws_29_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3924.4]
  wire [255:0] nv_ram_rws_29_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3924.4]
  wire  nv_ram_rws_30_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3927.4]
  wire  nv_ram_rws_30_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3927.4]
  wire  nv_ram_rws_30_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3927.4]
  wire [8:0] nv_ram_rws_30_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3927.4]
  wire [8:0] nv_ram_rws_30_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3927.4]
  wire [255:0] nv_ram_rws_30_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3927.4]
  wire [255:0] nv_ram_rws_30_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3927.4]
  wire  nv_ram_rws_31_io_clk; // @[NV_NVDLA_cbuf.scala 389:106:@3930.4]
  wire  nv_ram_rws_31_io_re; // @[NV_NVDLA_cbuf.scala 389:106:@3930.4]
  wire  nv_ram_rws_31_io_we; // @[NV_NVDLA_cbuf.scala 389:106:@3930.4]
  wire [8:0] nv_ram_rws_31_io_ra; // @[NV_NVDLA_cbuf.scala 389:106:@3930.4]
  wire [8:0] nv_ram_rws_31_io_wa; // @[NV_NVDLA_cbuf.scala 389:106:@3930.4]
  wire [255:0] nv_ram_rws_31_io_di; // @[NV_NVDLA_cbuf.scala 389:106:@3930.4]
  wire [255:0] nv_ram_rws_31_io_dout; // @[NV_NVDLA_cbuf.scala 389:106:@3930.4]
  wire  _T_178; // @[NV_NVDLA_cbuf.scala 26:38:@488.4]
  wire [3:0] _T_2665; // @[NV_NVDLA_cbuf.scala 35:72:@490.4]
  wire  _T_2667; // @[NV_NVDLA_cbuf.scala 35:123:@491.4]
  wire  _T_2668; // @[NV_NVDLA_cbuf.scala 34:69:@492.4]
  wire  _T_2669; // @[NV_NVDLA_cbuf.scala 36:71:@493.4]
  wire  _T_2672; // @[NV_NVDLA_cbuf.scala 35:130:@495.4]
  wire [3:0] _T_2673; // @[NV_NVDLA_cbuf.scala 35:72:@497.4]
  wire  _T_2675; // @[NV_NVDLA_cbuf.scala 35:123:@498.4]
  wire  _T_2676; // @[NV_NVDLA_cbuf.scala 34:69:@499.4]
  wire  _T_2677; // @[NV_NVDLA_cbuf.scala 36:71:@500.4]
  wire  _T_2680; // @[NV_NVDLA_cbuf.scala 35:130:@502.4]
  wire  _T_2685; // @[NV_NVDLA_cbuf.scala 36:71:@507.4]
  wire  _T_2688; // @[NV_NVDLA_cbuf.scala 35:130:@509.4]
  wire  _T_2693; // @[NV_NVDLA_cbuf.scala 36:71:@514.4]
  wire  _T_2696; // @[NV_NVDLA_cbuf.scala 35:130:@516.4]
  wire  _T_2699; // @[NV_NVDLA_cbuf.scala 35:123:@519.4]
  wire  _T_2700; // @[NV_NVDLA_cbuf.scala 34:69:@520.4]
  wire  _T_2704; // @[NV_NVDLA_cbuf.scala 35:130:@523.4]
  wire  _T_2707; // @[NV_NVDLA_cbuf.scala 35:123:@526.4]
  wire  _T_2708; // @[NV_NVDLA_cbuf.scala 34:69:@527.4]
  wire  _T_2712; // @[NV_NVDLA_cbuf.scala 35:130:@530.4]
  wire  _T_2720; // @[NV_NVDLA_cbuf.scala 35:130:@537.4]
  wire  _T_2728; // @[NV_NVDLA_cbuf.scala 35:130:@544.4]
  wire  _T_2731; // @[NV_NVDLA_cbuf.scala 35:123:@547.4]
  wire  _T_2732; // @[NV_NVDLA_cbuf.scala 34:69:@548.4]
  wire  _T_2736; // @[NV_NVDLA_cbuf.scala 35:130:@551.4]
  wire  _T_2739; // @[NV_NVDLA_cbuf.scala 35:123:@554.4]
  wire  _T_2740; // @[NV_NVDLA_cbuf.scala 34:69:@555.4]
  wire  _T_2744; // @[NV_NVDLA_cbuf.scala 35:130:@558.4]
  wire  _T_2752; // @[NV_NVDLA_cbuf.scala 35:130:@565.4]
  wire  _T_2760; // @[NV_NVDLA_cbuf.scala 35:130:@572.4]
  wire  _T_2763; // @[NV_NVDLA_cbuf.scala 35:123:@575.4]
  wire  _T_2764; // @[NV_NVDLA_cbuf.scala 34:69:@576.4]
  wire  _T_2768; // @[NV_NVDLA_cbuf.scala 35:130:@579.4]
  wire  _T_2771; // @[NV_NVDLA_cbuf.scala 35:123:@582.4]
  wire  _T_2772; // @[NV_NVDLA_cbuf.scala 34:69:@583.4]
  wire  _T_2776; // @[NV_NVDLA_cbuf.scala 35:130:@586.4]
  wire  _T_2784; // @[NV_NVDLA_cbuf.scala 35:130:@593.4]
  wire  _T_2792; // @[NV_NVDLA_cbuf.scala 35:130:@600.4]
  wire  _T_2795; // @[NV_NVDLA_cbuf.scala 35:123:@603.4]
  wire  _T_2796; // @[NV_NVDLA_cbuf.scala 34:69:@604.4]
  wire  _T_2800; // @[NV_NVDLA_cbuf.scala 35:130:@607.4]
  wire  _T_2803; // @[NV_NVDLA_cbuf.scala 35:123:@610.4]
  wire  _T_2804; // @[NV_NVDLA_cbuf.scala 34:69:@611.4]
  wire  _T_2808; // @[NV_NVDLA_cbuf.scala 35:130:@614.4]
  wire  _T_2816; // @[NV_NVDLA_cbuf.scala 35:130:@621.4]
  wire  _T_2824; // @[NV_NVDLA_cbuf.scala 35:130:@628.4]
  wire  _T_2827; // @[NV_NVDLA_cbuf.scala 35:123:@631.4]
  wire  _T_2828; // @[NV_NVDLA_cbuf.scala 34:69:@632.4]
  wire  _T_2832; // @[NV_NVDLA_cbuf.scala 35:130:@635.4]
  wire  _T_2835; // @[NV_NVDLA_cbuf.scala 35:123:@638.4]
  wire  _T_2836; // @[NV_NVDLA_cbuf.scala 34:69:@639.4]
  wire  _T_2840; // @[NV_NVDLA_cbuf.scala 35:130:@642.4]
  wire  _T_2848; // @[NV_NVDLA_cbuf.scala 35:130:@649.4]
  wire  _T_2856; // @[NV_NVDLA_cbuf.scala 35:130:@656.4]
  wire  _T_2859; // @[NV_NVDLA_cbuf.scala 35:123:@659.4]
  wire  _T_2860; // @[NV_NVDLA_cbuf.scala 34:69:@660.4]
  wire  _T_2864; // @[NV_NVDLA_cbuf.scala 35:130:@663.4]
  wire  _T_2867; // @[NV_NVDLA_cbuf.scala 35:123:@666.4]
  wire  _T_2868; // @[NV_NVDLA_cbuf.scala 34:69:@667.4]
  wire  _T_2872; // @[NV_NVDLA_cbuf.scala 35:130:@670.4]
  wire  _T_2880; // @[NV_NVDLA_cbuf.scala 35:130:@677.4]
  wire  _T_2888; // @[NV_NVDLA_cbuf.scala 35:130:@684.4]
  wire  _T_2891; // @[NV_NVDLA_cbuf.scala 35:123:@687.4]
  wire  _T_2892; // @[NV_NVDLA_cbuf.scala 34:69:@688.4]
  wire  _T_2896; // @[NV_NVDLA_cbuf.scala 35:130:@691.4]
  wire  _T_2899; // @[NV_NVDLA_cbuf.scala 35:123:@694.4]
  wire  _T_2900; // @[NV_NVDLA_cbuf.scala 34:69:@695.4]
  wire  _T_2904; // @[NV_NVDLA_cbuf.scala 35:130:@698.4]
  wire  _T_2912; // @[NV_NVDLA_cbuf.scala 35:130:@705.4]
  wire  _T_2920; // @[NV_NVDLA_cbuf.scala 35:130:@712.4]
  wire  _T_2923; // @[NV_NVDLA_cbuf.scala 35:123:@715.4]
  wire  _T_2924; // @[NV_NVDLA_cbuf.scala 34:69:@716.4]
  wire  _T_2928; // @[NV_NVDLA_cbuf.scala 35:130:@719.4]
  wire  _T_2931; // @[NV_NVDLA_cbuf.scala 35:123:@722.4]
  wire  _T_2932; // @[NV_NVDLA_cbuf.scala 34:69:@723.4]
  wire  _T_2936; // @[NV_NVDLA_cbuf.scala 35:130:@726.4]
  wire  _T_2944; // @[NV_NVDLA_cbuf.scala 35:130:@733.4]
  wire  _T_2952; // @[NV_NVDLA_cbuf.scala 35:130:@740.4]
  wire  _T_2955; // @[NV_NVDLA_cbuf.scala 35:123:@743.4]
  wire  _T_2956; // @[NV_NVDLA_cbuf.scala 34:69:@744.4]
  wire  _T_2960; // @[NV_NVDLA_cbuf.scala 35:130:@747.4]
  wire  _T_2963; // @[NV_NVDLA_cbuf.scala 35:123:@750.4]
  wire  _T_2964; // @[NV_NVDLA_cbuf.scala 34:69:@751.4]
  wire  _T_2968; // @[NV_NVDLA_cbuf.scala 35:130:@754.4]
  wire  _T_2976; // @[NV_NVDLA_cbuf.scala 35:130:@761.4]
  wire  _T_2984; // @[NV_NVDLA_cbuf.scala 35:130:@768.4]
  wire  _T_2987; // @[NV_NVDLA_cbuf.scala 35:123:@771.4]
  wire  _T_2988; // @[NV_NVDLA_cbuf.scala 34:69:@772.4]
  wire  _T_2992; // @[NV_NVDLA_cbuf.scala 35:130:@775.4]
  wire  _T_2995; // @[NV_NVDLA_cbuf.scala 35:123:@778.4]
  wire  _T_2996; // @[NV_NVDLA_cbuf.scala 34:69:@779.4]
  wire  _T_3000; // @[NV_NVDLA_cbuf.scala 35:130:@782.4]
  wire  _T_3008; // @[NV_NVDLA_cbuf.scala 35:130:@789.4]
  wire  _T_3016; // @[NV_NVDLA_cbuf.scala 35:130:@796.4]
  wire  _T_3019; // @[NV_NVDLA_cbuf.scala 35:123:@799.4]
  wire  _T_3020; // @[NV_NVDLA_cbuf.scala 34:69:@800.4]
  wire  _T_3024; // @[NV_NVDLA_cbuf.scala 35:130:@803.4]
  wire  _T_3027; // @[NV_NVDLA_cbuf.scala 35:123:@806.4]
  wire  _T_3028; // @[NV_NVDLA_cbuf.scala 34:69:@807.4]
  wire  _T_3032; // @[NV_NVDLA_cbuf.scala 35:130:@810.4]
  wire  _T_3040; // @[NV_NVDLA_cbuf.scala 35:130:@817.4]
  wire  _T_3048; // @[NV_NVDLA_cbuf.scala 35:130:@824.4]
  wire  _T_3051; // @[NV_NVDLA_cbuf.scala 35:123:@827.4]
  wire  _T_3052; // @[NV_NVDLA_cbuf.scala 34:69:@828.4]
  wire  _T_3056; // @[NV_NVDLA_cbuf.scala 35:130:@831.4]
  wire  _T_3059; // @[NV_NVDLA_cbuf.scala 35:123:@834.4]
  wire  _T_3060; // @[NV_NVDLA_cbuf.scala 34:69:@835.4]
  wire  _T_3064; // @[NV_NVDLA_cbuf.scala 35:130:@838.4]
  wire  _T_3072; // @[NV_NVDLA_cbuf.scala 35:130:@845.4]
  wire  _T_3080; // @[NV_NVDLA_cbuf.scala 35:130:@852.4]
  wire  _T_3083; // @[NV_NVDLA_cbuf.scala 35:123:@855.4]
  wire  _T_3084; // @[NV_NVDLA_cbuf.scala 34:69:@856.4]
  wire  _T_3088; // @[NV_NVDLA_cbuf.scala 35:130:@859.4]
  wire  _T_3091; // @[NV_NVDLA_cbuf.scala 35:123:@862.4]
  wire  _T_3092; // @[NV_NVDLA_cbuf.scala 34:69:@863.4]
  wire  _T_3096; // @[NV_NVDLA_cbuf.scala 35:130:@866.4]
  wire  _T_3104; // @[NV_NVDLA_cbuf.scala 35:130:@873.4]
  wire  _T_3112; // @[NV_NVDLA_cbuf.scala 35:130:@880.4]
  wire  _T_3115; // @[NV_NVDLA_cbuf.scala 35:123:@883.4]
  wire  _T_3116; // @[NV_NVDLA_cbuf.scala 34:69:@884.4]
  wire  _T_3120; // @[NV_NVDLA_cbuf.scala 35:130:@887.4]
  wire  _T_3123; // @[NV_NVDLA_cbuf.scala 35:123:@890.4]
  wire  _T_3124; // @[NV_NVDLA_cbuf.scala 34:69:@891.4]
  wire  _T_3128; // @[NV_NVDLA_cbuf.scala 35:130:@894.4]
  wire  _T_3136; // @[NV_NVDLA_cbuf.scala 35:130:@901.4]
  wire  _T_3144; // @[NV_NVDLA_cbuf.scala 35:130:@908.4]
  wire  _T_3147; // @[NV_NVDLA_cbuf.scala 35:123:@911.4]
  wire  _T_3148; // @[NV_NVDLA_cbuf.scala 34:69:@912.4]
  wire  _T_3152; // @[NV_NVDLA_cbuf.scala 35:130:@915.4]
  wire  _T_3155; // @[NV_NVDLA_cbuf.scala 35:123:@918.4]
  wire  _T_3156; // @[NV_NVDLA_cbuf.scala 34:69:@919.4]
  wire  _T_3160; // @[NV_NVDLA_cbuf.scala 35:130:@922.4]
  wire  _T_3168; // @[NV_NVDLA_cbuf.scala 35:130:@929.4]
  wire  _T_3176; // @[NV_NVDLA_cbuf.scala 35:130:@936.4]
  reg  _T_7112_0_0; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_0;
  reg  _T_7112_0_1; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_1;
  reg  _T_7112_1_0; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_2;
  reg  _T_7112_1_1; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_3;
  reg  _T_7112_2_0; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_4;
  reg  _T_7112_2_1; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_5;
  reg  _T_7112_3_0; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_6;
  reg  _T_7112_3_1; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_7;
  reg  _T_7112_4_0; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_8;
  reg  _T_7112_4_1; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_9;
  reg  _T_7112_5_0; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_10;
  reg  _T_7112_5_1; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_11;
  reg  _T_7112_6_0; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_12;
  reg  _T_7112_6_1; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_13;
  reg  _T_7112_7_0; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_14;
  reg  _T_7112_7_1; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_15;
  reg  _T_7112_8_0; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_16;
  reg  _T_7112_8_1; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_17;
  reg  _T_7112_9_0; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_18;
  reg  _T_7112_9_1; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_19;
  reg  _T_7112_10_0; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_20;
  reg  _T_7112_10_1; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_21;
  reg  _T_7112_11_0; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_22;
  reg  _T_7112_11_1; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_23;
  reg  _T_7112_12_0; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_24;
  reg  _T_7112_12_1; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_25;
  reg  _T_7112_13_0; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_26;
  reg  _T_7112_13_1; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_27;
  reg  _T_7112_14_0; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_28;
  reg  _T_7112_14_1; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_29;
  reg  _T_7112_15_0; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_30;
  reg  _T_7112_15_1; // @[NV_NVDLA_cbuf.scala 71:36:@1084.4]
  reg [31:0] _RAND_31;
  wire  _T_8151; // @[NV_NVDLA_cbuf.scala 74:72:@1085.4]
  wire  _T_8152; // @[NV_NVDLA_cbuf.scala 74:72:@1087.4]
  wire  _T_8153; // @[NV_NVDLA_cbuf.scala 74:72:@1089.4]
  wire  _T_8154; // @[NV_NVDLA_cbuf.scala 74:72:@1091.4]
  wire  _T_8155; // @[NV_NVDLA_cbuf.scala 74:72:@1093.4]
  wire  _T_8156; // @[NV_NVDLA_cbuf.scala 74:72:@1095.4]
  wire  _T_8157; // @[NV_NVDLA_cbuf.scala 74:72:@1097.4]
  wire  _T_8158; // @[NV_NVDLA_cbuf.scala 74:72:@1099.4]
  wire  _T_8159; // @[NV_NVDLA_cbuf.scala 74:72:@1101.4]
  wire  _T_8160; // @[NV_NVDLA_cbuf.scala 74:72:@1103.4]
  wire  _T_8161; // @[NV_NVDLA_cbuf.scala 74:72:@1105.4]
  wire  _T_8162; // @[NV_NVDLA_cbuf.scala 74:72:@1107.4]
  wire  _T_8163; // @[NV_NVDLA_cbuf.scala 74:72:@1109.4]
  wire  _T_8164; // @[NV_NVDLA_cbuf.scala 74:72:@1111.4]
  wire  _T_8165; // @[NV_NVDLA_cbuf.scala 74:72:@1113.4]
  wire  _T_8166; // @[NV_NVDLA_cbuf.scala 74:72:@1115.4]
  wire  _T_8167; // @[NV_NVDLA_cbuf.scala 74:72:@1117.4]
  wire  _T_8168; // @[NV_NVDLA_cbuf.scala 74:72:@1119.4]
  wire  _T_8169; // @[NV_NVDLA_cbuf.scala 74:72:@1121.4]
  wire  _T_8170; // @[NV_NVDLA_cbuf.scala 74:72:@1123.4]
  wire  _T_8171; // @[NV_NVDLA_cbuf.scala 74:72:@1125.4]
  wire  _T_8172; // @[NV_NVDLA_cbuf.scala 74:72:@1127.4]
  wire  _T_8173; // @[NV_NVDLA_cbuf.scala 74:72:@1129.4]
  wire  _T_8174; // @[NV_NVDLA_cbuf.scala 74:72:@1131.4]
  wire  _T_8175; // @[NV_NVDLA_cbuf.scala 74:72:@1133.4]
  wire  _T_8176; // @[NV_NVDLA_cbuf.scala 74:72:@1135.4]
  wire  _T_8177; // @[NV_NVDLA_cbuf.scala 74:72:@1137.4]
  wire  _T_8178; // @[NV_NVDLA_cbuf.scala 74:72:@1139.4]
  wire  _T_8179; // @[NV_NVDLA_cbuf.scala 74:72:@1141.4]
  wire  _T_8180; // @[NV_NVDLA_cbuf.scala 74:72:@1143.4]
  wire  _T_8181; // @[NV_NVDLA_cbuf.scala 74:72:@1145.4]
  wire  _T_8182; // @[NV_NVDLA_cbuf.scala 74:72:@1147.4]
  reg [12:0] _T_8201_0; // @[NV_NVDLA_cbuf.scala 79:38:@1152.4]
  reg [31:0] _RAND_32;
  reg [12:0] _T_8201_1; // @[NV_NVDLA_cbuf.scala 79:38:@1152.4]
  reg [31:0] _RAND_33;
  reg [255:0] _T_8215_0; // @[NV_NVDLA_cbuf.scala 80:34:@1153.4]
  reg [255:0] _RAND_34;
  reg [255:0] _T_8215_1; // @[NV_NVDLA_cbuf.scala 80:34:@1153.4]
  reg [255:0] _RAND_35;
  reg  _T_9669_0_0; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_36;
  reg  _T_9669_0_1; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_37;
  reg  _T_9669_1_0; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_38;
  reg  _T_9669_1_1; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_39;
  reg  _T_9669_2_0; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_40;
  reg  _T_9669_2_1; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_41;
  reg  _T_9669_3_0; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_42;
  reg  _T_9669_3_1; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_43;
  reg  _T_9669_4_0; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_44;
  reg  _T_9669_4_1; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_45;
  reg  _T_9669_5_0; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_46;
  reg  _T_9669_5_1; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_47;
  reg  _T_9669_6_0; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_48;
  reg  _T_9669_6_1; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_49;
  reg  _T_9669_7_0; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_50;
  reg  _T_9669_7_1; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_51;
  reg  _T_9669_8_0; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_52;
  reg  _T_9669_8_1; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_53;
  reg  _T_9669_9_0; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_54;
  reg  _T_9669_9_1; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_55;
  reg  _T_9669_10_0; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_56;
  reg  _T_9669_10_1; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_57;
  reg  _T_9669_11_0; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_58;
  reg  _T_9669_11_1; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_59;
  reg  _T_9669_12_0; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_60;
  reg  _T_9669_12_1; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_61;
  reg  _T_9669_13_0; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_62;
  reg  _T_9669_13_1; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_63;
  reg  _T_9669_14_0; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_64;
  reg  _T_9669_14_1; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_65;
  reg  _T_9669_15_0; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_66;
  reg  _T_9669_15_1; // @[NV_NVDLA_cbuf.scala 86:32:@1239.4]
  reg [31:0] _RAND_67;
  wire  _T_10708; // @[NV_NVDLA_cbuf.scala 89:68:@1240.4]
  wire  _T_10709; // @[NV_NVDLA_cbuf.scala 89:68:@1242.4]
  wire  _T_10710; // @[NV_NVDLA_cbuf.scala 89:68:@1244.4]
  wire  _T_10711; // @[NV_NVDLA_cbuf.scala 89:68:@1246.4]
  wire  _T_10712; // @[NV_NVDLA_cbuf.scala 89:68:@1248.4]
  wire  _T_10713; // @[NV_NVDLA_cbuf.scala 89:68:@1250.4]
  wire  _T_10714; // @[NV_NVDLA_cbuf.scala 89:68:@1252.4]
  wire  _T_10715; // @[NV_NVDLA_cbuf.scala 89:68:@1254.4]
  wire  _T_10716; // @[NV_NVDLA_cbuf.scala 89:68:@1256.4]
  wire  _T_10717; // @[NV_NVDLA_cbuf.scala 89:68:@1258.4]
  wire  _T_10718; // @[NV_NVDLA_cbuf.scala 89:68:@1260.4]
  wire  _T_10719; // @[NV_NVDLA_cbuf.scala 89:68:@1262.4]
  wire  _T_10720; // @[NV_NVDLA_cbuf.scala 89:68:@1264.4]
  wire  _T_10721; // @[NV_NVDLA_cbuf.scala 89:68:@1266.4]
  wire  _T_10722; // @[NV_NVDLA_cbuf.scala 89:68:@1268.4]
  wire  _T_10723; // @[NV_NVDLA_cbuf.scala 89:68:@1270.4]
  wire  _T_10724; // @[NV_NVDLA_cbuf.scala 89:68:@1272.4]
  wire  _T_10725; // @[NV_NVDLA_cbuf.scala 89:68:@1274.4]
  wire  _T_10726; // @[NV_NVDLA_cbuf.scala 89:68:@1276.4]
  wire  _T_10727; // @[NV_NVDLA_cbuf.scala 89:68:@1278.4]
  wire  _T_10728; // @[NV_NVDLA_cbuf.scala 89:68:@1280.4]
  wire  _T_10729; // @[NV_NVDLA_cbuf.scala 89:68:@1282.4]
  wire  _T_10730; // @[NV_NVDLA_cbuf.scala 89:68:@1284.4]
  wire  _T_10731; // @[NV_NVDLA_cbuf.scala 89:68:@1286.4]
  wire  _T_10732; // @[NV_NVDLA_cbuf.scala 89:68:@1288.4]
  wire  _T_10733; // @[NV_NVDLA_cbuf.scala 89:68:@1290.4]
  wire  _T_10734; // @[NV_NVDLA_cbuf.scala 89:68:@1292.4]
  wire  _T_10735; // @[NV_NVDLA_cbuf.scala 89:68:@1294.4]
  wire  _T_10736; // @[NV_NVDLA_cbuf.scala 89:68:@1296.4]
  wire  _T_10737; // @[NV_NVDLA_cbuf.scala 89:68:@1298.4]
  wire  _T_10738; // @[NV_NVDLA_cbuf.scala 89:68:@1300.4]
  wire  _T_10739; // @[NV_NVDLA_cbuf.scala 89:68:@1302.4]
  wire [12:0] _T_11345; // @[Bitwise.scala 72:12:@1309.4]
  wire [12:0] _T_11346; // @[NV_NVDLA_cbuf.scala 101:94:@1310.4]
  wire [255:0] _T_11350; // @[Bitwise.scala 72:12:@1313.4]
  wire [255:0] _T_11351; // @[NV_NVDLA_cbuf.scala 102:97:@1314.4]
  wire [12:0] _T_11355; // @[Bitwise.scala 72:12:@1317.4]
  wire [12:0] _T_11356; // @[NV_NVDLA_cbuf.scala 101:94:@1318.4]
  wire [255:0] _T_11360; // @[Bitwise.scala 72:12:@1321.4]
  wire [255:0] _T_11361; // @[NV_NVDLA_cbuf.scala 102:97:@1322.4]
  wire [12:0] _T_11362; // @[NV_NVDLA_cbuf.scala 104:68:@1324.4]
  wire [12:0] _T_11367; // @[Bitwise.scala 72:12:@1329.4]
  wire [12:0] _T_11368; // @[NV_NVDLA_cbuf.scala 101:94:@1330.4]
  wire [255:0] _T_11372; // @[Bitwise.scala 72:12:@1333.4]
  wire [255:0] _T_11373; // @[NV_NVDLA_cbuf.scala 102:97:@1334.4]
  wire [12:0] _T_11377; // @[Bitwise.scala 72:12:@1337.4]
  wire [12:0] _T_11378; // @[NV_NVDLA_cbuf.scala 101:94:@1338.4]
  wire [255:0] _T_11382; // @[Bitwise.scala 72:12:@1341.4]
  wire [255:0] _T_11383; // @[NV_NVDLA_cbuf.scala 102:97:@1342.4]
  wire [12:0] _T_11384; // @[NV_NVDLA_cbuf.scala 104:68:@1344.4]
  wire [12:0] _T_11389; // @[Bitwise.scala 72:12:@1349.4]
  wire [12:0] _T_11390; // @[NV_NVDLA_cbuf.scala 101:94:@1350.4]
  wire [255:0] _T_11394; // @[Bitwise.scala 72:12:@1353.4]
  wire [255:0] _T_11395; // @[NV_NVDLA_cbuf.scala 102:97:@1354.4]
  wire [12:0] _T_11399; // @[Bitwise.scala 72:12:@1357.4]
  wire [12:0] _T_11400; // @[NV_NVDLA_cbuf.scala 101:94:@1358.4]
  wire [255:0] _T_11404; // @[Bitwise.scala 72:12:@1361.4]
  wire [255:0] _T_11405; // @[NV_NVDLA_cbuf.scala 102:97:@1362.4]
  wire [12:0] _T_11406; // @[NV_NVDLA_cbuf.scala 104:68:@1364.4]
  wire [12:0] _T_11411; // @[Bitwise.scala 72:12:@1369.4]
  wire [12:0] _T_11412; // @[NV_NVDLA_cbuf.scala 101:94:@1370.4]
  wire [255:0] _T_11416; // @[Bitwise.scala 72:12:@1373.4]
  wire [255:0] _T_11417; // @[NV_NVDLA_cbuf.scala 102:97:@1374.4]
  wire [12:0] _T_11421; // @[Bitwise.scala 72:12:@1377.4]
  wire [12:0] _T_11422; // @[NV_NVDLA_cbuf.scala 101:94:@1378.4]
  wire [255:0] _T_11426; // @[Bitwise.scala 72:12:@1381.4]
  wire [255:0] _T_11427; // @[NV_NVDLA_cbuf.scala 102:97:@1382.4]
  wire [12:0] _T_11428; // @[NV_NVDLA_cbuf.scala 104:68:@1384.4]
  wire [12:0] _T_11433; // @[Bitwise.scala 72:12:@1389.4]
  wire [12:0] _T_11434; // @[NV_NVDLA_cbuf.scala 101:94:@1390.4]
  wire [255:0] _T_11438; // @[Bitwise.scala 72:12:@1393.4]
  wire [255:0] _T_11439; // @[NV_NVDLA_cbuf.scala 102:97:@1394.4]
  wire [12:0] _T_11443; // @[Bitwise.scala 72:12:@1397.4]
  wire [12:0] _T_11444; // @[NV_NVDLA_cbuf.scala 101:94:@1398.4]
  wire [255:0] _T_11448; // @[Bitwise.scala 72:12:@1401.4]
  wire [255:0] _T_11449; // @[NV_NVDLA_cbuf.scala 102:97:@1402.4]
  wire [12:0] _T_11450; // @[NV_NVDLA_cbuf.scala 104:68:@1404.4]
  wire [12:0] _T_11455; // @[Bitwise.scala 72:12:@1409.4]
  wire [12:0] _T_11456; // @[NV_NVDLA_cbuf.scala 101:94:@1410.4]
  wire [255:0] _T_11460; // @[Bitwise.scala 72:12:@1413.4]
  wire [255:0] _T_11461; // @[NV_NVDLA_cbuf.scala 102:97:@1414.4]
  wire [12:0] _T_11465; // @[Bitwise.scala 72:12:@1417.4]
  wire [12:0] _T_11466; // @[NV_NVDLA_cbuf.scala 101:94:@1418.4]
  wire [255:0] _T_11470; // @[Bitwise.scala 72:12:@1421.4]
  wire [255:0] _T_11471; // @[NV_NVDLA_cbuf.scala 102:97:@1422.4]
  wire [12:0] _T_11472; // @[NV_NVDLA_cbuf.scala 104:68:@1424.4]
  wire [12:0] _T_11477; // @[Bitwise.scala 72:12:@1429.4]
  wire [12:0] _T_11478; // @[NV_NVDLA_cbuf.scala 101:94:@1430.4]
  wire [255:0] _T_11482; // @[Bitwise.scala 72:12:@1433.4]
  wire [255:0] _T_11483; // @[NV_NVDLA_cbuf.scala 102:97:@1434.4]
  wire [12:0] _T_11487; // @[Bitwise.scala 72:12:@1437.4]
  wire [12:0] _T_11488; // @[NV_NVDLA_cbuf.scala 101:94:@1438.4]
  wire [255:0] _T_11492; // @[Bitwise.scala 72:12:@1441.4]
  wire [255:0] _T_11493; // @[NV_NVDLA_cbuf.scala 102:97:@1442.4]
  wire [12:0] _T_11494; // @[NV_NVDLA_cbuf.scala 104:68:@1444.4]
  wire [12:0] _T_11499; // @[Bitwise.scala 72:12:@1449.4]
  wire [12:0] _T_11500; // @[NV_NVDLA_cbuf.scala 101:94:@1450.4]
  wire [255:0] _T_11504; // @[Bitwise.scala 72:12:@1453.4]
  wire [255:0] _T_11505; // @[NV_NVDLA_cbuf.scala 102:97:@1454.4]
  wire [12:0] _T_11509; // @[Bitwise.scala 72:12:@1457.4]
  wire [12:0] _T_11510; // @[NV_NVDLA_cbuf.scala 101:94:@1458.4]
  wire [255:0] _T_11514; // @[Bitwise.scala 72:12:@1461.4]
  wire [255:0] _T_11515; // @[NV_NVDLA_cbuf.scala 102:97:@1462.4]
  wire [12:0] _T_11516; // @[NV_NVDLA_cbuf.scala 104:68:@1464.4]
  wire [12:0] _T_11521; // @[Bitwise.scala 72:12:@1469.4]
  wire [12:0] _T_11522; // @[NV_NVDLA_cbuf.scala 101:94:@1470.4]
  wire [255:0] _T_11526; // @[Bitwise.scala 72:12:@1473.4]
  wire [255:0] _T_11527; // @[NV_NVDLA_cbuf.scala 102:97:@1474.4]
  wire [12:0] _T_11531; // @[Bitwise.scala 72:12:@1477.4]
  wire [12:0] _T_11532; // @[NV_NVDLA_cbuf.scala 101:94:@1478.4]
  wire [255:0] _T_11536; // @[Bitwise.scala 72:12:@1481.4]
  wire [255:0] _T_11537; // @[NV_NVDLA_cbuf.scala 102:97:@1482.4]
  wire [12:0] _T_11538; // @[NV_NVDLA_cbuf.scala 104:68:@1484.4]
  wire [12:0] _T_11543; // @[Bitwise.scala 72:12:@1489.4]
  wire [12:0] _T_11544; // @[NV_NVDLA_cbuf.scala 101:94:@1490.4]
  wire [255:0] _T_11548; // @[Bitwise.scala 72:12:@1493.4]
  wire [255:0] _T_11549; // @[NV_NVDLA_cbuf.scala 102:97:@1494.4]
  wire [12:0] _T_11553; // @[Bitwise.scala 72:12:@1497.4]
  wire [12:0] _T_11554; // @[NV_NVDLA_cbuf.scala 101:94:@1498.4]
  wire [255:0] _T_11558; // @[Bitwise.scala 72:12:@1501.4]
  wire [255:0] _T_11559; // @[NV_NVDLA_cbuf.scala 102:97:@1502.4]
  wire [12:0] _T_11560; // @[NV_NVDLA_cbuf.scala 104:68:@1504.4]
  wire [12:0] _T_11565; // @[Bitwise.scala 72:12:@1509.4]
  wire [12:0] _T_11566; // @[NV_NVDLA_cbuf.scala 101:94:@1510.4]
  wire [255:0] _T_11570; // @[Bitwise.scala 72:12:@1513.4]
  wire [255:0] _T_11571; // @[NV_NVDLA_cbuf.scala 102:97:@1514.4]
  wire [12:0] _T_11575; // @[Bitwise.scala 72:12:@1517.4]
  wire [12:0] _T_11576; // @[NV_NVDLA_cbuf.scala 101:94:@1518.4]
  wire [255:0] _T_11580; // @[Bitwise.scala 72:12:@1521.4]
  wire [255:0] _T_11581; // @[NV_NVDLA_cbuf.scala 102:97:@1522.4]
  wire [12:0] _T_11582; // @[NV_NVDLA_cbuf.scala 104:68:@1524.4]
  wire [12:0] _T_11587; // @[Bitwise.scala 72:12:@1529.4]
  wire [12:0] _T_11588; // @[NV_NVDLA_cbuf.scala 101:94:@1530.4]
  wire [255:0] _T_11592; // @[Bitwise.scala 72:12:@1533.4]
  wire [255:0] _T_11593; // @[NV_NVDLA_cbuf.scala 102:97:@1534.4]
  wire [12:0] _T_11597; // @[Bitwise.scala 72:12:@1537.4]
  wire [12:0] _T_11598; // @[NV_NVDLA_cbuf.scala 101:94:@1538.4]
  wire [255:0] _T_11602; // @[Bitwise.scala 72:12:@1541.4]
  wire [255:0] _T_11603; // @[NV_NVDLA_cbuf.scala 102:97:@1542.4]
  wire [12:0] _T_11604; // @[NV_NVDLA_cbuf.scala 104:68:@1544.4]
  wire [12:0] _T_11609; // @[Bitwise.scala 72:12:@1549.4]
  wire [12:0] _T_11610; // @[NV_NVDLA_cbuf.scala 101:94:@1550.4]
  wire [255:0] _T_11614; // @[Bitwise.scala 72:12:@1553.4]
  wire [255:0] _T_11615; // @[NV_NVDLA_cbuf.scala 102:97:@1554.4]
  wire [12:0] _T_11619; // @[Bitwise.scala 72:12:@1557.4]
  wire [12:0] _T_11620; // @[NV_NVDLA_cbuf.scala 101:94:@1558.4]
  wire [255:0] _T_11624; // @[Bitwise.scala 72:12:@1561.4]
  wire [255:0] _T_11625; // @[NV_NVDLA_cbuf.scala 102:97:@1562.4]
  wire [12:0] _T_11626; // @[NV_NVDLA_cbuf.scala 104:68:@1564.4]
  wire [12:0] _T_11631; // @[Bitwise.scala 72:12:@1569.4]
  wire [12:0] _T_11632; // @[NV_NVDLA_cbuf.scala 101:94:@1570.4]
  wire [255:0] _T_11636; // @[Bitwise.scala 72:12:@1573.4]
  wire [255:0] _T_11637; // @[NV_NVDLA_cbuf.scala 102:97:@1574.4]
  wire [12:0] _T_11641; // @[Bitwise.scala 72:12:@1577.4]
  wire [12:0] _T_11642; // @[NV_NVDLA_cbuf.scala 101:94:@1578.4]
  wire [255:0] _T_11646; // @[Bitwise.scala 72:12:@1581.4]
  wire [255:0] _T_11647; // @[NV_NVDLA_cbuf.scala 102:97:@1582.4]
  wire [12:0] _T_11648; // @[NV_NVDLA_cbuf.scala 104:68:@1584.4]
  wire [12:0] _T_11653; // @[Bitwise.scala 72:12:@1589.4]
  wire [12:0] _T_11654; // @[NV_NVDLA_cbuf.scala 101:94:@1590.4]
  wire [255:0] _T_11658; // @[Bitwise.scala 72:12:@1593.4]
  wire [255:0] _T_11659; // @[NV_NVDLA_cbuf.scala 102:97:@1594.4]
  wire [12:0] _T_11663; // @[Bitwise.scala 72:12:@1597.4]
  wire [12:0] _T_11664; // @[NV_NVDLA_cbuf.scala 101:94:@1598.4]
  wire [255:0] _T_11668; // @[Bitwise.scala 72:12:@1601.4]
  wire [255:0] _T_11669; // @[NV_NVDLA_cbuf.scala 102:97:@1602.4]
  wire [12:0] _T_11670; // @[NV_NVDLA_cbuf.scala 104:68:@1604.4]
  wire [12:0] _T_11675; // @[Bitwise.scala 72:12:@1609.4]
  wire [12:0] _T_11676; // @[NV_NVDLA_cbuf.scala 101:94:@1610.4]
  wire [255:0] _T_11680; // @[Bitwise.scala 72:12:@1613.4]
  wire [255:0] _T_11681; // @[NV_NVDLA_cbuf.scala 102:97:@1614.4]
  wire [12:0] _T_11685; // @[Bitwise.scala 72:12:@1617.4]
  wire [12:0] _T_11686; // @[NV_NVDLA_cbuf.scala 101:94:@1618.4]
  wire [255:0] _T_11690; // @[Bitwise.scala 72:12:@1621.4]
  wire [255:0] _T_11691; // @[NV_NVDLA_cbuf.scala 102:97:@1622.4]
  wire [12:0] _T_11692; // @[NV_NVDLA_cbuf.scala 104:68:@1624.4]
  wire [8:0] _T_12252; // @[NV_NVDLA_cbuf.scala 114:63:@1630.4]
  wire [8:0] _T_12254; // @[NV_NVDLA_cbuf.scala 114:63:@1636.4]
  wire [8:0] _T_12256; // @[NV_NVDLA_cbuf.scala 114:63:@1642.4]
  wire [8:0] _T_12258; // @[NV_NVDLA_cbuf.scala 114:63:@1648.4]
  wire [8:0] _T_12260; // @[NV_NVDLA_cbuf.scala 114:63:@1654.4]
  wire [8:0] _T_12262; // @[NV_NVDLA_cbuf.scala 114:63:@1660.4]
  wire [8:0] _T_12264; // @[NV_NVDLA_cbuf.scala 114:63:@1666.4]
  wire [8:0] _T_12266; // @[NV_NVDLA_cbuf.scala 114:63:@1672.4]
  wire [8:0] _T_12268; // @[NV_NVDLA_cbuf.scala 114:63:@1678.4]
  wire [8:0] _T_12270; // @[NV_NVDLA_cbuf.scala 114:63:@1684.4]
  wire [8:0] _T_12272; // @[NV_NVDLA_cbuf.scala 114:63:@1690.4]
  wire [8:0] _T_12274; // @[NV_NVDLA_cbuf.scala 114:63:@1696.4]
  wire [8:0] _T_12276; // @[NV_NVDLA_cbuf.scala 114:63:@1702.4]
  wire [8:0] _T_12278; // @[NV_NVDLA_cbuf.scala 114:63:@1708.4]
  wire [8:0] _T_12280; // @[NV_NVDLA_cbuf.scala 114:63:@1714.4]
  wire [8:0] _T_12282; // @[NV_NVDLA_cbuf.scala 114:63:@1720.4]
  reg [8:0] _T_13733_0_0; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_68;
  reg [8:0] _T_13733_0_1; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_69;
  reg [8:0] _T_13733_1_0; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_70;
  reg [8:0] _T_13733_1_1; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_71;
  reg [8:0] _T_13733_2_0; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_72;
  reg [8:0] _T_13733_2_1; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_73;
  reg [8:0] _T_13733_3_0; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_74;
  reg [8:0] _T_13733_3_1; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_75;
  reg [8:0] _T_13733_4_0; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_76;
  reg [8:0] _T_13733_4_1; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_77;
  reg [8:0] _T_13733_5_0; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_78;
  reg [8:0] _T_13733_5_1; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_79;
  reg [8:0] _T_13733_6_0; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_80;
  reg [8:0] _T_13733_6_1; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_81;
  reg [8:0] _T_13733_7_0; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_82;
  reg [8:0] _T_13733_7_1; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_83;
  reg [8:0] _T_13733_8_0; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_84;
  reg [8:0] _T_13733_8_1; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_85;
  reg [8:0] _T_13733_9_0; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_86;
  reg [8:0] _T_13733_9_1; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_87;
  reg [8:0] _T_13733_10_0; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_88;
  reg [8:0] _T_13733_10_1; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_89;
  reg [8:0] _T_13733_11_0; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_90;
  reg [8:0] _T_13733_11_1; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_91;
  reg [8:0] _T_13733_12_0; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_92;
  reg [8:0] _T_13733_12_1; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_93;
  reg [8:0] _T_13733_13_0; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_94;
  reg [8:0] _T_13733_13_1; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_95;
  reg [8:0] _T_13733_14_0; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_96;
  reg [8:0] _T_13733_14_1; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_97;
  reg [8:0] _T_13733_15_0; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_98;
  reg [8:0] _T_13733_15_1; // @[NV_NVDLA_cbuf.scala 125:38:@1807.4]
  reg [31:0] _RAND_99;
  reg [255:0] _T_14845_0_0; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_100;
  reg [255:0] _T_14845_0_1; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_101;
  reg [255:0] _T_14845_1_0; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_102;
  reg [255:0] _T_14845_1_1; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_103;
  reg [255:0] _T_14845_2_0; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_104;
  reg [255:0] _T_14845_2_1; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_105;
  reg [255:0] _T_14845_3_0; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_106;
  reg [255:0] _T_14845_3_1; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_107;
  reg [255:0] _T_14845_4_0; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_108;
  reg [255:0] _T_14845_4_1; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_109;
  reg [255:0] _T_14845_5_0; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_110;
  reg [255:0] _T_14845_5_1; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_111;
  reg [255:0] _T_14845_6_0; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_112;
  reg [255:0] _T_14845_6_1; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_113;
  reg [255:0] _T_14845_7_0; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_114;
  reg [255:0] _T_14845_7_1; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_115;
  reg [255:0] _T_14845_8_0; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_116;
  reg [255:0] _T_14845_8_1; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_117;
  reg [255:0] _T_14845_9_0; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_118;
  reg [255:0] _T_14845_9_1; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_119;
  reg [255:0] _T_14845_10_0; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_120;
  reg [255:0] _T_14845_10_1; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_121;
  reg [255:0] _T_14845_11_0; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_122;
  reg [255:0] _T_14845_11_1; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_123;
  reg [255:0] _T_14845_12_0; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_124;
  reg [255:0] _T_14845_12_1; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_125;
  reg [255:0] _T_14845_13_0; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_126;
  reg [255:0] _T_14845_13_1; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_127;
  reg [255:0] _T_14845_14_0; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_128;
  reg [255:0] _T_14845_14_1; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_129;
  reg [255:0] _T_14845_15_0; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_130;
  reg [255:0] _T_14845_15_1; // @[NV_NVDLA_cbuf.scala 126:34:@1808.4]
  reg [255:0] _RAND_131;
  reg  _T_16500_0_0; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_132;
  reg  _T_16500_0_1; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_133;
  reg  _T_16500_1_0; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_134;
  reg  _T_16500_1_1; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_135;
  reg  _T_16500_2_0; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_136;
  reg  _T_16500_2_1; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_137;
  reg  _T_16500_3_0; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_138;
  reg  _T_16500_3_1; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_139;
  reg  _T_16500_4_0; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_140;
  reg  _T_16500_4_1; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_141;
  reg  _T_16500_5_0; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_142;
  reg  _T_16500_5_1; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_143;
  reg  _T_16500_6_0; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_144;
  reg  _T_16500_6_1; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_145;
  reg  _T_16500_7_0; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_146;
  reg  _T_16500_7_1; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_147;
  reg  _T_16500_8_0; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_148;
  reg  _T_16500_8_1; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_149;
  reg  _T_16500_9_0; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_150;
  reg  _T_16500_9_1; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_151;
  reg  _T_16500_10_0; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_152;
  reg  _T_16500_10_1; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_153;
  reg  _T_16500_11_0; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_154;
  reg  _T_16500_11_1; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_155;
  reg  _T_16500_12_0; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_156;
  reg  _T_16500_12_1; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_157;
  reg  _T_16500_13_0; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_158;
  reg  _T_16500_13_1; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_159;
  reg  _T_16500_14_0; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_160;
  reg  _T_16500_14_1; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_161;
  reg  _T_16500_15_0; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_162;
  reg  _T_16500_15_1; // @[NV_NVDLA_cbuf.scala 127:36:@1890.4]
  reg [31:0] _RAND_163;
  wire [3:0] _T_19410; // @[NV_NVDLA_cbuf.scala 140:107:@1988.4]
  wire  _T_19412; // @[NV_NVDLA_cbuf.scala 140:158:@1989.4]
  wire  _T_19413; // @[NV_NVDLA_cbuf.scala 140:78:@1990.4]
  wire  _T_19420; // @[NV_NVDLA_cbuf.scala 140:158:@1997.4]
  wire  _T_19421; // @[NV_NVDLA_cbuf.scala 140:78:@1998.4]
  wire  _T_19428; // @[NV_NVDLA_cbuf.scala 140:158:@2005.4]
  wire  _T_19429; // @[NV_NVDLA_cbuf.scala 140:78:@2006.4]
  wire  _T_19436; // @[NV_NVDLA_cbuf.scala 140:158:@2013.4]
  wire  _T_19437; // @[NV_NVDLA_cbuf.scala 140:78:@2014.4]
  wire  _T_19444; // @[NV_NVDLA_cbuf.scala 140:158:@2021.4]
  wire  _T_19445; // @[NV_NVDLA_cbuf.scala 140:78:@2022.4]
  wire  _T_19452; // @[NV_NVDLA_cbuf.scala 140:158:@2029.4]
  wire  _T_19453; // @[NV_NVDLA_cbuf.scala 140:78:@2030.4]
  wire  _T_19460; // @[NV_NVDLA_cbuf.scala 140:158:@2037.4]
  wire  _T_19461; // @[NV_NVDLA_cbuf.scala 140:78:@2038.4]
  wire  _T_19468; // @[NV_NVDLA_cbuf.scala 140:158:@2045.4]
  wire  _T_19469; // @[NV_NVDLA_cbuf.scala 140:78:@2046.4]
  wire  _T_19476; // @[NV_NVDLA_cbuf.scala 140:158:@2053.4]
  wire  _T_19477; // @[NV_NVDLA_cbuf.scala 140:78:@2054.4]
  wire  _T_19484; // @[NV_NVDLA_cbuf.scala 140:158:@2061.4]
  wire  _T_19485; // @[NV_NVDLA_cbuf.scala 140:78:@2062.4]
  wire  _T_19492; // @[NV_NVDLA_cbuf.scala 140:158:@2069.4]
  wire  _T_19493; // @[NV_NVDLA_cbuf.scala 140:78:@2070.4]
  wire  _T_19500; // @[NV_NVDLA_cbuf.scala 140:158:@2077.4]
  wire  _T_19501; // @[NV_NVDLA_cbuf.scala 140:78:@2078.4]
  wire  _T_19508; // @[NV_NVDLA_cbuf.scala 140:158:@2085.4]
  wire  _T_19509; // @[NV_NVDLA_cbuf.scala 140:78:@2086.4]
  wire  _T_19516; // @[NV_NVDLA_cbuf.scala 140:158:@2093.4]
  wire  _T_19517; // @[NV_NVDLA_cbuf.scala 140:78:@2094.4]
  wire  _T_19524; // @[NV_NVDLA_cbuf.scala 140:158:@2101.4]
  wire  _T_19525; // @[NV_NVDLA_cbuf.scala 140:78:@2102.4]
  wire  _T_19532; // @[NV_NVDLA_cbuf.scala 140:158:@2109.4]
  wire  _T_19533; // @[NV_NVDLA_cbuf.scala 140:78:@2110.4]
  wire [8:0] _T_21412; // @[Bitwise.scala 72:12:@2118.4]
  wire [8:0] _T_21413; // @[NV_NVDLA_cbuf.scala 160:139:@2119.4]
  wire [8:0] _T_21414; // @[NV_NVDLA_cbuf.scala 160:111:@2120.4]
  wire [8:0] _T_21424; // @[Bitwise.scala 72:12:@2128.4]
  wire [8:0] _T_21426; // @[NV_NVDLA_cbuf.scala 160:111:@2130.4]
  wire [8:0] _T_21436; // @[Bitwise.scala 72:12:@2138.4]
  wire [8:0] _T_21438; // @[NV_NVDLA_cbuf.scala 160:111:@2140.4]
  wire [8:0] _T_21448; // @[Bitwise.scala 72:12:@2148.4]
  wire [8:0] _T_21450; // @[NV_NVDLA_cbuf.scala 160:111:@2150.4]
  wire [8:0] _T_21460; // @[Bitwise.scala 72:12:@2158.4]
  wire [8:0] _T_21462; // @[NV_NVDLA_cbuf.scala 160:111:@2160.4]
  wire [8:0] _T_21472; // @[Bitwise.scala 72:12:@2168.4]
  wire [8:0] _T_21474; // @[NV_NVDLA_cbuf.scala 160:111:@2170.4]
  wire [8:0] _T_21484; // @[Bitwise.scala 72:12:@2178.4]
  wire [8:0] _T_21486; // @[NV_NVDLA_cbuf.scala 160:111:@2180.4]
  wire [8:0] _T_21496; // @[Bitwise.scala 72:12:@2188.4]
  wire [8:0] _T_21498; // @[NV_NVDLA_cbuf.scala 160:111:@2190.4]
  wire [8:0] _T_21508; // @[Bitwise.scala 72:12:@2198.4]
  wire [8:0] _T_21510; // @[NV_NVDLA_cbuf.scala 160:111:@2200.4]
  wire [8:0] _T_21520; // @[Bitwise.scala 72:12:@2208.4]
  wire [8:0] _T_21522; // @[NV_NVDLA_cbuf.scala 160:111:@2210.4]
  wire [8:0] _T_21532; // @[Bitwise.scala 72:12:@2218.4]
  wire [8:0] _T_21534; // @[NV_NVDLA_cbuf.scala 160:111:@2220.4]
  wire [8:0] _T_21544; // @[Bitwise.scala 72:12:@2228.4]
  wire [8:0] _T_21546; // @[NV_NVDLA_cbuf.scala 160:111:@2230.4]
  wire [8:0] _T_21556; // @[Bitwise.scala 72:12:@2238.4]
  wire [8:0] _T_21558; // @[NV_NVDLA_cbuf.scala 160:111:@2240.4]
  wire [8:0] _T_21568; // @[Bitwise.scala 72:12:@2248.4]
  wire [8:0] _T_21570; // @[NV_NVDLA_cbuf.scala 160:111:@2250.4]
  wire [8:0] _T_21580; // @[Bitwise.scala 72:12:@2258.4]
  wire [8:0] _T_21582; // @[NV_NVDLA_cbuf.scala 160:111:@2260.4]
  wire [8:0] _T_21592; // @[Bitwise.scala 72:12:@2268.4]
  wire [8:0] _T_21594; // @[NV_NVDLA_cbuf.scala 160:111:@2270.4]
  reg  _T_39941_0_0_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_164;
  reg  _T_39941_0_1_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_165;
  reg  _T_39941_1_0_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_166;
  reg  _T_39941_1_1_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_167;
  reg  _T_39941_2_0_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_168;
  reg  _T_39941_2_1_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_169;
  reg  _T_39941_3_0_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_170;
  reg  _T_39941_3_1_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_171;
  reg  _T_39941_4_0_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_172;
  reg  _T_39941_4_1_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_173;
  reg  _T_39941_5_0_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_174;
  reg  _T_39941_5_1_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_175;
  reg  _T_39941_6_0_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_176;
  reg  _T_39941_6_1_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_177;
  reg  _T_39941_7_0_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_178;
  reg  _T_39941_7_1_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_179;
  reg  _T_39941_8_0_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_180;
  reg  _T_39941_8_1_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_181;
  reg  _T_39941_9_0_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_182;
  reg  _T_39941_9_1_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_183;
  reg  _T_39941_10_0_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_184;
  reg  _T_39941_10_1_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_185;
  reg  _T_39941_11_0_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_186;
  reg  _T_39941_11_1_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_187;
  reg  _T_39941_12_0_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_188;
  reg  _T_39941_12_1_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_189;
  reg  _T_39941_13_0_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_190;
  reg  _T_39941_13_1_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_191;
  reg  _T_39941_14_0_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_192;
  reg  _T_39941_14_1_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_193;
  reg  _T_39941_15_0_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_194;
  reg  _T_39941_15_1_0; // @[NV_NVDLA_cbuf.scala 170:41:@2422.4]
  reg [31:0] _RAND_195;
  reg  _T_72478_0_0_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_196;
  reg  _T_72478_0_1_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_197;
  reg  _T_72478_1_0_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_198;
  reg  _T_72478_1_1_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_199;
  reg  _T_72478_2_0_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_200;
  reg  _T_72478_2_1_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_201;
  reg  _T_72478_3_0_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_202;
  reg  _T_72478_3_1_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_203;
  reg  _T_72478_4_0_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_204;
  reg  _T_72478_4_1_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_205;
  reg  _T_72478_5_0_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_206;
  reg  _T_72478_5_1_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_207;
  reg  _T_72478_6_0_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_208;
  reg  _T_72478_6_1_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_209;
  reg  _T_72478_7_0_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_210;
  reg  _T_72478_7_1_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_211;
  reg  _T_72478_8_0_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_212;
  reg  _T_72478_8_1_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_213;
  reg  _T_72478_9_0_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_214;
  reg  _T_72478_9_1_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_215;
  reg  _T_72478_10_0_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_216;
  reg  _T_72478_10_1_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_217;
  reg  _T_72478_11_0_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_218;
  reg  _T_72478_11_1_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_219;
  reg  _T_72478_12_0_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_220;
  reg  _T_72478_12_1_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_221;
  reg  _T_72478_13_0_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_222;
  reg  _T_72478_13_1_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_223;
  reg  _T_72478_14_0_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_224;
  reg  _T_72478_14_1_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_225;
  reg  _T_72478_15_0_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_226;
  reg  _T_72478_15_1_0; // @[NV_NVDLA_cbuf.scala 171:41:@2568.4]
  reg [31:0] _RAND_227;
  wire [7:0] _T_86681; // @[NV_NVDLA_cbuf.scala 177:73:@2639.4]
  wire [15:0] _T_86689; // @[NV_NVDLA_cbuf.scala 177:73:@2647.4]
  wire [7:0] _T_86696; // @[NV_NVDLA_cbuf.scala 177:73:@2654.4]
  wire [31:0] _T_86705; // @[NV_NVDLA_cbuf.scala 177:73:@2663.4]
  reg  _T_86710; // @[Reg.scala 11:16:@2665.4]
  reg [31:0] _RAND_228;
  reg  _T_86712; // @[Reg.scala 11:16:@2669.4]
  reg [31:0] _RAND_229;
  reg  _T_86714; // @[Reg.scala 11:16:@2673.4]
  reg [31:0] _RAND_230;
  reg  _T_86716; // @[Reg.scala 11:16:@2677.4]
  reg [31:0] _RAND_231;
  wire [255:0] _T_87210; // @[Bitwise.scala 72:12:@2685.4]
  wire [255:0] _T_86790_0_1; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@3950.4]
  wire [255:0] _T_87211; // @[NV_NVDLA_cbuf.scala 197:68:@2686.4]
  wire [255:0] _T_87215; // @[Bitwise.scala 72:12:@2688.4]
  wire [255:0] _T_86790_0_0; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@3941.4]
  wire [255:0] _T_87216; // @[NV_NVDLA_cbuf.scala 198:65:@2689.4]
  wire [255:0] _T_87221; // @[Bitwise.scala 72:12:@2693.4]
  wire [255:0] _T_86790_1_1; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@3968.4]
  wire [255:0] _T_87222; // @[NV_NVDLA_cbuf.scala 197:68:@2694.4]
  wire [255:0] _T_87226; // @[Bitwise.scala 72:12:@2696.4]
  wire [255:0] _T_86790_1_0; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@3959.4]
  wire [255:0] _T_87227; // @[NV_NVDLA_cbuf.scala 198:65:@2697.4]
  wire [255:0] _T_87232; // @[Bitwise.scala 72:12:@2701.4]
  wire [255:0] _T_86790_2_1; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@3986.4]
  wire [255:0] _T_87233; // @[NV_NVDLA_cbuf.scala 197:68:@2702.4]
  wire [255:0] _T_87237; // @[Bitwise.scala 72:12:@2704.4]
  wire [255:0] _T_86790_2_0; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@3977.4]
  wire [255:0] _T_87238; // @[NV_NVDLA_cbuf.scala 198:65:@2705.4]
  wire [255:0] _T_87243; // @[Bitwise.scala 72:12:@2709.4]
  wire [255:0] _T_86790_3_1; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4004.4]
  wire [255:0] _T_87244; // @[NV_NVDLA_cbuf.scala 197:68:@2710.4]
  wire [255:0] _T_87248; // @[Bitwise.scala 72:12:@2712.4]
  wire [255:0] _T_86790_3_0; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@3995.4]
  wire [255:0] _T_87249; // @[NV_NVDLA_cbuf.scala 198:65:@2713.4]
  wire [255:0] _T_87254; // @[Bitwise.scala 72:12:@2717.4]
  wire [255:0] _T_86790_4_1; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4022.4]
  wire [255:0] _T_87255; // @[NV_NVDLA_cbuf.scala 197:68:@2718.4]
  wire [255:0] _T_87259; // @[Bitwise.scala 72:12:@2720.4]
  wire [255:0] _T_86790_4_0; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4013.4]
  wire [255:0] _T_87260; // @[NV_NVDLA_cbuf.scala 198:65:@2721.4]
  wire [255:0] _T_87265; // @[Bitwise.scala 72:12:@2725.4]
  wire [255:0] _T_86790_5_1; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4040.4]
  wire [255:0] _T_87266; // @[NV_NVDLA_cbuf.scala 197:68:@2726.4]
  wire [255:0] _T_87270; // @[Bitwise.scala 72:12:@2728.4]
  wire [255:0] _T_86790_5_0; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4031.4]
  wire [255:0] _T_87271; // @[NV_NVDLA_cbuf.scala 198:65:@2729.4]
  wire [255:0] _T_87276; // @[Bitwise.scala 72:12:@2733.4]
  wire [255:0] _T_86790_6_1; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4058.4]
  wire [255:0] _T_87277; // @[NV_NVDLA_cbuf.scala 197:68:@2734.4]
  wire [255:0] _T_87281; // @[Bitwise.scala 72:12:@2736.4]
  wire [255:0] _T_86790_6_0; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4049.4]
  wire [255:0] _T_87282; // @[NV_NVDLA_cbuf.scala 198:65:@2737.4]
  wire [255:0] _T_87287; // @[Bitwise.scala 72:12:@2741.4]
  wire [255:0] _T_86790_7_1; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4076.4]
  wire [255:0] _T_87288; // @[NV_NVDLA_cbuf.scala 197:68:@2742.4]
  wire [255:0] _T_87292; // @[Bitwise.scala 72:12:@2744.4]
  wire [255:0] _T_86790_7_0; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4067.4]
  wire [255:0] _T_87293; // @[NV_NVDLA_cbuf.scala 198:65:@2745.4]
  wire [255:0] _T_87298; // @[Bitwise.scala 72:12:@2749.4]
  wire [255:0] _T_86790_8_1; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4094.4]
  wire [255:0] _T_87299; // @[NV_NVDLA_cbuf.scala 197:68:@2750.4]
  wire [255:0] _T_87303; // @[Bitwise.scala 72:12:@2752.4]
  wire [255:0] _T_86790_8_0; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4085.4]
  wire [255:0] _T_87304; // @[NV_NVDLA_cbuf.scala 198:65:@2753.4]
  wire [255:0] _T_87309; // @[Bitwise.scala 72:12:@2757.4]
  wire [255:0] _T_86790_9_1; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4112.4]
  wire [255:0] _T_87310; // @[NV_NVDLA_cbuf.scala 197:68:@2758.4]
  wire [255:0] _T_87314; // @[Bitwise.scala 72:12:@2760.4]
  wire [255:0] _T_86790_9_0; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4103.4]
  wire [255:0] _T_87315; // @[NV_NVDLA_cbuf.scala 198:65:@2761.4]
  wire [255:0] _T_87320; // @[Bitwise.scala 72:12:@2765.4]
  wire [255:0] _T_86790_10_1; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4130.4]
  wire [255:0] _T_87321; // @[NV_NVDLA_cbuf.scala 197:68:@2766.4]
  wire [255:0] _T_87325; // @[Bitwise.scala 72:12:@2768.4]
  wire [255:0] _T_86790_10_0; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4121.4]
  wire [255:0] _T_87326; // @[NV_NVDLA_cbuf.scala 198:65:@2769.4]
  wire [255:0] _T_87331; // @[Bitwise.scala 72:12:@2773.4]
  wire [255:0] _T_86790_11_1; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4148.4]
  wire [255:0] _T_87332; // @[NV_NVDLA_cbuf.scala 197:68:@2774.4]
  wire [255:0] _T_87336; // @[Bitwise.scala 72:12:@2776.4]
  wire [255:0] _T_86790_11_0; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4139.4]
  wire [255:0] _T_87337; // @[NV_NVDLA_cbuf.scala 198:65:@2777.4]
  wire [255:0] _T_87342; // @[Bitwise.scala 72:12:@2781.4]
  wire [255:0] _T_86790_12_1; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4166.4]
  wire [255:0] _T_87343; // @[NV_NVDLA_cbuf.scala 197:68:@2782.4]
  wire [255:0] _T_87347; // @[Bitwise.scala 72:12:@2784.4]
  wire [255:0] _T_86790_12_0; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4157.4]
  wire [255:0] _T_87348; // @[NV_NVDLA_cbuf.scala 198:65:@2785.4]
  wire [255:0] _T_87353; // @[Bitwise.scala 72:12:@2789.4]
  wire [255:0] _T_86790_13_1; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4184.4]
  wire [255:0] _T_87354; // @[NV_NVDLA_cbuf.scala 197:68:@2790.4]
  wire [255:0] _T_87358; // @[Bitwise.scala 72:12:@2792.4]
  wire [255:0] _T_86790_13_0; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4175.4]
  wire [255:0] _T_87359; // @[NV_NVDLA_cbuf.scala 198:65:@2793.4]
  wire [255:0] _T_87364; // @[Bitwise.scala 72:12:@2797.4]
  wire [255:0] _T_86790_14_1; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4202.4]
  wire [255:0] _T_87365; // @[NV_NVDLA_cbuf.scala 197:68:@2798.4]
  wire [255:0] _T_87369; // @[Bitwise.scala 72:12:@2800.4]
  wire [255:0] _T_86790_14_0; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4193.4]
  wire [255:0] _T_87370; // @[NV_NVDLA_cbuf.scala 198:65:@2801.4]
  wire [255:0] _T_87375; // @[Bitwise.scala 72:12:@2805.4]
  wire [255:0] _T_86790_15_1; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4220.4]
  wire [255:0] _T_87376; // @[NV_NVDLA_cbuf.scala 197:68:@2806.4]
  wire [255:0] _T_87380; // @[Bitwise.scala 72:12:@2808.4]
  wire [255:0] _T_86790_15_0; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4211.4]
  wire [255:0] _T_87381; // @[NV_NVDLA_cbuf.scala 198:65:@2809.4]
  reg [511:0] _T_87674_0_0; // @[NV_NVDLA_cbuf.scala 233:39:@2812.4]
  reg [511:0] _RAND_232;
  reg [511:0] _T_87674_1_0; // @[NV_NVDLA_cbuf.scala 233:39:@2812.4]
  reg [511:0] _RAND_233;
  reg [511:0] _T_87674_2_0; // @[NV_NVDLA_cbuf.scala 233:39:@2812.4]
  reg [511:0] _RAND_234;
  reg [511:0] _T_87674_3_0; // @[NV_NVDLA_cbuf.scala 233:39:@2812.4]
  reg [511:0] _RAND_235;
  reg [511:0] _T_87674_4_0; // @[NV_NVDLA_cbuf.scala 233:39:@2812.4]
  reg [511:0] _RAND_236;
  reg [511:0] _T_87674_5_0; // @[NV_NVDLA_cbuf.scala 233:39:@2812.4]
  reg [511:0] _RAND_237;
  reg [511:0] _T_87674_6_0; // @[NV_NVDLA_cbuf.scala 233:39:@2812.4]
  reg [511:0] _RAND_238;
  reg [511:0] _T_87674_7_0; // @[NV_NVDLA_cbuf.scala 233:39:@2812.4]
  reg [511:0] _RAND_239;
  reg [511:0] _T_87674_8_0; // @[NV_NVDLA_cbuf.scala 233:39:@2812.4]
  reg [511:0] _RAND_240;
  reg [511:0] _T_87674_9_0; // @[NV_NVDLA_cbuf.scala 233:39:@2812.4]
  reg [511:0] _RAND_241;
  reg [511:0] _T_87674_10_0; // @[NV_NVDLA_cbuf.scala 233:39:@2812.4]
  reg [511:0] _RAND_242;
  reg [511:0] _T_87674_11_0; // @[NV_NVDLA_cbuf.scala 233:39:@2812.4]
  reg [511:0] _RAND_243;
  reg [511:0] _T_87674_12_0; // @[NV_NVDLA_cbuf.scala 233:39:@2812.4]
  reg [511:0] _RAND_244;
  reg [511:0] _T_87674_13_0; // @[NV_NVDLA_cbuf.scala 233:39:@2812.4]
  reg [511:0] _RAND_245;
  reg [511:0] _T_87674_14_0; // @[NV_NVDLA_cbuf.scala 233:39:@2812.4]
  reg [511:0] _RAND_246;
  reg [511:0] _T_87674_15_0; // @[NV_NVDLA_cbuf.scala 233:39:@2812.4]
  reg [511:0] _RAND_247;
  reg [511:0] _T_88155_0_0; // @[NV_NVDLA_cbuf.scala 235:35:@2829.4]
  reg [511:0] _RAND_248;
  reg [511:0] _T_88155_1_0; // @[NV_NVDLA_cbuf.scala 235:35:@2829.4]
  reg [511:0] _RAND_249;
  reg [511:0] _T_88155_2_0; // @[NV_NVDLA_cbuf.scala 235:35:@2829.4]
  reg [511:0] _RAND_250;
  reg [511:0] _T_88155_3_0; // @[NV_NVDLA_cbuf.scala 235:35:@2829.4]
  reg [511:0] _RAND_251;
  wire [511:0] _T_88202; // @[NV_NVDLA_cbuf.scala 237:67:@2830.4]
  wire [511:0] _T_88203; // @[NV_NVDLA_cbuf.scala 237:98:@2831.4]
  wire [511:0] _T_88205; // @[NV_NVDLA_cbuf.scala 237:67:@2834.4]
  wire [511:0] _T_88206; // @[NV_NVDLA_cbuf.scala 237:98:@2835.4]
  wire [511:0] _T_88208; // @[NV_NVDLA_cbuf.scala 237:67:@2838.4]
  wire [511:0] _T_88209; // @[NV_NVDLA_cbuf.scala 237:98:@2839.4]
  wire [511:0] _T_88211; // @[NV_NVDLA_cbuf.scala 237:67:@2842.4]
  wire [511:0] _T_88212; // @[NV_NVDLA_cbuf.scala 237:98:@2843.4]
  reg [511:0] _T_88225_0_0; // @[NV_NVDLA_cbuf.scala 240:35:@2846.4]
  reg [511:0] _RAND_252;
  wire [511:0] _T_88245; // @[NV_NVDLA_cbuf.scala 242:67:@2847.4]
  wire [511:0] _T_88246; // @[NV_NVDLA_cbuf.scala 242:98:@2848.4]
  reg [511:0] _T_88249; // @[NV_NVDLA_cbuf.scala 246:35:@2851.4]
  reg [511:0] _RAND_253;
  wire [3:0] _T_88529; // @[NV_NVDLA_cbuf.scala 265:100:@2855.4]
  wire  _T_88531; // @[NV_NVDLA_cbuf.scala 265:151:@2856.4]
  wire  _T_88532; // @[NV_NVDLA_cbuf.scala 265:72:@2857.4]
  wire  _T_88539; // @[NV_NVDLA_cbuf.scala 265:151:@2864.4]
  wire  _T_88540; // @[NV_NVDLA_cbuf.scala 265:72:@2865.4]
  wire  _T_88547; // @[NV_NVDLA_cbuf.scala 265:151:@2872.4]
  wire  _T_88548; // @[NV_NVDLA_cbuf.scala 265:72:@2873.4]
  wire  _T_88555; // @[NV_NVDLA_cbuf.scala 265:151:@2880.4]
  wire  _T_88556; // @[NV_NVDLA_cbuf.scala 265:72:@2881.4]
  wire  _T_88563; // @[NV_NVDLA_cbuf.scala 265:151:@2888.4]
  wire  _T_88564; // @[NV_NVDLA_cbuf.scala 265:72:@2889.4]
  wire  _T_88571; // @[NV_NVDLA_cbuf.scala 265:151:@2896.4]
  wire  _T_88572; // @[NV_NVDLA_cbuf.scala 265:72:@2897.4]
  wire  _T_88579; // @[NV_NVDLA_cbuf.scala 265:151:@2904.4]
  wire  _T_88580; // @[NV_NVDLA_cbuf.scala 265:72:@2905.4]
  wire  _T_88587; // @[NV_NVDLA_cbuf.scala 265:151:@2912.4]
  wire  _T_88588; // @[NV_NVDLA_cbuf.scala 265:72:@2913.4]
  wire  _T_88595; // @[NV_NVDLA_cbuf.scala 265:151:@2920.4]
  wire  _T_88596; // @[NV_NVDLA_cbuf.scala 265:72:@2921.4]
  wire  _T_88603; // @[NV_NVDLA_cbuf.scala 265:151:@2928.4]
  wire  _T_88604; // @[NV_NVDLA_cbuf.scala 265:72:@2929.4]
  wire  _T_88611; // @[NV_NVDLA_cbuf.scala 265:151:@2936.4]
  wire  _T_88612; // @[NV_NVDLA_cbuf.scala 265:72:@2937.4]
  wire  _T_88619; // @[NV_NVDLA_cbuf.scala 265:151:@2944.4]
  wire  _T_88620; // @[NV_NVDLA_cbuf.scala 265:72:@2945.4]
  wire  _T_88627; // @[NV_NVDLA_cbuf.scala 265:151:@2952.4]
  wire  _T_88628; // @[NV_NVDLA_cbuf.scala 265:72:@2953.4]
  wire  _T_88635; // @[NV_NVDLA_cbuf.scala 265:151:@2960.4]
  wire  _T_88636; // @[NV_NVDLA_cbuf.scala 265:72:@2961.4]
  wire  _T_88643; // @[NV_NVDLA_cbuf.scala 265:151:@2968.4]
  wire  _T_88644; // @[NV_NVDLA_cbuf.scala 265:72:@2969.4]
  wire  _T_88651; // @[NV_NVDLA_cbuf.scala 265:151:@2976.4]
  wire  _T_88652; // @[NV_NVDLA_cbuf.scala 265:72:@2977.4]
  wire [8:0] _T_88939; // @[Bitwise.scala 72:12:@2985.4]
  wire [8:0] _T_88940; // @[NV_NVDLA_cbuf.scala 285:128:@2986.4]
  wire [8:0] _T_88941; // @[NV_NVDLA_cbuf.scala 285:101:@2987.4]
  wire [8:0] _T_88951; // @[Bitwise.scala 72:12:@2995.4]
  wire [8:0] _T_88953; // @[NV_NVDLA_cbuf.scala 285:101:@2997.4]
  wire [8:0] _T_88963; // @[Bitwise.scala 72:12:@3005.4]
  wire [8:0] _T_88965; // @[NV_NVDLA_cbuf.scala 285:101:@3007.4]
  wire [8:0] _T_88975; // @[Bitwise.scala 72:12:@3015.4]
  wire [8:0] _T_88977; // @[NV_NVDLA_cbuf.scala 285:101:@3017.4]
  wire [8:0] _T_88987; // @[Bitwise.scala 72:12:@3025.4]
  wire [8:0] _T_88989; // @[NV_NVDLA_cbuf.scala 285:101:@3027.4]
  wire [8:0] _T_88999; // @[Bitwise.scala 72:12:@3035.4]
  wire [8:0] _T_89001; // @[NV_NVDLA_cbuf.scala 285:101:@3037.4]
  wire [8:0] _T_89011; // @[Bitwise.scala 72:12:@3045.4]
  wire [8:0] _T_89013; // @[NV_NVDLA_cbuf.scala 285:101:@3047.4]
  wire [8:0] _T_89023; // @[Bitwise.scala 72:12:@3055.4]
  wire [8:0] _T_89025; // @[NV_NVDLA_cbuf.scala 285:101:@3057.4]
  wire [8:0] _T_89035; // @[Bitwise.scala 72:12:@3065.4]
  wire [8:0] _T_89037; // @[NV_NVDLA_cbuf.scala 285:101:@3067.4]
  wire [8:0] _T_89047; // @[Bitwise.scala 72:12:@3075.4]
  wire [8:0] _T_89049; // @[NV_NVDLA_cbuf.scala 285:101:@3077.4]
  wire [8:0] _T_89059; // @[Bitwise.scala 72:12:@3085.4]
  wire [8:0] _T_89061; // @[NV_NVDLA_cbuf.scala 285:101:@3087.4]
  wire [8:0] _T_89071; // @[Bitwise.scala 72:12:@3095.4]
  wire [8:0] _T_89073; // @[NV_NVDLA_cbuf.scala 285:101:@3097.4]
  wire [8:0] _T_89083; // @[Bitwise.scala 72:12:@3105.4]
  wire [8:0] _T_89085; // @[NV_NVDLA_cbuf.scala 285:101:@3107.4]
  wire [8:0] _T_89095; // @[Bitwise.scala 72:12:@3115.4]
  wire [8:0] _T_89097; // @[NV_NVDLA_cbuf.scala 285:101:@3117.4]
  wire [8:0] _T_89107; // @[Bitwise.scala 72:12:@3125.4]
  wire [8:0] _T_89109; // @[NV_NVDLA_cbuf.scala 285:101:@3127.4]
  wire [8:0] _T_89119; // @[Bitwise.scala 72:12:@3135.4]
  wire [8:0] _T_89121; // @[NV_NVDLA_cbuf.scala 285:101:@3137.4]
  reg  _T_89522_0_0; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_254;
  reg  _T_89522_0_1; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_255;
  reg  _T_89522_1_0; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_256;
  reg  _T_89522_1_1; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_257;
  reg  _T_89522_2_0; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_258;
  reg  _T_89522_2_1; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_259;
  reg  _T_89522_3_0; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_260;
  reg  _T_89522_3_1; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_261;
  reg  _T_89522_4_0; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_262;
  reg  _T_89522_4_1; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_263;
  reg  _T_89522_5_0; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_264;
  reg  _T_89522_5_1; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_265;
  reg  _T_89522_6_0; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_266;
  reg  _T_89522_6_1; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_267;
  reg  _T_89522_7_0; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_268;
  reg  _T_89522_7_1; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_269;
  reg  _T_89522_8_0; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_270;
  reg  _T_89522_8_1; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_271;
  reg  _T_89522_9_0; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_272;
  reg  _T_89522_9_1; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_273;
  reg  _T_89522_10_0; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_274;
  reg  _T_89522_10_1; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_275;
  reg  _T_89522_11_0; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_276;
  reg  _T_89522_11_1; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_277;
  reg  _T_89522_12_0; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_278;
  reg  _T_89522_12_1; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_279;
  reg  _T_89522_13_0; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_280;
  reg  _T_89522_13_1; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_281;
  reg  _T_89522_14_0; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_282;
  reg  _T_89522_14_1; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_283;
  reg  _T_89522_15_0; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_284;
  reg  _T_89522_15_1; // @[Reg.scala 11:16:@3144.4]
  reg [31:0] _RAND_285;
  reg  _T_91073_0_0; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_286;
  reg  _T_91073_0_1; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_287;
  reg  _T_91073_1_0; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_288;
  reg  _T_91073_1_1; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_289;
  reg  _T_91073_2_0; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_290;
  reg  _T_91073_2_1; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_291;
  reg  _T_91073_3_0; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_292;
  reg  _T_91073_3_1; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_293;
  reg  _T_91073_4_0; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_294;
  reg  _T_91073_4_1; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_295;
  reg  _T_91073_5_0; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_296;
  reg  _T_91073_5_1; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_297;
  reg  _T_91073_6_0; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_298;
  reg  _T_91073_6_1; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_299;
  reg  _T_91073_7_0; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_300;
  reg  _T_91073_7_1; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_301;
  reg  _T_91073_8_0; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_302;
  reg  _T_91073_8_1; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_303;
  reg  _T_91073_9_0; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_304;
  reg  _T_91073_9_1; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_305;
  reg  _T_91073_10_0; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_306;
  reg  _T_91073_10_1; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_307;
  reg  _T_91073_11_0; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_308;
  reg  _T_91073_11_1; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_309;
  reg  _T_91073_12_0; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_310;
  reg  _T_91073_12_1; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_311;
  reg  _T_91073_13_0; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_312;
  reg  _T_91073_13_1; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_313;
  reg  _T_91073_14_0; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_314;
  reg  _T_91073_14_1; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_315;
  reg  _T_91073_15_0; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_316;
  reg  _T_91073_15_1; // @[Reg.scala 11:16:@3179.4]
  reg [31:0] _RAND_317;
  wire [7:0] _T_92339; // @[NV_NVDLA_cbuf.scala 298:70:@3220.4]
  wire [15:0] _T_92347; // @[NV_NVDLA_cbuf.scala 298:70:@3228.4]
  wire [7:0] _T_92354; // @[NV_NVDLA_cbuf.scala 298:70:@3235.4]
  wire [31:0] _T_92363; // @[NV_NVDLA_cbuf.scala 298:70:@3244.4]
  reg  _T_92368; // @[Reg.scala 11:16:@3246.4]
  reg [31:0] _RAND_318;
  reg  _T_92370; // @[Reg.scala 11:16:@3250.4]
  reg [31:0] _RAND_319;
  reg  _T_92372; // @[Reg.scala 11:16:@3254.4]
  reg [31:0] _RAND_320;
  reg  _T_92374; // @[Reg.scala 11:16:@3258.4]
  reg [31:0] _RAND_321;
  wire [255:0] _T_92400; // @[Bitwise.scala 72:12:@3265.4]
  wire [255:0] _T_92401; // @[NV_NVDLA_cbuf.scala 315:63:@3266.4]
  wire [255:0] _T_92405; // @[Bitwise.scala 72:12:@3268.4]
  wire [255:0] _T_92406; // @[NV_NVDLA_cbuf.scala 316:61:@3269.4]
  wire [255:0] _T_92411; // @[Bitwise.scala 72:12:@3273.4]
  wire [255:0] _T_92412; // @[NV_NVDLA_cbuf.scala 315:63:@3274.4]
  wire [255:0] _T_92416; // @[Bitwise.scala 72:12:@3276.4]
  wire [255:0] _T_92417; // @[NV_NVDLA_cbuf.scala 316:61:@3277.4]
  wire [255:0] _T_92422; // @[Bitwise.scala 72:12:@3281.4]
  wire [255:0] _T_92423; // @[NV_NVDLA_cbuf.scala 315:63:@3282.4]
  wire [255:0] _T_92427; // @[Bitwise.scala 72:12:@3284.4]
  wire [255:0] _T_92428; // @[NV_NVDLA_cbuf.scala 316:61:@3285.4]
  wire [255:0] _T_92433; // @[Bitwise.scala 72:12:@3289.4]
  wire [255:0] _T_92434; // @[NV_NVDLA_cbuf.scala 315:63:@3290.4]
  wire [255:0] _T_92438; // @[Bitwise.scala 72:12:@3292.4]
  wire [255:0] _T_92439; // @[NV_NVDLA_cbuf.scala 316:61:@3293.4]
  wire [255:0] _T_92444; // @[Bitwise.scala 72:12:@3297.4]
  wire [255:0] _T_92445; // @[NV_NVDLA_cbuf.scala 315:63:@3298.4]
  wire [255:0] _T_92449; // @[Bitwise.scala 72:12:@3300.4]
  wire [255:0] _T_92450; // @[NV_NVDLA_cbuf.scala 316:61:@3301.4]
  wire [255:0] _T_92455; // @[Bitwise.scala 72:12:@3305.4]
  wire [255:0] _T_92456; // @[NV_NVDLA_cbuf.scala 315:63:@3306.4]
  wire [255:0] _T_92460; // @[Bitwise.scala 72:12:@3308.4]
  wire [255:0] _T_92461; // @[NV_NVDLA_cbuf.scala 316:61:@3309.4]
  wire [255:0] _T_92466; // @[Bitwise.scala 72:12:@3313.4]
  wire [255:0] _T_92467; // @[NV_NVDLA_cbuf.scala 315:63:@3314.4]
  wire [255:0] _T_92471; // @[Bitwise.scala 72:12:@3316.4]
  wire [255:0] _T_92472; // @[NV_NVDLA_cbuf.scala 316:61:@3317.4]
  wire [255:0] _T_92477; // @[Bitwise.scala 72:12:@3321.4]
  wire [255:0] _T_92478; // @[NV_NVDLA_cbuf.scala 315:63:@3322.4]
  wire [255:0] _T_92482; // @[Bitwise.scala 72:12:@3324.4]
  wire [255:0] _T_92483; // @[NV_NVDLA_cbuf.scala 316:61:@3325.4]
  wire [255:0] _T_92488; // @[Bitwise.scala 72:12:@3329.4]
  wire [255:0] _T_92489; // @[NV_NVDLA_cbuf.scala 315:63:@3330.4]
  wire [255:0] _T_92493; // @[Bitwise.scala 72:12:@3332.4]
  wire [255:0] _T_92494; // @[NV_NVDLA_cbuf.scala 316:61:@3333.4]
  wire [255:0] _T_92499; // @[Bitwise.scala 72:12:@3337.4]
  wire [255:0] _T_92500; // @[NV_NVDLA_cbuf.scala 315:63:@3338.4]
  wire [255:0] _T_92504; // @[Bitwise.scala 72:12:@3340.4]
  wire [255:0] _T_92505; // @[NV_NVDLA_cbuf.scala 316:61:@3341.4]
  wire [255:0] _T_92510; // @[Bitwise.scala 72:12:@3345.4]
  wire [255:0] _T_92511; // @[NV_NVDLA_cbuf.scala 315:63:@3346.4]
  wire [255:0] _T_92515; // @[Bitwise.scala 72:12:@3348.4]
  wire [255:0] _T_92516; // @[NV_NVDLA_cbuf.scala 316:61:@3349.4]
  wire [255:0] _T_92521; // @[Bitwise.scala 72:12:@3353.4]
  wire [255:0] _T_92522; // @[NV_NVDLA_cbuf.scala 315:63:@3354.4]
  wire [255:0] _T_92526; // @[Bitwise.scala 72:12:@3356.4]
  wire [255:0] _T_92527; // @[NV_NVDLA_cbuf.scala 316:61:@3357.4]
  wire [255:0] _T_92532; // @[Bitwise.scala 72:12:@3361.4]
  wire [255:0] _T_92533; // @[NV_NVDLA_cbuf.scala 315:63:@3362.4]
  wire [255:0] _T_92537; // @[Bitwise.scala 72:12:@3364.4]
  wire [255:0] _T_92538; // @[NV_NVDLA_cbuf.scala 316:61:@3365.4]
  wire [255:0] _T_92543; // @[Bitwise.scala 72:12:@3369.4]
  wire [255:0] _T_92544; // @[NV_NVDLA_cbuf.scala 315:63:@3370.4]
  wire [255:0] _T_92548; // @[Bitwise.scala 72:12:@3372.4]
  wire [255:0] _T_92549; // @[NV_NVDLA_cbuf.scala 316:61:@3373.4]
  wire [255:0] _T_92554; // @[Bitwise.scala 72:12:@3377.4]
  wire [255:0] _T_92555; // @[NV_NVDLA_cbuf.scala 315:63:@3378.4]
  wire [255:0] _T_92559; // @[Bitwise.scala 72:12:@3380.4]
  wire [255:0] _T_92560; // @[NV_NVDLA_cbuf.scala 316:61:@3381.4]
  wire [255:0] _T_92565; // @[Bitwise.scala 72:12:@3385.4]
  wire [255:0] _T_92566; // @[NV_NVDLA_cbuf.scala 315:63:@3386.4]
  wire [255:0] _T_92570; // @[Bitwise.scala 72:12:@3388.4]
  wire [255:0] _T_92571; // @[NV_NVDLA_cbuf.scala 316:61:@3389.4]
  reg [511:0] _T_92609_0; // @[NV_NVDLA_cbuf.scala 350:37:@3392.4]
  reg [511:0] _RAND_322;
  reg [511:0] _T_92609_1; // @[NV_NVDLA_cbuf.scala 350:37:@3392.4]
  reg [511:0] _RAND_323;
  reg [511:0] _T_92609_2; // @[NV_NVDLA_cbuf.scala 350:37:@3392.4]
  reg [511:0] _RAND_324;
  reg [511:0] _T_92609_3; // @[NV_NVDLA_cbuf.scala 350:37:@3392.4]
  reg [511:0] _RAND_325;
  reg [511:0] _T_92609_4; // @[NV_NVDLA_cbuf.scala 350:37:@3392.4]
  reg [511:0] _RAND_326;
  reg [511:0] _T_92609_5; // @[NV_NVDLA_cbuf.scala 350:37:@3392.4]
  reg [511:0] _RAND_327;
  reg [511:0] _T_92609_6; // @[NV_NVDLA_cbuf.scala 350:37:@3392.4]
  reg [511:0] _RAND_328;
  reg [511:0] _T_92609_7; // @[NV_NVDLA_cbuf.scala 350:37:@3392.4]
  reg [511:0] _RAND_329;
  reg [511:0] _T_92609_8; // @[NV_NVDLA_cbuf.scala 350:37:@3392.4]
  reg [511:0] _RAND_330;
  reg [511:0] _T_92609_9; // @[NV_NVDLA_cbuf.scala 350:37:@3392.4]
  reg [511:0] _RAND_331;
  reg [511:0] _T_92609_10; // @[NV_NVDLA_cbuf.scala 350:37:@3392.4]
  reg [511:0] _RAND_332;
  reg [511:0] _T_92609_11; // @[NV_NVDLA_cbuf.scala 350:37:@3392.4]
  reg [511:0] _RAND_333;
  reg [511:0] _T_92609_12; // @[NV_NVDLA_cbuf.scala 350:37:@3392.4]
  reg [511:0] _RAND_334;
  reg [511:0] _T_92609_13; // @[NV_NVDLA_cbuf.scala 350:37:@3392.4]
  reg [511:0] _RAND_335;
  reg [511:0] _T_92609_14; // @[NV_NVDLA_cbuf.scala 350:37:@3392.4]
  reg [511:0] _RAND_336;
  reg [511:0] _T_92609_15; // @[NV_NVDLA_cbuf.scala 350:37:@3392.4]
  reg [511:0] _RAND_337;
  reg [511:0] _T_92665_0; // @[NV_NVDLA_cbuf.scala 352:33:@3409.4]
  reg [511:0] _RAND_338;
  reg [511:0] _T_92665_1; // @[NV_NVDLA_cbuf.scala 352:33:@3409.4]
  reg [511:0] _RAND_339;
  reg [511:0] _T_92665_2; // @[NV_NVDLA_cbuf.scala 352:33:@3409.4]
  reg [511:0] _RAND_340;
  reg [511:0] _T_92665_3; // @[NV_NVDLA_cbuf.scala 352:33:@3409.4]
  reg [511:0] _RAND_341;
  wire [511:0] _T_92672; // @[NV_NVDLA_cbuf.scala 354:57:@3410.4]
  wire [511:0] _T_92673; // @[NV_NVDLA_cbuf.scala 354:83:@3411.4]
  wire [511:0] _T_92675; // @[NV_NVDLA_cbuf.scala 354:57:@3414.4]
  wire [511:0] _T_92676; // @[NV_NVDLA_cbuf.scala 354:83:@3415.4]
  wire [511:0] _T_92678; // @[NV_NVDLA_cbuf.scala 354:57:@3418.4]
  wire [511:0] _T_92679; // @[NV_NVDLA_cbuf.scala 354:83:@3419.4]
  wire [511:0] _T_92681; // @[NV_NVDLA_cbuf.scala 354:57:@3422.4]
  wire [511:0] _T_92682; // @[NV_NVDLA_cbuf.scala 354:83:@3423.4]
  reg [511:0] _T_92687_0; // @[NV_NVDLA_cbuf.scala 357:33:@3426.4]
  reg [511:0] _RAND_342;
  wire [511:0] _T_92691; // @[NV_NVDLA_cbuf.scala 359:57:@3427.4]
  wire [511:0] _T_92692; // @[NV_NVDLA_cbuf.scala 359:83:@3428.4]
  reg [511:0] _T_92695; // @[NV_NVDLA_cbuf.scala 362:33:@3431.4]
  reg [511:0] _RAND_343;
  reg  _T_94145_0_0; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_344;
  reg  _T_94145_0_1; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_345;
  reg  _T_94145_1_0; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_346;
  reg  _T_94145_1_1; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_347;
  reg  _T_94145_2_0; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_348;
  reg  _T_94145_2_1; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_349;
  reg  _T_94145_3_0; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_350;
  reg  _T_94145_3_1; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_351;
  reg  _T_94145_4_0; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_352;
  reg  _T_94145_4_1; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_353;
  reg  _T_94145_5_0; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_354;
  reg  _T_94145_5_1; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_355;
  reg  _T_94145_6_0; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_356;
  reg  _T_94145_6_1; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_357;
  reg  _T_94145_7_0; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_358;
  reg  _T_94145_7_1; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_359;
  reg  _T_94145_8_0; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_360;
  reg  _T_94145_8_1; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_361;
  reg  _T_94145_9_0; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_362;
  reg  _T_94145_9_1; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_363;
  reg  _T_94145_10_0; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_364;
  reg  _T_94145_10_1; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_365;
  reg  _T_94145_11_0; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_366;
  reg  _T_94145_11_1; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_367;
  reg  _T_94145_12_0; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_368;
  reg  _T_94145_12_1; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_369;
  reg  _T_94145_13_0; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_370;
  reg  _T_94145_13_1; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_371;
  reg  _T_94145_14_0; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_372;
  reg  _T_94145_14_1; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_373;
  reg  _T_94145_15_0; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_374;
  reg  _T_94145_15_1; // @[NV_NVDLA_cbuf.scala 377:36:@3515.4]
  reg [31:0] _RAND_375;
  reg [8:0] _T_95257_0_0; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_376;
  reg [8:0] _T_95257_0_1; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_377;
  reg [8:0] _T_95257_1_0; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_378;
  reg [8:0] _T_95257_1_1; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_379;
  reg [8:0] _T_95257_2_0; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_380;
  reg [8:0] _T_95257_2_1; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_381;
  reg [8:0] _T_95257_3_0; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_382;
  reg [8:0] _T_95257_3_1; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_383;
  reg [8:0] _T_95257_4_0; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_384;
  reg [8:0] _T_95257_4_1; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_385;
  reg [8:0] _T_95257_5_0; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_386;
  reg [8:0] _T_95257_5_1; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_387;
  reg [8:0] _T_95257_6_0; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_388;
  reg [8:0] _T_95257_6_1; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_389;
  reg [8:0] _T_95257_7_0; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_390;
  reg [8:0] _T_95257_7_1; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_391;
  reg [8:0] _T_95257_8_0; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_392;
  reg [8:0] _T_95257_8_1; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_393;
  reg [8:0] _T_95257_9_0; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_394;
  reg [8:0] _T_95257_9_1; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_395;
  reg [8:0] _T_95257_10_0; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_396;
  reg [8:0] _T_95257_10_1; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_397;
  reg [8:0] _T_95257_11_0; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_398;
  reg [8:0] _T_95257_11_1; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_399;
  reg [8:0] _T_95257_12_0; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_400;
  reg [8:0] _T_95257_12_1; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_401;
  reg [8:0] _T_95257_13_0; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_402;
  reg [8:0] _T_95257_13_1; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_403;
  reg [8:0] _T_95257_14_0; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_404;
  reg [8:0] _T_95257_14_1; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_405;
  reg [8:0] _T_95257_15_0; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_406;
  reg [8:0] _T_95257_15_1; // @[NV_NVDLA_cbuf.scala 378:34:@3516.4]
  reg [31:0] _RAND_407;
  wire  _T_95463; // @[NV_NVDLA_cbuf.scala 382:68:@3517.4]
  wire [8:0] _T_95468; // @[NV_NVDLA_cbuf.scala 383:103:@3521.4]
  wire [8:0] _T_95473; // @[NV_NVDLA_cbuf.scala 384:98:@3524.4]
  wire  _T_95487; // @[NV_NVDLA_cbuf.scala 382:68:@3537.4]
  wire [8:0] _T_95492; // @[NV_NVDLA_cbuf.scala 383:103:@3541.4]
  wire [8:0] _T_95497; // @[NV_NVDLA_cbuf.scala 384:98:@3544.4]
  wire  _T_95511; // @[NV_NVDLA_cbuf.scala 382:68:@3557.4]
  wire [8:0] _T_95516; // @[NV_NVDLA_cbuf.scala 383:103:@3561.4]
  wire [8:0] _T_95521; // @[NV_NVDLA_cbuf.scala 384:98:@3564.4]
  wire  _T_95535; // @[NV_NVDLA_cbuf.scala 382:68:@3577.4]
  wire [8:0] _T_95540; // @[NV_NVDLA_cbuf.scala 383:103:@3581.4]
  wire [8:0] _T_95545; // @[NV_NVDLA_cbuf.scala 384:98:@3584.4]
  wire  _T_95559; // @[NV_NVDLA_cbuf.scala 382:68:@3597.4]
  wire [8:0] _T_95564; // @[NV_NVDLA_cbuf.scala 383:103:@3601.4]
  wire [8:0] _T_95569; // @[NV_NVDLA_cbuf.scala 384:98:@3604.4]
  wire  _T_95583; // @[NV_NVDLA_cbuf.scala 382:68:@3617.4]
  wire [8:0] _T_95588; // @[NV_NVDLA_cbuf.scala 383:103:@3621.4]
  wire [8:0] _T_95593; // @[NV_NVDLA_cbuf.scala 384:98:@3624.4]
  wire  _T_95607; // @[NV_NVDLA_cbuf.scala 382:68:@3637.4]
  wire [8:0] _T_95612; // @[NV_NVDLA_cbuf.scala 383:103:@3641.4]
  wire [8:0] _T_95617; // @[NV_NVDLA_cbuf.scala 384:98:@3644.4]
  wire  _T_95631; // @[NV_NVDLA_cbuf.scala 382:68:@3657.4]
  wire [8:0] _T_95636; // @[NV_NVDLA_cbuf.scala 383:103:@3661.4]
  wire [8:0] _T_95641; // @[NV_NVDLA_cbuf.scala 384:98:@3664.4]
  wire  _T_95655; // @[NV_NVDLA_cbuf.scala 382:68:@3677.4]
  wire [8:0] _T_95660; // @[NV_NVDLA_cbuf.scala 383:103:@3681.4]
  wire [8:0] _T_95665; // @[NV_NVDLA_cbuf.scala 384:98:@3684.4]
  wire  _T_95679; // @[NV_NVDLA_cbuf.scala 382:68:@3697.4]
  wire [8:0] _T_95684; // @[NV_NVDLA_cbuf.scala 383:103:@3701.4]
  wire [8:0] _T_95689; // @[NV_NVDLA_cbuf.scala 384:98:@3704.4]
  wire  _T_95703; // @[NV_NVDLA_cbuf.scala 382:68:@3717.4]
  wire [8:0] _T_95708; // @[NV_NVDLA_cbuf.scala 383:103:@3721.4]
  wire [8:0] _T_95713; // @[NV_NVDLA_cbuf.scala 384:98:@3724.4]
  wire  _T_95727; // @[NV_NVDLA_cbuf.scala 382:68:@3737.4]
  wire [8:0] _T_95732; // @[NV_NVDLA_cbuf.scala 383:103:@3741.4]
  wire [8:0] _T_95737; // @[NV_NVDLA_cbuf.scala 384:98:@3744.4]
  wire  _T_95751; // @[NV_NVDLA_cbuf.scala 382:68:@3757.4]
  wire [8:0] _T_95756; // @[NV_NVDLA_cbuf.scala 383:103:@3761.4]
  wire [8:0] _T_95761; // @[NV_NVDLA_cbuf.scala 384:98:@3764.4]
  wire  _T_95775; // @[NV_NVDLA_cbuf.scala 382:68:@3777.4]
  wire [8:0] _T_95780; // @[NV_NVDLA_cbuf.scala 383:103:@3781.4]
  wire [8:0] _T_95785; // @[NV_NVDLA_cbuf.scala 384:98:@3784.4]
  wire  _T_95799; // @[NV_NVDLA_cbuf.scala 382:68:@3797.4]
  wire [8:0] _T_95804; // @[NV_NVDLA_cbuf.scala 383:103:@3801.4]
  wire [8:0] _T_95809; // @[NV_NVDLA_cbuf.scala 384:98:@3804.4]
  wire  _T_95823; // @[NV_NVDLA_cbuf.scala 382:68:@3817.4]
  wire [8:0] _T_95828; // @[NV_NVDLA_cbuf.scala 383:103:@3821.4]
  wire [8:0] _T_95833; // @[NV_NVDLA_cbuf.scala 384:98:@3824.4]
  nv_ram_rws nv_ram_rws ( // @[NV_NVDLA_cbuf.scala 389:106:@3837.4]
    .io_clk(nv_ram_rws_io_clk),
    .io_re(nv_ram_rws_io_re),
    .io_we(nv_ram_rws_io_we),
    .io_ra(nv_ram_rws_io_ra),
    .io_wa(nv_ram_rws_io_wa),
    .io_di(nv_ram_rws_io_di),
    .io_dout(nv_ram_rws_io_dout)
  );
  nv_ram_rws nv_ram_rws_1 ( // @[NV_NVDLA_cbuf.scala 389:106:@3840.4]
    .io_clk(nv_ram_rws_1_io_clk),
    .io_re(nv_ram_rws_1_io_re),
    .io_we(nv_ram_rws_1_io_we),
    .io_ra(nv_ram_rws_1_io_ra),
    .io_wa(nv_ram_rws_1_io_wa),
    .io_di(nv_ram_rws_1_io_di),
    .io_dout(nv_ram_rws_1_io_dout)
  );
  nv_ram_rws nv_ram_rws_2 ( // @[NV_NVDLA_cbuf.scala 389:106:@3843.4]
    .io_clk(nv_ram_rws_2_io_clk),
    .io_re(nv_ram_rws_2_io_re),
    .io_we(nv_ram_rws_2_io_we),
    .io_ra(nv_ram_rws_2_io_ra),
    .io_wa(nv_ram_rws_2_io_wa),
    .io_di(nv_ram_rws_2_io_di),
    .io_dout(nv_ram_rws_2_io_dout)
  );
  nv_ram_rws nv_ram_rws_3 ( // @[NV_NVDLA_cbuf.scala 389:106:@3846.4]
    .io_clk(nv_ram_rws_3_io_clk),
    .io_re(nv_ram_rws_3_io_re),
    .io_we(nv_ram_rws_3_io_we),
    .io_ra(nv_ram_rws_3_io_ra),
    .io_wa(nv_ram_rws_3_io_wa),
    .io_di(nv_ram_rws_3_io_di),
    .io_dout(nv_ram_rws_3_io_dout)
  );
  nv_ram_rws nv_ram_rws_4 ( // @[NV_NVDLA_cbuf.scala 389:106:@3849.4]
    .io_clk(nv_ram_rws_4_io_clk),
    .io_re(nv_ram_rws_4_io_re),
    .io_we(nv_ram_rws_4_io_we),
    .io_ra(nv_ram_rws_4_io_ra),
    .io_wa(nv_ram_rws_4_io_wa),
    .io_di(nv_ram_rws_4_io_di),
    .io_dout(nv_ram_rws_4_io_dout)
  );
  nv_ram_rws nv_ram_rws_5 ( // @[NV_NVDLA_cbuf.scala 389:106:@3852.4]
    .io_clk(nv_ram_rws_5_io_clk),
    .io_re(nv_ram_rws_5_io_re),
    .io_we(nv_ram_rws_5_io_we),
    .io_ra(nv_ram_rws_5_io_ra),
    .io_wa(nv_ram_rws_5_io_wa),
    .io_di(nv_ram_rws_5_io_di),
    .io_dout(nv_ram_rws_5_io_dout)
  );
  nv_ram_rws nv_ram_rws_6 ( // @[NV_NVDLA_cbuf.scala 389:106:@3855.4]
    .io_clk(nv_ram_rws_6_io_clk),
    .io_re(nv_ram_rws_6_io_re),
    .io_we(nv_ram_rws_6_io_we),
    .io_ra(nv_ram_rws_6_io_ra),
    .io_wa(nv_ram_rws_6_io_wa),
    .io_di(nv_ram_rws_6_io_di),
    .io_dout(nv_ram_rws_6_io_dout)
  );
  nv_ram_rws nv_ram_rws_7 ( // @[NV_NVDLA_cbuf.scala 389:106:@3858.4]
    .io_clk(nv_ram_rws_7_io_clk),
    .io_re(nv_ram_rws_7_io_re),
    .io_we(nv_ram_rws_7_io_we),
    .io_ra(nv_ram_rws_7_io_ra),
    .io_wa(nv_ram_rws_7_io_wa),
    .io_di(nv_ram_rws_7_io_di),
    .io_dout(nv_ram_rws_7_io_dout)
  );
  nv_ram_rws nv_ram_rws_8 ( // @[NV_NVDLA_cbuf.scala 389:106:@3861.4]
    .io_clk(nv_ram_rws_8_io_clk),
    .io_re(nv_ram_rws_8_io_re),
    .io_we(nv_ram_rws_8_io_we),
    .io_ra(nv_ram_rws_8_io_ra),
    .io_wa(nv_ram_rws_8_io_wa),
    .io_di(nv_ram_rws_8_io_di),
    .io_dout(nv_ram_rws_8_io_dout)
  );
  nv_ram_rws nv_ram_rws_9 ( // @[NV_NVDLA_cbuf.scala 389:106:@3864.4]
    .io_clk(nv_ram_rws_9_io_clk),
    .io_re(nv_ram_rws_9_io_re),
    .io_we(nv_ram_rws_9_io_we),
    .io_ra(nv_ram_rws_9_io_ra),
    .io_wa(nv_ram_rws_9_io_wa),
    .io_di(nv_ram_rws_9_io_di),
    .io_dout(nv_ram_rws_9_io_dout)
  );
  nv_ram_rws nv_ram_rws_10 ( // @[NV_NVDLA_cbuf.scala 389:106:@3867.4]
    .io_clk(nv_ram_rws_10_io_clk),
    .io_re(nv_ram_rws_10_io_re),
    .io_we(nv_ram_rws_10_io_we),
    .io_ra(nv_ram_rws_10_io_ra),
    .io_wa(nv_ram_rws_10_io_wa),
    .io_di(nv_ram_rws_10_io_di),
    .io_dout(nv_ram_rws_10_io_dout)
  );
  nv_ram_rws nv_ram_rws_11 ( // @[NV_NVDLA_cbuf.scala 389:106:@3870.4]
    .io_clk(nv_ram_rws_11_io_clk),
    .io_re(nv_ram_rws_11_io_re),
    .io_we(nv_ram_rws_11_io_we),
    .io_ra(nv_ram_rws_11_io_ra),
    .io_wa(nv_ram_rws_11_io_wa),
    .io_di(nv_ram_rws_11_io_di),
    .io_dout(nv_ram_rws_11_io_dout)
  );
  nv_ram_rws nv_ram_rws_12 ( // @[NV_NVDLA_cbuf.scala 389:106:@3873.4]
    .io_clk(nv_ram_rws_12_io_clk),
    .io_re(nv_ram_rws_12_io_re),
    .io_we(nv_ram_rws_12_io_we),
    .io_ra(nv_ram_rws_12_io_ra),
    .io_wa(nv_ram_rws_12_io_wa),
    .io_di(nv_ram_rws_12_io_di),
    .io_dout(nv_ram_rws_12_io_dout)
  );
  nv_ram_rws nv_ram_rws_13 ( // @[NV_NVDLA_cbuf.scala 389:106:@3876.4]
    .io_clk(nv_ram_rws_13_io_clk),
    .io_re(nv_ram_rws_13_io_re),
    .io_we(nv_ram_rws_13_io_we),
    .io_ra(nv_ram_rws_13_io_ra),
    .io_wa(nv_ram_rws_13_io_wa),
    .io_di(nv_ram_rws_13_io_di),
    .io_dout(nv_ram_rws_13_io_dout)
  );
  nv_ram_rws nv_ram_rws_14 ( // @[NV_NVDLA_cbuf.scala 389:106:@3879.4]
    .io_clk(nv_ram_rws_14_io_clk),
    .io_re(nv_ram_rws_14_io_re),
    .io_we(nv_ram_rws_14_io_we),
    .io_ra(nv_ram_rws_14_io_ra),
    .io_wa(nv_ram_rws_14_io_wa),
    .io_di(nv_ram_rws_14_io_di),
    .io_dout(nv_ram_rws_14_io_dout)
  );
  nv_ram_rws nv_ram_rws_15 ( // @[NV_NVDLA_cbuf.scala 389:106:@3882.4]
    .io_clk(nv_ram_rws_15_io_clk),
    .io_re(nv_ram_rws_15_io_re),
    .io_we(nv_ram_rws_15_io_we),
    .io_ra(nv_ram_rws_15_io_ra),
    .io_wa(nv_ram_rws_15_io_wa),
    .io_di(nv_ram_rws_15_io_di),
    .io_dout(nv_ram_rws_15_io_dout)
  );
  nv_ram_rws nv_ram_rws_16 ( // @[NV_NVDLA_cbuf.scala 389:106:@3885.4]
    .io_clk(nv_ram_rws_16_io_clk),
    .io_re(nv_ram_rws_16_io_re),
    .io_we(nv_ram_rws_16_io_we),
    .io_ra(nv_ram_rws_16_io_ra),
    .io_wa(nv_ram_rws_16_io_wa),
    .io_di(nv_ram_rws_16_io_di),
    .io_dout(nv_ram_rws_16_io_dout)
  );
  nv_ram_rws nv_ram_rws_17 ( // @[NV_NVDLA_cbuf.scala 389:106:@3888.4]
    .io_clk(nv_ram_rws_17_io_clk),
    .io_re(nv_ram_rws_17_io_re),
    .io_we(nv_ram_rws_17_io_we),
    .io_ra(nv_ram_rws_17_io_ra),
    .io_wa(nv_ram_rws_17_io_wa),
    .io_di(nv_ram_rws_17_io_di),
    .io_dout(nv_ram_rws_17_io_dout)
  );
  nv_ram_rws nv_ram_rws_18 ( // @[NV_NVDLA_cbuf.scala 389:106:@3891.4]
    .io_clk(nv_ram_rws_18_io_clk),
    .io_re(nv_ram_rws_18_io_re),
    .io_we(nv_ram_rws_18_io_we),
    .io_ra(nv_ram_rws_18_io_ra),
    .io_wa(nv_ram_rws_18_io_wa),
    .io_di(nv_ram_rws_18_io_di),
    .io_dout(nv_ram_rws_18_io_dout)
  );
  nv_ram_rws nv_ram_rws_19 ( // @[NV_NVDLA_cbuf.scala 389:106:@3894.4]
    .io_clk(nv_ram_rws_19_io_clk),
    .io_re(nv_ram_rws_19_io_re),
    .io_we(nv_ram_rws_19_io_we),
    .io_ra(nv_ram_rws_19_io_ra),
    .io_wa(nv_ram_rws_19_io_wa),
    .io_di(nv_ram_rws_19_io_di),
    .io_dout(nv_ram_rws_19_io_dout)
  );
  nv_ram_rws nv_ram_rws_20 ( // @[NV_NVDLA_cbuf.scala 389:106:@3897.4]
    .io_clk(nv_ram_rws_20_io_clk),
    .io_re(nv_ram_rws_20_io_re),
    .io_we(nv_ram_rws_20_io_we),
    .io_ra(nv_ram_rws_20_io_ra),
    .io_wa(nv_ram_rws_20_io_wa),
    .io_di(nv_ram_rws_20_io_di),
    .io_dout(nv_ram_rws_20_io_dout)
  );
  nv_ram_rws nv_ram_rws_21 ( // @[NV_NVDLA_cbuf.scala 389:106:@3900.4]
    .io_clk(nv_ram_rws_21_io_clk),
    .io_re(nv_ram_rws_21_io_re),
    .io_we(nv_ram_rws_21_io_we),
    .io_ra(nv_ram_rws_21_io_ra),
    .io_wa(nv_ram_rws_21_io_wa),
    .io_di(nv_ram_rws_21_io_di),
    .io_dout(nv_ram_rws_21_io_dout)
  );
  nv_ram_rws nv_ram_rws_22 ( // @[NV_NVDLA_cbuf.scala 389:106:@3903.4]
    .io_clk(nv_ram_rws_22_io_clk),
    .io_re(nv_ram_rws_22_io_re),
    .io_we(nv_ram_rws_22_io_we),
    .io_ra(nv_ram_rws_22_io_ra),
    .io_wa(nv_ram_rws_22_io_wa),
    .io_di(nv_ram_rws_22_io_di),
    .io_dout(nv_ram_rws_22_io_dout)
  );
  nv_ram_rws nv_ram_rws_23 ( // @[NV_NVDLA_cbuf.scala 389:106:@3906.4]
    .io_clk(nv_ram_rws_23_io_clk),
    .io_re(nv_ram_rws_23_io_re),
    .io_we(nv_ram_rws_23_io_we),
    .io_ra(nv_ram_rws_23_io_ra),
    .io_wa(nv_ram_rws_23_io_wa),
    .io_di(nv_ram_rws_23_io_di),
    .io_dout(nv_ram_rws_23_io_dout)
  );
  nv_ram_rws nv_ram_rws_24 ( // @[NV_NVDLA_cbuf.scala 389:106:@3909.4]
    .io_clk(nv_ram_rws_24_io_clk),
    .io_re(nv_ram_rws_24_io_re),
    .io_we(nv_ram_rws_24_io_we),
    .io_ra(nv_ram_rws_24_io_ra),
    .io_wa(nv_ram_rws_24_io_wa),
    .io_di(nv_ram_rws_24_io_di),
    .io_dout(nv_ram_rws_24_io_dout)
  );
  nv_ram_rws nv_ram_rws_25 ( // @[NV_NVDLA_cbuf.scala 389:106:@3912.4]
    .io_clk(nv_ram_rws_25_io_clk),
    .io_re(nv_ram_rws_25_io_re),
    .io_we(nv_ram_rws_25_io_we),
    .io_ra(nv_ram_rws_25_io_ra),
    .io_wa(nv_ram_rws_25_io_wa),
    .io_di(nv_ram_rws_25_io_di),
    .io_dout(nv_ram_rws_25_io_dout)
  );
  nv_ram_rws nv_ram_rws_26 ( // @[NV_NVDLA_cbuf.scala 389:106:@3915.4]
    .io_clk(nv_ram_rws_26_io_clk),
    .io_re(nv_ram_rws_26_io_re),
    .io_we(nv_ram_rws_26_io_we),
    .io_ra(nv_ram_rws_26_io_ra),
    .io_wa(nv_ram_rws_26_io_wa),
    .io_di(nv_ram_rws_26_io_di),
    .io_dout(nv_ram_rws_26_io_dout)
  );
  nv_ram_rws nv_ram_rws_27 ( // @[NV_NVDLA_cbuf.scala 389:106:@3918.4]
    .io_clk(nv_ram_rws_27_io_clk),
    .io_re(nv_ram_rws_27_io_re),
    .io_we(nv_ram_rws_27_io_we),
    .io_ra(nv_ram_rws_27_io_ra),
    .io_wa(nv_ram_rws_27_io_wa),
    .io_di(nv_ram_rws_27_io_di),
    .io_dout(nv_ram_rws_27_io_dout)
  );
  nv_ram_rws nv_ram_rws_28 ( // @[NV_NVDLA_cbuf.scala 389:106:@3921.4]
    .io_clk(nv_ram_rws_28_io_clk),
    .io_re(nv_ram_rws_28_io_re),
    .io_we(nv_ram_rws_28_io_we),
    .io_ra(nv_ram_rws_28_io_ra),
    .io_wa(nv_ram_rws_28_io_wa),
    .io_di(nv_ram_rws_28_io_di),
    .io_dout(nv_ram_rws_28_io_dout)
  );
  nv_ram_rws nv_ram_rws_29 ( // @[NV_NVDLA_cbuf.scala 389:106:@3924.4]
    .io_clk(nv_ram_rws_29_io_clk),
    .io_re(nv_ram_rws_29_io_re),
    .io_we(nv_ram_rws_29_io_we),
    .io_ra(nv_ram_rws_29_io_ra),
    .io_wa(nv_ram_rws_29_io_wa),
    .io_di(nv_ram_rws_29_io_di),
    .io_dout(nv_ram_rws_29_io_dout)
  );
  nv_ram_rws nv_ram_rws_30 ( // @[NV_NVDLA_cbuf.scala 389:106:@3927.4]
    .io_clk(nv_ram_rws_30_io_clk),
    .io_re(nv_ram_rws_30_io_re),
    .io_we(nv_ram_rws_30_io_we),
    .io_ra(nv_ram_rws_30_io_ra),
    .io_wa(nv_ram_rws_30_io_wa),
    .io_di(nv_ram_rws_30_io_di),
    .io_dout(nv_ram_rws_30_io_dout)
  );
  nv_ram_rws nv_ram_rws_31 ( // @[NV_NVDLA_cbuf.scala 389:106:@3930.4]
    .io_clk(nv_ram_rws_31_io_clk),
    .io_re(nv_ram_rws_31_io_re),
    .io_we(nv_ram_rws_31_io_we),
    .io_ra(nv_ram_rws_31_io_ra),
    .io_wa(nv_ram_rws_31_io_wa),
    .io_di(nv_ram_rws_31_io_di),
    .io_dout(nv_ram_rws_31_io_dout)
  );
  assign _T_178 = io_nvdla_core_rstn == 1'h0; // @[NV_NVDLA_cbuf.scala 26:38:@488.4]
  assign _T_2665 = io_cdma2buf_wr_addr_0[12:9]; // @[NV_NVDLA_cbuf.scala 35:72:@490.4]
  assign _T_2667 = _T_2665 == 4'h0; // @[NV_NVDLA_cbuf.scala 35:123:@491.4]
  assign _T_2668 = io_cdma2buf_wr_en_0 & _T_2667; // @[NV_NVDLA_cbuf.scala 34:69:@492.4]
  assign _T_2669 = io_cdma2buf_wr_sel_0[0]; // @[NV_NVDLA_cbuf.scala 36:71:@493.4]
  assign _T_2672 = _T_2668 & _T_2669; // @[NV_NVDLA_cbuf.scala 35:130:@495.4]
  assign _T_2673 = io_cdma2buf_wr_addr_1[12:9]; // @[NV_NVDLA_cbuf.scala 35:72:@497.4]
  assign _T_2675 = _T_2673 == 4'h0; // @[NV_NVDLA_cbuf.scala 35:123:@498.4]
  assign _T_2676 = io_cdma2buf_wr_en_1 & _T_2675; // @[NV_NVDLA_cbuf.scala 34:69:@499.4]
  assign _T_2677 = io_cdma2buf_wr_sel_1[0]; // @[NV_NVDLA_cbuf.scala 36:71:@500.4]
  assign _T_2680 = _T_2676 & _T_2677; // @[NV_NVDLA_cbuf.scala 35:130:@502.4]
  assign _T_2685 = io_cdma2buf_wr_sel_0[1]; // @[NV_NVDLA_cbuf.scala 36:71:@507.4]
  assign _T_2688 = _T_2668 & _T_2685; // @[NV_NVDLA_cbuf.scala 35:130:@509.4]
  assign _T_2693 = io_cdma2buf_wr_sel_1[1]; // @[NV_NVDLA_cbuf.scala 36:71:@514.4]
  assign _T_2696 = _T_2676 & _T_2693; // @[NV_NVDLA_cbuf.scala 35:130:@516.4]
  assign _T_2699 = _T_2665 == 4'h1; // @[NV_NVDLA_cbuf.scala 35:123:@519.4]
  assign _T_2700 = io_cdma2buf_wr_en_0 & _T_2699; // @[NV_NVDLA_cbuf.scala 34:69:@520.4]
  assign _T_2704 = _T_2700 & _T_2669; // @[NV_NVDLA_cbuf.scala 35:130:@523.4]
  assign _T_2707 = _T_2673 == 4'h1; // @[NV_NVDLA_cbuf.scala 35:123:@526.4]
  assign _T_2708 = io_cdma2buf_wr_en_1 & _T_2707; // @[NV_NVDLA_cbuf.scala 34:69:@527.4]
  assign _T_2712 = _T_2708 & _T_2677; // @[NV_NVDLA_cbuf.scala 35:130:@530.4]
  assign _T_2720 = _T_2700 & _T_2685; // @[NV_NVDLA_cbuf.scala 35:130:@537.4]
  assign _T_2728 = _T_2708 & _T_2693; // @[NV_NVDLA_cbuf.scala 35:130:@544.4]
  assign _T_2731 = _T_2665 == 4'h2; // @[NV_NVDLA_cbuf.scala 35:123:@547.4]
  assign _T_2732 = io_cdma2buf_wr_en_0 & _T_2731; // @[NV_NVDLA_cbuf.scala 34:69:@548.4]
  assign _T_2736 = _T_2732 & _T_2669; // @[NV_NVDLA_cbuf.scala 35:130:@551.4]
  assign _T_2739 = _T_2673 == 4'h2; // @[NV_NVDLA_cbuf.scala 35:123:@554.4]
  assign _T_2740 = io_cdma2buf_wr_en_1 & _T_2739; // @[NV_NVDLA_cbuf.scala 34:69:@555.4]
  assign _T_2744 = _T_2740 & _T_2677; // @[NV_NVDLA_cbuf.scala 35:130:@558.4]
  assign _T_2752 = _T_2732 & _T_2685; // @[NV_NVDLA_cbuf.scala 35:130:@565.4]
  assign _T_2760 = _T_2740 & _T_2693; // @[NV_NVDLA_cbuf.scala 35:130:@572.4]
  assign _T_2763 = _T_2665 == 4'h3; // @[NV_NVDLA_cbuf.scala 35:123:@575.4]
  assign _T_2764 = io_cdma2buf_wr_en_0 & _T_2763; // @[NV_NVDLA_cbuf.scala 34:69:@576.4]
  assign _T_2768 = _T_2764 & _T_2669; // @[NV_NVDLA_cbuf.scala 35:130:@579.4]
  assign _T_2771 = _T_2673 == 4'h3; // @[NV_NVDLA_cbuf.scala 35:123:@582.4]
  assign _T_2772 = io_cdma2buf_wr_en_1 & _T_2771; // @[NV_NVDLA_cbuf.scala 34:69:@583.4]
  assign _T_2776 = _T_2772 & _T_2677; // @[NV_NVDLA_cbuf.scala 35:130:@586.4]
  assign _T_2784 = _T_2764 & _T_2685; // @[NV_NVDLA_cbuf.scala 35:130:@593.4]
  assign _T_2792 = _T_2772 & _T_2693; // @[NV_NVDLA_cbuf.scala 35:130:@600.4]
  assign _T_2795 = _T_2665 == 4'h4; // @[NV_NVDLA_cbuf.scala 35:123:@603.4]
  assign _T_2796 = io_cdma2buf_wr_en_0 & _T_2795; // @[NV_NVDLA_cbuf.scala 34:69:@604.4]
  assign _T_2800 = _T_2796 & _T_2669; // @[NV_NVDLA_cbuf.scala 35:130:@607.4]
  assign _T_2803 = _T_2673 == 4'h4; // @[NV_NVDLA_cbuf.scala 35:123:@610.4]
  assign _T_2804 = io_cdma2buf_wr_en_1 & _T_2803; // @[NV_NVDLA_cbuf.scala 34:69:@611.4]
  assign _T_2808 = _T_2804 & _T_2677; // @[NV_NVDLA_cbuf.scala 35:130:@614.4]
  assign _T_2816 = _T_2796 & _T_2685; // @[NV_NVDLA_cbuf.scala 35:130:@621.4]
  assign _T_2824 = _T_2804 & _T_2693; // @[NV_NVDLA_cbuf.scala 35:130:@628.4]
  assign _T_2827 = _T_2665 == 4'h5; // @[NV_NVDLA_cbuf.scala 35:123:@631.4]
  assign _T_2828 = io_cdma2buf_wr_en_0 & _T_2827; // @[NV_NVDLA_cbuf.scala 34:69:@632.4]
  assign _T_2832 = _T_2828 & _T_2669; // @[NV_NVDLA_cbuf.scala 35:130:@635.4]
  assign _T_2835 = _T_2673 == 4'h5; // @[NV_NVDLA_cbuf.scala 35:123:@638.4]
  assign _T_2836 = io_cdma2buf_wr_en_1 & _T_2835; // @[NV_NVDLA_cbuf.scala 34:69:@639.4]
  assign _T_2840 = _T_2836 & _T_2677; // @[NV_NVDLA_cbuf.scala 35:130:@642.4]
  assign _T_2848 = _T_2828 & _T_2685; // @[NV_NVDLA_cbuf.scala 35:130:@649.4]
  assign _T_2856 = _T_2836 & _T_2693; // @[NV_NVDLA_cbuf.scala 35:130:@656.4]
  assign _T_2859 = _T_2665 == 4'h6; // @[NV_NVDLA_cbuf.scala 35:123:@659.4]
  assign _T_2860 = io_cdma2buf_wr_en_0 & _T_2859; // @[NV_NVDLA_cbuf.scala 34:69:@660.4]
  assign _T_2864 = _T_2860 & _T_2669; // @[NV_NVDLA_cbuf.scala 35:130:@663.4]
  assign _T_2867 = _T_2673 == 4'h6; // @[NV_NVDLA_cbuf.scala 35:123:@666.4]
  assign _T_2868 = io_cdma2buf_wr_en_1 & _T_2867; // @[NV_NVDLA_cbuf.scala 34:69:@667.4]
  assign _T_2872 = _T_2868 & _T_2677; // @[NV_NVDLA_cbuf.scala 35:130:@670.4]
  assign _T_2880 = _T_2860 & _T_2685; // @[NV_NVDLA_cbuf.scala 35:130:@677.4]
  assign _T_2888 = _T_2868 & _T_2693; // @[NV_NVDLA_cbuf.scala 35:130:@684.4]
  assign _T_2891 = _T_2665 == 4'h7; // @[NV_NVDLA_cbuf.scala 35:123:@687.4]
  assign _T_2892 = io_cdma2buf_wr_en_0 & _T_2891; // @[NV_NVDLA_cbuf.scala 34:69:@688.4]
  assign _T_2896 = _T_2892 & _T_2669; // @[NV_NVDLA_cbuf.scala 35:130:@691.4]
  assign _T_2899 = _T_2673 == 4'h7; // @[NV_NVDLA_cbuf.scala 35:123:@694.4]
  assign _T_2900 = io_cdma2buf_wr_en_1 & _T_2899; // @[NV_NVDLA_cbuf.scala 34:69:@695.4]
  assign _T_2904 = _T_2900 & _T_2677; // @[NV_NVDLA_cbuf.scala 35:130:@698.4]
  assign _T_2912 = _T_2892 & _T_2685; // @[NV_NVDLA_cbuf.scala 35:130:@705.4]
  assign _T_2920 = _T_2900 & _T_2693; // @[NV_NVDLA_cbuf.scala 35:130:@712.4]
  assign _T_2923 = _T_2665 == 4'h8; // @[NV_NVDLA_cbuf.scala 35:123:@715.4]
  assign _T_2924 = io_cdma2buf_wr_en_0 & _T_2923; // @[NV_NVDLA_cbuf.scala 34:69:@716.4]
  assign _T_2928 = _T_2924 & _T_2669; // @[NV_NVDLA_cbuf.scala 35:130:@719.4]
  assign _T_2931 = _T_2673 == 4'h8; // @[NV_NVDLA_cbuf.scala 35:123:@722.4]
  assign _T_2932 = io_cdma2buf_wr_en_1 & _T_2931; // @[NV_NVDLA_cbuf.scala 34:69:@723.4]
  assign _T_2936 = _T_2932 & _T_2677; // @[NV_NVDLA_cbuf.scala 35:130:@726.4]
  assign _T_2944 = _T_2924 & _T_2685; // @[NV_NVDLA_cbuf.scala 35:130:@733.4]
  assign _T_2952 = _T_2932 & _T_2693; // @[NV_NVDLA_cbuf.scala 35:130:@740.4]
  assign _T_2955 = _T_2665 == 4'h9; // @[NV_NVDLA_cbuf.scala 35:123:@743.4]
  assign _T_2956 = io_cdma2buf_wr_en_0 & _T_2955; // @[NV_NVDLA_cbuf.scala 34:69:@744.4]
  assign _T_2960 = _T_2956 & _T_2669; // @[NV_NVDLA_cbuf.scala 35:130:@747.4]
  assign _T_2963 = _T_2673 == 4'h9; // @[NV_NVDLA_cbuf.scala 35:123:@750.4]
  assign _T_2964 = io_cdma2buf_wr_en_1 & _T_2963; // @[NV_NVDLA_cbuf.scala 34:69:@751.4]
  assign _T_2968 = _T_2964 & _T_2677; // @[NV_NVDLA_cbuf.scala 35:130:@754.4]
  assign _T_2976 = _T_2956 & _T_2685; // @[NV_NVDLA_cbuf.scala 35:130:@761.4]
  assign _T_2984 = _T_2964 & _T_2693; // @[NV_NVDLA_cbuf.scala 35:130:@768.4]
  assign _T_2987 = _T_2665 == 4'ha; // @[NV_NVDLA_cbuf.scala 35:123:@771.4]
  assign _T_2988 = io_cdma2buf_wr_en_0 & _T_2987; // @[NV_NVDLA_cbuf.scala 34:69:@772.4]
  assign _T_2992 = _T_2988 & _T_2669; // @[NV_NVDLA_cbuf.scala 35:130:@775.4]
  assign _T_2995 = _T_2673 == 4'ha; // @[NV_NVDLA_cbuf.scala 35:123:@778.4]
  assign _T_2996 = io_cdma2buf_wr_en_1 & _T_2995; // @[NV_NVDLA_cbuf.scala 34:69:@779.4]
  assign _T_3000 = _T_2996 & _T_2677; // @[NV_NVDLA_cbuf.scala 35:130:@782.4]
  assign _T_3008 = _T_2988 & _T_2685; // @[NV_NVDLA_cbuf.scala 35:130:@789.4]
  assign _T_3016 = _T_2996 & _T_2693; // @[NV_NVDLA_cbuf.scala 35:130:@796.4]
  assign _T_3019 = _T_2665 == 4'hb; // @[NV_NVDLA_cbuf.scala 35:123:@799.4]
  assign _T_3020 = io_cdma2buf_wr_en_0 & _T_3019; // @[NV_NVDLA_cbuf.scala 34:69:@800.4]
  assign _T_3024 = _T_3020 & _T_2669; // @[NV_NVDLA_cbuf.scala 35:130:@803.4]
  assign _T_3027 = _T_2673 == 4'hb; // @[NV_NVDLA_cbuf.scala 35:123:@806.4]
  assign _T_3028 = io_cdma2buf_wr_en_1 & _T_3027; // @[NV_NVDLA_cbuf.scala 34:69:@807.4]
  assign _T_3032 = _T_3028 & _T_2677; // @[NV_NVDLA_cbuf.scala 35:130:@810.4]
  assign _T_3040 = _T_3020 & _T_2685; // @[NV_NVDLA_cbuf.scala 35:130:@817.4]
  assign _T_3048 = _T_3028 & _T_2693; // @[NV_NVDLA_cbuf.scala 35:130:@824.4]
  assign _T_3051 = _T_2665 == 4'hc; // @[NV_NVDLA_cbuf.scala 35:123:@827.4]
  assign _T_3052 = io_cdma2buf_wr_en_0 & _T_3051; // @[NV_NVDLA_cbuf.scala 34:69:@828.4]
  assign _T_3056 = _T_3052 & _T_2669; // @[NV_NVDLA_cbuf.scala 35:130:@831.4]
  assign _T_3059 = _T_2673 == 4'hc; // @[NV_NVDLA_cbuf.scala 35:123:@834.4]
  assign _T_3060 = io_cdma2buf_wr_en_1 & _T_3059; // @[NV_NVDLA_cbuf.scala 34:69:@835.4]
  assign _T_3064 = _T_3060 & _T_2677; // @[NV_NVDLA_cbuf.scala 35:130:@838.4]
  assign _T_3072 = _T_3052 & _T_2685; // @[NV_NVDLA_cbuf.scala 35:130:@845.4]
  assign _T_3080 = _T_3060 & _T_2693; // @[NV_NVDLA_cbuf.scala 35:130:@852.4]
  assign _T_3083 = _T_2665 == 4'hd; // @[NV_NVDLA_cbuf.scala 35:123:@855.4]
  assign _T_3084 = io_cdma2buf_wr_en_0 & _T_3083; // @[NV_NVDLA_cbuf.scala 34:69:@856.4]
  assign _T_3088 = _T_3084 & _T_2669; // @[NV_NVDLA_cbuf.scala 35:130:@859.4]
  assign _T_3091 = _T_2673 == 4'hd; // @[NV_NVDLA_cbuf.scala 35:123:@862.4]
  assign _T_3092 = io_cdma2buf_wr_en_1 & _T_3091; // @[NV_NVDLA_cbuf.scala 34:69:@863.4]
  assign _T_3096 = _T_3092 & _T_2677; // @[NV_NVDLA_cbuf.scala 35:130:@866.4]
  assign _T_3104 = _T_3084 & _T_2685; // @[NV_NVDLA_cbuf.scala 35:130:@873.4]
  assign _T_3112 = _T_3092 & _T_2693; // @[NV_NVDLA_cbuf.scala 35:130:@880.4]
  assign _T_3115 = _T_2665 == 4'he; // @[NV_NVDLA_cbuf.scala 35:123:@883.4]
  assign _T_3116 = io_cdma2buf_wr_en_0 & _T_3115; // @[NV_NVDLA_cbuf.scala 34:69:@884.4]
  assign _T_3120 = _T_3116 & _T_2669; // @[NV_NVDLA_cbuf.scala 35:130:@887.4]
  assign _T_3123 = _T_2673 == 4'he; // @[NV_NVDLA_cbuf.scala 35:123:@890.4]
  assign _T_3124 = io_cdma2buf_wr_en_1 & _T_3123; // @[NV_NVDLA_cbuf.scala 34:69:@891.4]
  assign _T_3128 = _T_3124 & _T_2677; // @[NV_NVDLA_cbuf.scala 35:130:@894.4]
  assign _T_3136 = _T_3116 & _T_2685; // @[NV_NVDLA_cbuf.scala 35:130:@901.4]
  assign _T_3144 = _T_3124 & _T_2693; // @[NV_NVDLA_cbuf.scala 35:130:@908.4]
  assign _T_3147 = _T_2665 == 4'hf; // @[NV_NVDLA_cbuf.scala 35:123:@911.4]
  assign _T_3148 = io_cdma2buf_wr_en_0 & _T_3147; // @[NV_NVDLA_cbuf.scala 34:69:@912.4]
  assign _T_3152 = _T_3148 & _T_2669; // @[NV_NVDLA_cbuf.scala 35:130:@915.4]
  assign _T_3155 = _T_2673 == 4'hf; // @[NV_NVDLA_cbuf.scala 35:123:@918.4]
  assign _T_3156 = io_cdma2buf_wr_en_1 & _T_3155; // @[NV_NVDLA_cbuf.scala 34:69:@919.4]
  assign _T_3160 = _T_3156 & _T_2677; // @[NV_NVDLA_cbuf.scala 35:130:@922.4]
  assign _T_3168 = _T_3148 & _T_2685; // @[NV_NVDLA_cbuf.scala 35:130:@929.4]
  assign _T_3176 = _T_3156 & _T_2693; // @[NV_NVDLA_cbuf.scala 35:130:@936.4]
  assign _T_8151 = _T_2672 | _T_2680; // @[NV_NVDLA_cbuf.scala 74:72:@1085.4]
  assign _T_8152 = _T_2688 | _T_2696; // @[NV_NVDLA_cbuf.scala 74:72:@1087.4]
  assign _T_8153 = _T_2704 | _T_2712; // @[NV_NVDLA_cbuf.scala 74:72:@1089.4]
  assign _T_8154 = _T_2720 | _T_2728; // @[NV_NVDLA_cbuf.scala 74:72:@1091.4]
  assign _T_8155 = _T_2736 | _T_2744; // @[NV_NVDLA_cbuf.scala 74:72:@1093.4]
  assign _T_8156 = _T_2752 | _T_2760; // @[NV_NVDLA_cbuf.scala 74:72:@1095.4]
  assign _T_8157 = _T_2768 | _T_2776; // @[NV_NVDLA_cbuf.scala 74:72:@1097.4]
  assign _T_8158 = _T_2784 | _T_2792; // @[NV_NVDLA_cbuf.scala 74:72:@1099.4]
  assign _T_8159 = _T_2800 | _T_2808; // @[NV_NVDLA_cbuf.scala 74:72:@1101.4]
  assign _T_8160 = _T_2816 | _T_2824; // @[NV_NVDLA_cbuf.scala 74:72:@1103.4]
  assign _T_8161 = _T_2832 | _T_2840; // @[NV_NVDLA_cbuf.scala 74:72:@1105.4]
  assign _T_8162 = _T_2848 | _T_2856; // @[NV_NVDLA_cbuf.scala 74:72:@1107.4]
  assign _T_8163 = _T_2864 | _T_2872; // @[NV_NVDLA_cbuf.scala 74:72:@1109.4]
  assign _T_8164 = _T_2880 | _T_2888; // @[NV_NVDLA_cbuf.scala 74:72:@1111.4]
  assign _T_8165 = _T_2896 | _T_2904; // @[NV_NVDLA_cbuf.scala 74:72:@1113.4]
  assign _T_8166 = _T_2912 | _T_2920; // @[NV_NVDLA_cbuf.scala 74:72:@1115.4]
  assign _T_8167 = _T_2928 | _T_2936; // @[NV_NVDLA_cbuf.scala 74:72:@1117.4]
  assign _T_8168 = _T_2944 | _T_2952; // @[NV_NVDLA_cbuf.scala 74:72:@1119.4]
  assign _T_8169 = _T_2960 | _T_2968; // @[NV_NVDLA_cbuf.scala 74:72:@1121.4]
  assign _T_8170 = _T_2976 | _T_2984; // @[NV_NVDLA_cbuf.scala 74:72:@1123.4]
  assign _T_8171 = _T_2992 | _T_3000; // @[NV_NVDLA_cbuf.scala 74:72:@1125.4]
  assign _T_8172 = _T_3008 | _T_3016; // @[NV_NVDLA_cbuf.scala 74:72:@1127.4]
  assign _T_8173 = _T_3024 | _T_3032; // @[NV_NVDLA_cbuf.scala 74:72:@1129.4]
  assign _T_8174 = _T_3040 | _T_3048; // @[NV_NVDLA_cbuf.scala 74:72:@1131.4]
  assign _T_8175 = _T_3056 | _T_3064; // @[NV_NVDLA_cbuf.scala 74:72:@1133.4]
  assign _T_8176 = _T_3072 | _T_3080; // @[NV_NVDLA_cbuf.scala 74:72:@1135.4]
  assign _T_8177 = _T_3088 | _T_3096; // @[NV_NVDLA_cbuf.scala 74:72:@1137.4]
  assign _T_8178 = _T_3104 | _T_3112; // @[NV_NVDLA_cbuf.scala 74:72:@1139.4]
  assign _T_8179 = _T_3120 | _T_3128; // @[NV_NVDLA_cbuf.scala 74:72:@1141.4]
  assign _T_8180 = _T_3136 | _T_3144; // @[NV_NVDLA_cbuf.scala 74:72:@1143.4]
  assign _T_8181 = _T_3152 | _T_3160; // @[NV_NVDLA_cbuf.scala 74:72:@1145.4]
  assign _T_8182 = _T_3168 | _T_3176; // @[NV_NVDLA_cbuf.scala 74:72:@1147.4]
  assign _T_10708 = _T_2672 | _T_2688; // @[NV_NVDLA_cbuf.scala 89:68:@1240.4]
  assign _T_10709 = _T_2704 | _T_2720; // @[NV_NVDLA_cbuf.scala 89:68:@1242.4]
  assign _T_10710 = _T_2736 | _T_2752; // @[NV_NVDLA_cbuf.scala 89:68:@1244.4]
  assign _T_10711 = _T_2768 | _T_2784; // @[NV_NVDLA_cbuf.scala 89:68:@1246.4]
  assign _T_10712 = _T_2800 | _T_2816; // @[NV_NVDLA_cbuf.scala 89:68:@1248.4]
  assign _T_10713 = _T_2832 | _T_2848; // @[NV_NVDLA_cbuf.scala 89:68:@1250.4]
  assign _T_10714 = _T_2864 | _T_2880; // @[NV_NVDLA_cbuf.scala 89:68:@1252.4]
  assign _T_10715 = _T_2896 | _T_2912; // @[NV_NVDLA_cbuf.scala 89:68:@1254.4]
  assign _T_10716 = _T_2928 | _T_2944; // @[NV_NVDLA_cbuf.scala 89:68:@1256.4]
  assign _T_10717 = _T_2960 | _T_2976; // @[NV_NVDLA_cbuf.scala 89:68:@1258.4]
  assign _T_10718 = _T_2992 | _T_3008; // @[NV_NVDLA_cbuf.scala 89:68:@1260.4]
  assign _T_10719 = _T_3024 | _T_3040; // @[NV_NVDLA_cbuf.scala 89:68:@1262.4]
  assign _T_10720 = _T_3056 | _T_3072; // @[NV_NVDLA_cbuf.scala 89:68:@1264.4]
  assign _T_10721 = _T_3088 | _T_3104; // @[NV_NVDLA_cbuf.scala 89:68:@1266.4]
  assign _T_10722 = _T_3120 | _T_3136; // @[NV_NVDLA_cbuf.scala 89:68:@1268.4]
  assign _T_10723 = _T_3152 | _T_3168; // @[NV_NVDLA_cbuf.scala 89:68:@1270.4]
  assign _T_10724 = _T_2680 | _T_2696; // @[NV_NVDLA_cbuf.scala 89:68:@1272.4]
  assign _T_10725 = _T_2712 | _T_2728; // @[NV_NVDLA_cbuf.scala 89:68:@1274.4]
  assign _T_10726 = _T_2744 | _T_2760; // @[NV_NVDLA_cbuf.scala 89:68:@1276.4]
  assign _T_10727 = _T_2776 | _T_2792; // @[NV_NVDLA_cbuf.scala 89:68:@1278.4]
  assign _T_10728 = _T_2808 | _T_2824; // @[NV_NVDLA_cbuf.scala 89:68:@1280.4]
  assign _T_10729 = _T_2840 | _T_2856; // @[NV_NVDLA_cbuf.scala 89:68:@1282.4]
  assign _T_10730 = _T_2872 | _T_2888; // @[NV_NVDLA_cbuf.scala 89:68:@1284.4]
  assign _T_10731 = _T_2904 | _T_2920; // @[NV_NVDLA_cbuf.scala 89:68:@1286.4]
  assign _T_10732 = _T_2936 | _T_2952; // @[NV_NVDLA_cbuf.scala 89:68:@1288.4]
  assign _T_10733 = _T_2968 | _T_2984; // @[NV_NVDLA_cbuf.scala 89:68:@1290.4]
  assign _T_10734 = _T_3000 | _T_3016; // @[NV_NVDLA_cbuf.scala 89:68:@1292.4]
  assign _T_10735 = _T_3032 | _T_3048; // @[NV_NVDLA_cbuf.scala 89:68:@1294.4]
  assign _T_10736 = _T_3064 | _T_3080; // @[NV_NVDLA_cbuf.scala 89:68:@1296.4]
  assign _T_10737 = _T_3096 | _T_3112; // @[NV_NVDLA_cbuf.scala 89:68:@1298.4]
  assign _T_10738 = _T_3128 | _T_3144; // @[NV_NVDLA_cbuf.scala 89:68:@1300.4]
  assign _T_10739 = _T_3160 | _T_3176; // @[NV_NVDLA_cbuf.scala 89:68:@1302.4]
  assign _T_11345 = _T_9669_0_0 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1309.4]
  assign _T_11346 = _T_11345 & _T_8201_0; // @[NV_NVDLA_cbuf.scala 101:94:@1310.4]
  assign _T_11350 = _T_9669_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1313.4]
  assign _T_11351 = _T_11350 & _T_8215_0; // @[NV_NVDLA_cbuf.scala 102:97:@1314.4]
  assign _T_11355 = _T_9669_0_1 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1317.4]
  assign _T_11356 = _T_11355 & _T_8201_1; // @[NV_NVDLA_cbuf.scala 101:94:@1318.4]
  assign _T_11360 = _T_9669_0_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1321.4]
  assign _T_11361 = _T_11360 & _T_8215_1; // @[NV_NVDLA_cbuf.scala 102:97:@1322.4]
  assign _T_11362 = _T_11346 | _T_11356; // @[NV_NVDLA_cbuf.scala 104:68:@1324.4]
  assign _T_11367 = _T_9669_1_0 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1329.4]
  assign _T_11368 = _T_11367 & _T_8201_0; // @[NV_NVDLA_cbuf.scala 101:94:@1330.4]
  assign _T_11372 = _T_9669_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1333.4]
  assign _T_11373 = _T_11372 & _T_8215_0; // @[NV_NVDLA_cbuf.scala 102:97:@1334.4]
  assign _T_11377 = _T_9669_1_1 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1337.4]
  assign _T_11378 = _T_11377 & _T_8201_1; // @[NV_NVDLA_cbuf.scala 101:94:@1338.4]
  assign _T_11382 = _T_9669_1_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1341.4]
  assign _T_11383 = _T_11382 & _T_8215_1; // @[NV_NVDLA_cbuf.scala 102:97:@1342.4]
  assign _T_11384 = _T_11368 | _T_11378; // @[NV_NVDLA_cbuf.scala 104:68:@1344.4]
  assign _T_11389 = _T_9669_2_0 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1349.4]
  assign _T_11390 = _T_11389 & _T_8201_0; // @[NV_NVDLA_cbuf.scala 101:94:@1350.4]
  assign _T_11394 = _T_9669_2_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1353.4]
  assign _T_11395 = _T_11394 & _T_8215_0; // @[NV_NVDLA_cbuf.scala 102:97:@1354.4]
  assign _T_11399 = _T_9669_2_1 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1357.4]
  assign _T_11400 = _T_11399 & _T_8201_1; // @[NV_NVDLA_cbuf.scala 101:94:@1358.4]
  assign _T_11404 = _T_9669_2_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1361.4]
  assign _T_11405 = _T_11404 & _T_8215_1; // @[NV_NVDLA_cbuf.scala 102:97:@1362.4]
  assign _T_11406 = _T_11390 | _T_11400; // @[NV_NVDLA_cbuf.scala 104:68:@1364.4]
  assign _T_11411 = _T_9669_3_0 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1369.4]
  assign _T_11412 = _T_11411 & _T_8201_0; // @[NV_NVDLA_cbuf.scala 101:94:@1370.4]
  assign _T_11416 = _T_9669_3_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1373.4]
  assign _T_11417 = _T_11416 & _T_8215_0; // @[NV_NVDLA_cbuf.scala 102:97:@1374.4]
  assign _T_11421 = _T_9669_3_1 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1377.4]
  assign _T_11422 = _T_11421 & _T_8201_1; // @[NV_NVDLA_cbuf.scala 101:94:@1378.4]
  assign _T_11426 = _T_9669_3_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1381.4]
  assign _T_11427 = _T_11426 & _T_8215_1; // @[NV_NVDLA_cbuf.scala 102:97:@1382.4]
  assign _T_11428 = _T_11412 | _T_11422; // @[NV_NVDLA_cbuf.scala 104:68:@1384.4]
  assign _T_11433 = _T_9669_4_0 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1389.4]
  assign _T_11434 = _T_11433 & _T_8201_0; // @[NV_NVDLA_cbuf.scala 101:94:@1390.4]
  assign _T_11438 = _T_9669_4_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1393.4]
  assign _T_11439 = _T_11438 & _T_8215_0; // @[NV_NVDLA_cbuf.scala 102:97:@1394.4]
  assign _T_11443 = _T_9669_4_1 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1397.4]
  assign _T_11444 = _T_11443 & _T_8201_1; // @[NV_NVDLA_cbuf.scala 101:94:@1398.4]
  assign _T_11448 = _T_9669_4_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1401.4]
  assign _T_11449 = _T_11448 & _T_8215_1; // @[NV_NVDLA_cbuf.scala 102:97:@1402.4]
  assign _T_11450 = _T_11434 | _T_11444; // @[NV_NVDLA_cbuf.scala 104:68:@1404.4]
  assign _T_11455 = _T_9669_5_0 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1409.4]
  assign _T_11456 = _T_11455 & _T_8201_0; // @[NV_NVDLA_cbuf.scala 101:94:@1410.4]
  assign _T_11460 = _T_9669_5_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1413.4]
  assign _T_11461 = _T_11460 & _T_8215_0; // @[NV_NVDLA_cbuf.scala 102:97:@1414.4]
  assign _T_11465 = _T_9669_5_1 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1417.4]
  assign _T_11466 = _T_11465 & _T_8201_1; // @[NV_NVDLA_cbuf.scala 101:94:@1418.4]
  assign _T_11470 = _T_9669_5_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1421.4]
  assign _T_11471 = _T_11470 & _T_8215_1; // @[NV_NVDLA_cbuf.scala 102:97:@1422.4]
  assign _T_11472 = _T_11456 | _T_11466; // @[NV_NVDLA_cbuf.scala 104:68:@1424.4]
  assign _T_11477 = _T_9669_6_0 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1429.4]
  assign _T_11478 = _T_11477 & _T_8201_0; // @[NV_NVDLA_cbuf.scala 101:94:@1430.4]
  assign _T_11482 = _T_9669_6_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1433.4]
  assign _T_11483 = _T_11482 & _T_8215_0; // @[NV_NVDLA_cbuf.scala 102:97:@1434.4]
  assign _T_11487 = _T_9669_6_1 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1437.4]
  assign _T_11488 = _T_11487 & _T_8201_1; // @[NV_NVDLA_cbuf.scala 101:94:@1438.4]
  assign _T_11492 = _T_9669_6_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1441.4]
  assign _T_11493 = _T_11492 & _T_8215_1; // @[NV_NVDLA_cbuf.scala 102:97:@1442.4]
  assign _T_11494 = _T_11478 | _T_11488; // @[NV_NVDLA_cbuf.scala 104:68:@1444.4]
  assign _T_11499 = _T_9669_7_0 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1449.4]
  assign _T_11500 = _T_11499 & _T_8201_0; // @[NV_NVDLA_cbuf.scala 101:94:@1450.4]
  assign _T_11504 = _T_9669_7_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1453.4]
  assign _T_11505 = _T_11504 & _T_8215_0; // @[NV_NVDLA_cbuf.scala 102:97:@1454.4]
  assign _T_11509 = _T_9669_7_1 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1457.4]
  assign _T_11510 = _T_11509 & _T_8201_1; // @[NV_NVDLA_cbuf.scala 101:94:@1458.4]
  assign _T_11514 = _T_9669_7_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1461.4]
  assign _T_11515 = _T_11514 & _T_8215_1; // @[NV_NVDLA_cbuf.scala 102:97:@1462.4]
  assign _T_11516 = _T_11500 | _T_11510; // @[NV_NVDLA_cbuf.scala 104:68:@1464.4]
  assign _T_11521 = _T_9669_8_0 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1469.4]
  assign _T_11522 = _T_11521 & _T_8201_0; // @[NV_NVDLA_cbuf.scala 101:94:@1470.4]
  assign _T_11526 = _T_9669_8_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1473.4]
  assign _T_11527 = _T_11526 & _T_8215_0; // @[NV_NVDLA_cbuf.scala 102:97:@1474.4]
  assign _T_11531 = _T_9669_8_1 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1477.4]
  assign _T_11532 = _T_11531 & _T_8201_1; // @[NV_NVDLA_cbuf.scala 101:94:@1478.4]
  assign _T_11536 = _T_9669_8_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1481.4]
  assign _T_11537 = _T_11536 & _T_8215_1; // @[NV_NVDLA_cbuf.scala 102:97:@1482.4]
  assign _T_11538 = _T_11522 | _T_11532; // @[NV_NVDLA_cbuf.scala 104:68:@1484.4]
  assign _T_11543 = _T_9669_9_0 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1489.4]
  assign _T_11544 = _T_11543 & _T_8201_0; // @[NV_NVDLA_cbuf.scala 101:94:@1490.4]
  assign _T_11548 = _T_9669_9_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1493.4]
  assign _T_11549 = _T_11548 & _T_8215_0; // @[NV_NVDLA_cbuf.scala 102:97:@1494.4]
  assign _T_11553 = _T_9669_9_1 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1497.4]
  assign _T_11554 = _T_11553 & _T_8201_1; // @[NV_NVDLA_cbuf.scala 101:94:@1498.4]
  assign _T_11558 = _T_9669_9_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1501.4]
  assign _T_11559 = _T_11558 & _T_8215_1; // @[NV_NVDLA_cbuf.scala 102:97:@1502.4]
  assign _T_11560 = _T_11544 | _T_11554; // @[NV_NVDLA_cbuf.scala 104:68:@1504.4]
  assign _T_11565 = _T_9669_10_0 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1509.4]
  assign _T_11566 = _T_11565 & _T_8201_0; // @[NV_NVDLA_cbuf.scala 101:94:@1510.4]
  assign _T_11570 = _T_9669_10_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1513.4]
  assign _T_11571 = _T_11570 & _T_8215_0; // @[NV_NVDLA_cbuf.scala 102:97:@1514.4]
  assign _T_11575 = _T_9669_10_1 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1517.4]
  assign _T_11576 = _T_11575 & _T_8201_1; // @[NV_NVDLA_cbuf.scala 101:94:@1518.4]
  assign _T_11580 = _T_9669_10_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1521.4]
  assign _T_11581 = _T_11580 & _T_8215_1; // @[NV_NVDLA_cbuf.scala 102:97:@1522.4]
  assign _T_11582 = _T_11566 | _T_11576; // @[NV_NVDLA_cbuf.scala 104:68:@1524.4]
  assign _T_11587 = _T_9669_11_0 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1529.4]
  assign _T_11588 = _T_11587 & _T_8201_0; // @[NV_NVDLA_cbuf.scala 101:94:@1530.4]
  assign _T_11592 = _T_9669_11_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1533.4]
  assign _T_11593 = _T_11592 & _T_8215_0; // @[NV_NVDLA_cbuf.scala 102:97:@1534.4]
  assign _T_11597 = _T_9669_11_1 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1537.4]
  assign _T_11598 = _T_11597 & _T_8201_1; // @[NV_NVDLA_cbuf.scala 101:94:@1538.4]
  assign _T_11602 = _T_9669_11_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1541.4]
  assign _T_11603 = _T_11602 & _T_8215_1; // @[NV_NVDLA_cbuf.scala 102:97:@1542.4]
  assign _T_11604 = _T_11588 | _T_11598; // @[NV_NVDLA_cbuf.scala 104:68:@1544.4]
  assign _T_11609 = _T_9669_12_0 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1549.4]
  assign _T_11610 = _T_11609 & _T_8201_0; // @[NV_NVDLA_cbuf.scala 101:94:@1550.4]
  assign _T_11614 = _T_9669_12_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1553.4]
  assign _T_11615 = _T_11614 & _T_8215_0; // @[NV_NVDLA_cbuf.scala 102:97:@1554.4]
  assign _T_11619 = _T_9669_12_1 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1557.4]
  assign _T_11620 = _T_11619 & _T_8201_1; // @[NV_NVDLA_cbuf.scala 101:94:@1558.4]
  assign _T_11624 = _T_9669_12_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1561.4]
  assign _T_11625 = _T_11624 & _T_8215_1; // @[NV_NVDLA_cbuf.scala 102:97:@1562.4]
  assign _T_11626 = _T_11610 | _T_11620; // @[NV_NVDLA_cbuf.scala 104:68:@1564.4]
  assign _T_11631 = _T_9669_13_0 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1569.4]
  assign _T_11632 = _T_11631 & _T_8201_0; // @[NV_NVDLA_cbuf.scala 101:94:@1570.4]
  assign _T_11636 = _T_9669_13_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1573.4]
  assign _T_11637 = _T_11636 & _T_8215_0; // @[NV_NVDLA_cbuf.scala 102:97:@1574.4]
  assign _T_11641 = _T_9669_13_1 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1577.4]
  assign _T_11642 = _T_11641 & _T_8201_1; // @[NV_NVDLA_cbuf.scala 101:94:@1578.4]
  assign _T_11646 = _T_9669_13_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1581.4]
  assign _T_11647 = _T_11646 & _T_8215_1; // @[NV_NVDLA_cbuf.scala 102:97:@1582.4]
  assign _T_11648 = _T_11632 | _T_11642; // @[NV_NVDLA_cbuf.scala 104:68:@1584.4]
  assign _T_11653 = _T_9669_14_0 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1589.4]
  assign _T_11654 = _T_11653 & _T_8201_0; // @[NV_NVDLA_cbuf.scala 101:94:@1590.4]
  assign _T_11658 = _T_9669_14_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1593.4]
  assign _T_11659 = _T_11658 & _T_8215_0; // @[NV_NVDLA_cbuf.scala 102:97:@1594.4]
  assign _T_11663 = _T_9669_14_1 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1597.4]
  assign _T_11664 = _T_11663 & _T_8201_1; // @[NV_NVDLA_cbuf.scala 101:94:@1598.4]
  assign _T_11668 = _T_9669_14_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1601.4]
  assign _T_11669 = _T_11668 & _T_8215_1; // @[NV_NVDLA_cbuf.scala 102:97:@1602.4]
  assign _T_11670 = _T_11654 | _T_11664; // @[NV_NVDLA_cbuf.scala 104:68:@1604.4]
  assign _T_11675 = _T_9669_15_0 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1609.4]
  assign _T_11676 = _T_11675 & _T_8201_0; // @[NV_NVDLA_cbuf.scala 101:94:@1610.4]
  assign _T_11680 = _T_9669_15_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1613.4]
  assign _T_11681 = _T_11680 & _T_8215_0; // @[NV_NVDLA_cbuf.scala 102:97:@1614.4]
  assign _T_11685 = _T_9669_15_1 ? 13'h1fff : 13'h0; // @[Bitwise.scala 72:12:@1617.4]
  assign _T_11686 = _T_11685 & _T_8201_1; // @[NV_NVDLA_cbuf.scala 101:94:@1618.4]
  assign _T_11690 = _T_9669_15_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@1621.4]
  assign _T_11691 = _T_11690 & _T_8215_1; // @[NV_NVDLA_cbuf.scala 102:97:@1622.4]
  assign _T_11692 = _T_11676 | _T_11686; // @[NV_NVDLA_cbuf.scala 104:68:@1624.4]
  assign _T_12252 = _T_11362[8:0]; // @[NV_NVDLA_cbuf.scala 114:63:@1630.4]
  assign _T_12254 = _T_11384[8:0]; // @[NV_NVDLA_cbuf.scala 114:63:@1636.4]
  assign _T_12256 = _T_11406[8:0]; // @[NV_NVDLA_cbuf.scala 114:63:@1642.4]
  assign _T_12258 = _T_11428[8:0]; // @[NV_NVDLA_cbuf.scala 114:63:@1648.4]
  assign _T_12260 = _T_11450[8:0]; // @[NV_NVDLA_cbuf.scala 114:63:@1654.4]
  assign _T_12262 = _T_11472[8:0]; // @[NV_NVDLA_cbuf.scala 114:63:@1660.4]
  assign _T_12264 = _T_11494[8:0]; // @[NV_NVDLA_cbuf.scala 114:63:@1666.4]
  assign _T_12266 = _T_11516[8:0]; // @[NV_NVDLA_cbuf.scala 114:63:@1672.4]
  assign _T_12268 = _T_11538[8:0]; // @[NV_NVDLA_cbuf.scala 114:63:@1678.4]
  assign _T_12270 = _T_11560[8:0]; // @[NV_NVDLA_cbuf.scala 114:63:@1684.4]
  assign _T_12272 = _T_11582[8:0]; // @[NV_NVDLA_cbuf.scala 114:63:@1690.4]
  assign _T_12274 = _T_11604[8:0]; // @[NV_NVDLA_cbuf.scala 114:63:@1696.4]
  assign _T_12276 = _T_11626[8:0]; // @[NV_NVDLA_cbuf.scala 114:63:@1702.4]
  assign _T_12278 = _T_11648[8:0]; // @[NV_NVDLA_cbuf.scala 114:63:@1708.4]
  assign _T_12280 = _T_11670[8:0]; // @[NV_NVDLA_cbuf.scala 114:63:@1714.4]
  assign _T_12282 = _T_11692[8:0]; // @[NV_NVDLA_cbuf.scala 114:63:@1720.4]
  assign _T_19410 = io_sc2buf_dat_rd_addr_bits[12:9]; // @[NV_NVDLA_cbuf.scala 140:107:@1988.4]
  assign _T_19412 = _T_19410 == 4'h0; // @[NV_NVDLA_cbuf.scala 140:158:@1989.4]
  assign _T_19413 = io_sc2buf_dat_rd_addr_valid & _T_19412; // @[NV_NVDLA_cbuf.scala 140:78:@1990.4]
  assign _T_19420 = _T_19410 == 4'h1; // @[NV_NVDLA_cbuf.scala 140:158:@1997.4]
  assign _T_19421 = io_sc2buf_dat_rd_addr_valid & _T_19420; // @[NV_NVDLA_cbuf.scala 140:78:@1998.4]
  assign _T_19428 = _T_19410 == 4'h2; // @[NV_NVDLA_cbuf.scala 140:158:@2005.4]
  assign _T_19429 = io_sc2buf_dat_rd_addr_valid & _T_19428; // @[NV_NVDLA_cbuf.scala 140:78:@2006.4]
  assign _T_19436 = _T_19410 == 4'h3; // @[NV_NVDLA_cbuf.scala 140:158:@2013.4]
  assign _T_19437 = io_sc2buf_dat_rd_addr_valid & _T_19436; // @[NV_NVDLA_cbuf.scala 140:78:@2014.4]
  assign _T_19444 = _T_19410 == 4'h4; // @[NV_NVDLA_cbuf.scala 140:158:@2021.4]
  assign _T_19445 = io_sc2buf_dat_rd_addr_valid & _T_19444; // @[NV_NVDLA_cbuf.scala 140:78:@2022.4]
  assign _T_19452 = _T_19410 == 4'h5; // @[NV_NVDLA_cbuf.scala 140:158:@2029.4]
  assign _T_19453 = io_sc2buf_dat_rd_addr_valid & _T_19452; // @[NV_NVDLA_cbuf.scala 140:78:@2030.4]
  assign _T_19460 = _T_19410 == 4'h6; // @[NV_NVDLA_cbuf.scala 140:158:@2037.4]
  assign _T_19461 = io_sc2buf_dat_rd_addr_valid & _T_19460; // @[NV_NVDLA_cbuf.scala 140:78:@2038.4]
  assign _T_19468 = _T_19410 == 4'h7; // @[NV_NVDLA_cbuf.scala 140:158:@2045.4]
  assign _T_19469 = io_sc2buf_dat_rd_addr_valid & _T_19468; // @[NV_NVDLA_cbuf.scala 140:78:@2046.4]
  assign _T_19476 = _T_19410 == 4'h8; // @[NV_NVDLA_cbuf.scala 140:158:@2053.4]
  assign _T_19477 = io_sc2buf_dat_rd_addr_valid & _T_19476; // @[NV_NVDLA_cbuf.scala 140:78:@2054.4]
  assign _T_19484 = _T_19410 == 4'h9; // @[NV_NVDLA_cbuf.scala 140:158:@2061.4]
  assign _T_19485 = io_sc2buf_dat_rd_addr_valid & _T_19484; // @[NV_NVDLA_cbuf.scala 140:78:@2062.4]
  assign _T_19492 = _T_19410 == 4'ha; // @[NV_NVDLA_cbuf.scala 140:158:@2069.4]
  assign _T_19493 = io_sc2buf_dat_rd_addr_valid & _T_19492; // @[NV_NVDLA_cbuf.scala 140:78:@2070.4]
  assign _T_19500 = _T_19410 == 4'hb; // @[NV_NVDLA_cbuf.scala 140:158:@2077.4]
  assign _T_19501 = io_sc2buf_dat_rd_addr_valid & _T_19500; // @[NV_NVDLA_cbuf.scala 140:78:@2078.4]
  assign _T_19508 = _T_19410 == 4'hc; // @[NV_NVDLA_cbuf.scala 140:158:@2085.4]
  assign _T_19509 = io_sc2buf_dat_rd_addr_valid & _T_19508; // @[NV_NVDLA_cbuf.scala 140:78:@2086.4]
  assign _T_19516 = _T_19410 == 4'hd; // @[NV_NVDLA_cbuf.scala 140:158:@2093.4]
  assign _T_19517 = io_sc2buf_dat_rd_addr_valid & _T_19516; // @[NV_NVDLA_cbuf.scala 140:78:@2094.4]
  assign _T_19524 = _T_19410 == 4'he; // @[NV_NVDLA_cbuf.scala 140:158:@2101.4]
  assign _T_19525 = io_sc2buf_dat_rd_addr_valid & _T_19524; // @[NV_NVDLA_cbuf.scala 140:78:@2102.4]
  assign _T_19532 = _T_19410 == 4'hf; // @[NV_NVDLA_cbuf.scala 140:158:@2109.4]
  assign _T_19533 = io_sc2buf_dat_rd_addr_valid & _T_19532; // @[NV_NVDLA_cbuf.scala 140:78:@2110.4]
  assign _T_21412 = _T_19413 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2118.4]
  assign _T_21413 = io_sc2buf_dat_rd_addr_bits[8:0]; // @[NV_NVDLA_cbuf.scala 160:139:@2119.4]
  assign _T_21414 = _T_21412 & _T_21413; // @[NV_NVDLA_cbuf.scala 160:111:@2120.4]
  assign _T_21424 = _T_19421 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2128.4]
  assign _T_21426 = _T_21424 & _T_21413; // @[NV_NVDLA_cbuf.scala 160:111:@2130.4]
  assign _T_21436 = _T_19429 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2138.4]
  assign _T_21438 = _T_21436 & _T_21413; // @[NV_NVDLA_cbuf.scala 160:111:@2140.4]
  assign _T_21448 = _T_19437 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2148.4]
  assign _T_21450 = _T_21448 & _T_21413; // @[NV_NVDLA_cbuf.scala 160:111:@2150.4]
  assign _T_21460 = _T_19445 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2158.4]
  assign _T_21462 = _T_21460 & _T_21413; // @[NV_NVDLA_cbuf.scala 160:111:@2160.4]
  assign _T_21472 = _T_19453 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2168.4]
  assign _T_21474 = _T_21472 & _T_21413; // @[NV_NVDLA_cbuf.scala 160:111:@2170.4]
  assign _T_21484 = _T_19461 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2178.4]
  assign _T_21486 = _T_21484 & _T_21413; // @[NV_NVDLA_cbuf.scala 160:111:@2180.4]
  assign _T_21496 = _T_19469 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2188.4]
  assign _T_21498 = _T_21496 & _T_21413; // @[NV_NVDLA_cbuf.scala 160:111:@2190.4]
  assign _T_21508 = _T_19477 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2198.4]
  assign _T_21510 = _T_21508 & _T_21413; // @[NV_NVDLA_cbuf.scala 160:111:@2200.4]
  assign _T_21520 = _T_19485 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2208.4]
  assign _T_21522 = _T_21520 & _T_21413; // @[NV_NVDLA_cbuf.scala 160:111:@2210.4]
  assign _T_21532 = _T_19493 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2218.4]
  assign _T_21534 = _T_21532 & _T_21413; // @[NV_NVDLA_cbuf.scala 160:111:@2220.4]
  assign _T_21544 = _T_19501 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2228.4]
  assign _T_21546 = _T_21544 & _T_21413; // @[NV_NVDLA_cbuf.scala 160:111:@2230.4]
  assign _T_21556 = _T_19509 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2238.4]
  assign _T_21558 = _T_21556 & _T_21413; // @[NV_NVDLA_cbuf.scala 160:111:@2240.4]
  assign _T_21568 = _T_19517 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2248.4]
  assign _T_21570 = _T_21568 & _T_21413; // @[NV_NVDLA_cbuf.scala 160:111:@2250.4]
  assign _T_21580 = _T_19525 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2258.4]
  assign _T_21582 = _T_21580 & _T_21413; // @[NV_NVDLA_cbuf.scala 160:111:@2260.4]
  assign _T_21592 = _T_19533 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2268.4]
  assign _T_21594 = _T_21592 & _T_21413; // @[NV_NVDLA_cbuf.scala 160:111:@2270.4]
  assign _T_86681 = {_T_72478_3_1_0,_T_72478_3_0_0,_T_72478_2_1_0,_T_72478_2_0_0,_T_72478_1_1_0,_T_72478_1_0_0,_T_72478_0_1_0,_T_72478_0_0_0}; // @[NV_NVDLA_cbuf.scala 177:73:@2639.4]
  assign _T_86689 = {_T_72478_7_1_0,_T_72478_7_0_0,_T_72478_6_1_0,_T_72478_6_0_0,_T_72478_5_1_0,_T_72478_5_0_0,_T_72478_4_1_0,_T_72478_4_0_0,_T_86681}; // @[NV_NVDLA_cbuf.scala 177:73:@2647.4]
  assign _T_86696 = {_T_72478_11_1_0,_T_72478_11_0_0,_T_72478_10_1_0,_T_72478_10_0_0,_T_72478_9_1_0,_T_72478_9_0_0,_T_72478_8_1_0,_T_72478_8_0_0}; // @[NV_NVDLA_cbuf.scala 177:73:@2654.4]
  assign _T_86705 = {_T_72478_15_1_0,_T_72478_15_0_0,_T_72478_14_1_0,_T_72478_14_0_0,_T_72478_13_1_0,_T_72478_13_0_0,_T_72478_12_1_0,_T_72478_12_0_0,_T_86696,_T_86689}; // @[NV_NVDLA_cbuf.scala 177:73:@2663.4]
  assign _T_87210 = _T_72478_0_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2685.4]
  assign _T_86790_0_1 = nv_ram_rws_1_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@3950.4]
  assign _T_87211 = _T_86790_0_1 & _T_87210; // @[NV_NVDLA_cbuf.scala 197:68:@2686.4]
  assign _T_87215 = _T_72478_0_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2688.4]
  assign _T_86790_0_0 = nv_ram_rws_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@3941.4]
  assign _T_87216 = _T_86790_0_0 & _T_87215; // @[NV_NVDLA_cbuf.scala 198:65:@2689.4]
  assign _T_87221 = _T_72478_1_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2693.4]
  assign _T_86790_1_1 = nv_ram_rws_3_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@3968.4]
  assign _T_87222 = _T_86790_1_1 & _T_87221; // @[NV_NVDLA_cbuf.scala 197:68:@2694.4]
  assign _T_87226 = _T_72478_1_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2696.4]
  assign _T_86790_1_0 = nv_ram_rws_2_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@3959.4]
  assign _T_87227 = _T_86790_1_0 & _T_87226; // @[NV_NVDLA_cbuf.scala 198:65:@2697.4]
  assign _T_87232 = _T_72478_2_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2701.4]
  assign _T_86790_2_1 = nv_ram_rws_5_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@3986.4]
  assign _T_87233 = _T_86790_2_1 & _T_87232; // @[NV_NVDLA_cbuf.scala 197:68:@2702.4]
  assign _T_87237 = _T_72478_2_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2704.4]
  assign _T_86790_2_0 = nv_ram_rws_4_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@3977.4]
  assign _T_87238 = _T_86790_2_0 & _T_87237; // @[NV_NVDLA_cbuf.scala 198:65:@2705.4]
  assign _T_87243 = _T_72478_3_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2709.4]
  assign _T_86790_3_1 = nv_ram_rws_7_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4004.4]
  assign _T_87244 = _T_86790_3_1 & _T_87243; // @[NV_NVDLA_cbuf.scala 197:68:@2710.4]
  assign _T_87248 = _T_72478_3_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2712.4]
  assign _T_86790_3_0 = nv_ram_rws_6_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@3995.4]
  assign _T_87249 = _T_86790_3_0 & _T_87248; // @[NV_NVDLA_cbuf.scala 198:65:@2713.4]
  assign _T_87254 = _T_72478_4_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2717.4]
  assign _T_86790_4_1 = nv_ram_rws_9_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4022.4]
  assign _T_87255 = _T_86790_4_1 & _T_87254; // @[NV_NVDLA_cbuf.scala 197:68:@2718.4]
  assign _T_87259 = _T_72478_4_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2720.4]
  assign _T_86790_4_0 = nv_ram_rws_8_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4013.4]
  assign _T_87260 = _T_86790_4_0 & _T_87259; // @[NV_NVDLA_cbuf.scala 198:65:@2721.4]
  assign _T_87265 = _T_72478_5_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2725.4]
  assign _T_86790_5_1 = nv_ram_rws_11_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4040.4]
  assign _T_87266 = _T_86790_5_1 & _T_87265; // @[NV_NVDLA_cbuf.scala 197:68:@2726.4]
  assign _T_87270 = _T_72478_5_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2728.4]
  assign _T_86790_5_0 = nv_ram_rws_10_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4031.4]
  assign _T_87271 = _T_86790_5_0 & _T_87270; // @[NV_NVDLA_cbuf.scala 198:65:@2729.4]
  assign _T_87276 = _T_72478_6_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2733.4]
  assign _T_86790_6_1 = nv_ram_rws_13_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4058.4]
  assign _T_87277 = _T_86790_6_1 & _T_87276; // @[NV_NVDLA_cbuf.scala 197:68:@2734.4]
  assign _T_87281 = _T_72478_6_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2736.4]
  assign _T_86790_6_0 = nv_ram_rws_12_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4049.4]
  assign _T_87282 = _T_86790_6_0 & _T_87281; // @[NV_NVDLA_cbuf.scala 198:65:@2737.4]
  assign _T_87287 = _T_72478_7_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2741.4]
  assign _T_86790_7_1 = nv_ram_rws_15_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4076.4]
  assign _T_87288 = _T_86790_7_1 & _T_87287; // @[NV_NVDLA_cbuf.scala 197:68:@2742.4]
  assign _T_87292 = _T_72478_7_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2744.4]
  assign _T_86790_7_0 = nv_ram_rws_14_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4067.4]
  assign _T_87293 = _T_86790_7_0 & _T_87292; // @[NV_NVDLA_cbuf.scala 198:65:@2745.4]
  assign _T_87298 = _T_72478_8_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2749.4]
  assign _T_86790_8_1 = nv_ram_rws_17_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4094.4]
  assign _T_87299 = _T_86790_8_1 & _T_87298; // @[NV_NVDLA_cbuf.scala 197:68:@2750.4]
  assign _T_87303 = _T_72478_8_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2752.4]
  assign _T_86790_8_0 = nv_ram_rws_16_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4085.4]
  assign _T_87304 = _T_86790_8_0 & _T_87303; // @[NV_NVDLA_cbuf.scala 198:65:@2753.4]
  assign _T_87309 = _T_72478_9_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2757.4]
  assign _T_86790_9_1 = nv_ram_rws_19_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4112.4]
  assign _T_87310 = _T_86790_9_1 & _T_87309; // @[NV_NVDLA_cbuf.scala 197:68:@2758.4]
  assign _T_87314 = _T_72478_9_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2760.4]
  assign _T_86790_9_0 = nv_ram_rws_18_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4103.4]
  assign _T_87315 = _T_86790_9_0 & _T_87314; // @[NV_NVDLA_cbuf.scala 198:65:@2761.4]
  assign _T_87320 = _T_72478_10_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2765.4]
  assign _T_86790_10_1 = nv_ram_rws_21_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4130.4]
  assign _T_87321 = _T_86790_10_1 & _T_87320; // @[NV_NVDLA_cbuf.scala 197:68:@2766.4]
  assign _T_87325 = _T_72478_10_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2768.4]
  assign _T_86790_10_0 = nv_ram_rws_20_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4121.4]
  assign _T_87326 = _T_86790_10_0 & _T_87325; // @[NV_NVDLA_cbuf.scala 198:65:@2769.4]
  assign _T_87331 = _T_72478_11_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2773.4]
  assign _T_86790_11_1 = nv_ram_rws_23_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4148.4]
  assign _T_87332 = _T_86790_11_1 & _T_87331; // @[NV_NVDLA_cbuf.scala 197:68:@2774.4]
  assign _T_87336 = _T_72478_11_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2776.4]
  assign _T_86790_11_0 = nv_ram_rws_22_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4139.4]
  assign _T_87337 = _T_86790_11_0 & _T_87336; // @[NV_NVDLA_cbuf.scala 198:65:@2777.4]
  assign _T_87342 = _T_72478_12_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2781.4]
  assign _T_86790_12_1 = nv_ram_rws_25_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4166.4]
  assign _T_87343 = _T_86790_12_1 & _T_87342; // @[NV_NVDLA_cbuf.scala 197:68:@2782.4]
  assign _T_87347 = _T_72478_12_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2784.4]
  assign _T_86790_12_0 = nv_ram_rws_24_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4157.4]
  assign _T_87348 = _T_86790_12_0 & _T_87347; // @[NV_NVDLA_cbuf.scala 198:65:@2785.4]
  assign _T_87353 = _T_72478_13_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2789.4]
  assign _T_86790_13_1 = nv_ram_rws_27_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4184.4]
  assign _T_87354 = _T_86790_13_1 & _T_87353; // @[NV_NVDLA_cbuf.scala 197:68:@2790.4]
  assign _T_87358 = _T_72478_13_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2792.4]
  assign _T_86790_13_0 = nv_ram_rws_26_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4175.4]
  assign _T_87359 = _T_86790_13_0 & _T_87358; // @[NV_NVDLA_cbuf.scala 198:65:@2793.4]
  assign _T_87364 = _T_72478_14_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2797.4]
  assign _T_86790_14_1 = nv_ram_rws_29_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4202.4]
  assign _T_87365 = _T_86790_14_1 & _T_87364; // @[NV_NVDLA_cbuf.scala 197:68:@2798.4]
  assign _T_87369 = _T_72478_14_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2800.4]
  assign _T_86790_14_0 = nv_ram_rws_28_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4193.4]
  assign _T_87370 = _T_86790_14_0 & _T_87369; // @[NV_NVDLA_cbuf.scala 198:65:@2801.4]
  assign _T_87375 = _T_72478_15_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2805.4]
  assign _T_86790_15_1 = nv_ram_rws_31_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4220.4]
  assign _T_87376 = _T_86790_15_1 & _T_87375; // @[NV_NVDLA_cbuf.scala 197:68:@2806.4]
  assign _T_87380 = _T_72478_15_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@2808.4]
  assign _T_86790_15_0 = nv_ram_rws_30_io_dout; // @[NV_NVDLA_cbuf.scala 179:32:@2682.4 NV_NVDLA_cbuf.scala 399:35:@4211.4]
  assign _T_87381 = _T_86790_15_0 & _T_87380; // @[NV_NVDLA_cbuf.scala 198:65:@2809.4]
  assign _T_88202 = _T_87674_0_0 | _T_87674_1_0; // @[NV_NVDLA_cbuf.scala 237:67:@2830.4]
  assign _T_88203 = _T_88202 | _T_87674_2_0; // @[NV_NVDLA_cbuf.scala 237:98:@2831.4]
  assign _T_88205 = _T_87674_4_0 | _T_87674_5_0; // @[NV_NVDLA_cbuf.scala 237:67:@2834.4]
  assign _T_88206 = _T_88205 | _T_87674_6_0; // @[NV_NVDLA_cbuf.scala 237:98:@2835.4]
  assign _T_88208 = _T_87674_8_0 | _T_87674_9_0; // @[NV_NVDLA_cbuf.scala 237:67:@2838.4]
  assign _T_88209 = _T_88208 | _T_87674_10_0; // @[NV_NVDLA_cbuf.scala 237:98:@2839.4]
  assign _T_88211 = _T_87674_12_0 | _T_87674_13_0; // @[NV_NVDLA_cbuf.scala 237:67:@2842.4]
  assign _T_88212 = _T_88211 | _T_87674_14_0; // @[NV_NVDLA_cbuf.scala 237:98:@2843.4]
  assign _T_88245 = _T_88155_0_0 | _T_88155_1_0; // @[NV_NVDLA_cbuf.scala 242:67:@2847.4]
  assign _T_88246 = _T_88245 | _T_88155_2_0; // @[NV_NVDLA_cbuf.scala 242:98:@2848.4]
  assign _T_88529 = io_sc2buf_wt_rd_addr_bits[12:9]; // @[NV_NVDLA_cbuf.scala 265:100:@2855.4]
  assign _T_88531 = _T_88529 == 4'h0; // @[NV_NVDLA_cbuf.scala 265:151:@2856.4]
  assign _T_88532 = io_sc2buf_wt_rd_addr_valid & _T_88531; // @[NV_NVDLA_cbuf.scala 265:72:@2857.4]
  assign _T_88539 = _T_88529 == 4'h1; // @[NV_NVDLA_cbuf.scala 265:151:@2864.4]
  assign _T_88540 = io_sc2buf_wt_rd_addr_valid & _T_88539; // @[NV_NVDLA_cbuf.scala 265:72:@2865.4]
  assign _T_88547 = _T_88529 == 4'h2; // @[NV_NVDLA_cbuf.scala 265:151:@2872.4]
  assign _T_88548 = io_sc2buf_wt_rd_addr_valid & _T_88547; // @[NV_NVDLA_cbuf.scala 265:72:@2873.4]
  assign _T_88555 = _T_88529 == 4'h3; // @[NV_NVDLA_cbuf.scala 265:151:@2880.4]
  assign _T_88556 = io_sc2buf_wt_rd_addr_valid & _T_88555; // @[NV_NVDLA_cbuf.scala 265:72:@2881.4]
  assign _T_88563 = _T_88529 == 4'h4; // @[NV_NVDLA_cbuf.scala 265:151:@2888.4]
  assign _T_88564 = io_sc2buf_wt_rd_addr_valid & _T_88563; // @[NV_NVDLA_cbuf.scala 265:72:@2889.4]
  assign _T_88571 = _T_88529 == 4'h5; // @[NV_NVDLA_cbuf.scala 265:151:@2896.4]
  assign _T_88572 = io_sc2buf_wt_rd_addr_valid & _T_88571; // @[NV_NVDLA_cbuf.scala 265:72:@2897.4]
  assign _T_88579 = _T_88529 == 4'h6; // @[NV_NVDLA_cbuf.scala 265:151:@2904.4]
  assign _T_88580 = io_sc2buf_wt_rd_addr_valid & _T_88579; // @[NV_NVDLA_cbuf.scala 265:72:@2905.4]
  assign _T_88587 = _T_88529 == 4'h7; // @[NV_NVDLA_cbuf.scala 265:151:@2912.4]
  assign _T_88588 = io_sc2buf_wt_rd_addr_valid & _T_88587; // @[NV_NVDLA_cbuf.scala 265:72:@2913.4]
  assign _T_88595 = _T_88529 == 4'h8; // @[NV_NVDLA_cbuf.scala 265:151:@2920.4]
  assign _T_88596 = io_sc2buf_wt_rd_addr_valid & _T_88595; // @[NV_NVDLA_cbuf.scala 265:72:@2921.4]
  assign _T_88603 = _T_88529 == 4'h9; // @[NV_NVDLA_cbuf.scala 265:151:@2928.4]
  assign _T_88604 = io_sc2buf_wt_rd_addr_valid & _T_88603; // @[NV_NVDLA_cbuf.scala 265:72:@2929.4]
  assign _T_88611 = _T_88529 == 4'ha; // @[NV_NVDLA_cbuf.scala 265:151:@2936.4]
  assign _T_88612 = io_sc2buf_wt_rd_addr_valid & _T_88611; // @[NV_NVDLA_cbuf.scala 265:72:@2937.4]
  assign _T_88619 = _T_88529 == 4'hb; // @[NV_NVDLA_cbuf.scala 265:151:@2944.4]
  assign _T_88620 = io_sc2buf_wt_rd_addr_valid & _T_88619; // @[NV_NVDLA_cbuf.scala 265:72:@2945.4]
  assign _T_88627 = _T_88529 == 4'hc; // @[NV_NVDLA_cbuf.scala 265:151:@2952.4]
  assign _T_88628 = io_sc2buf_wt_rd_addr_valid & _T_88627; // @[NV_NVDLA_cbuf.scala 265:72:@2953.4]
  assign _T_88635 = _T_88529 == 4'hd; // @[NV_NVDLA_cbuf.scala 265:151:@2960.4]
  assign _T_88636 = io_sc2buf_wt_rd_addr_valid & _T_88635; // @[NV_NVDLA_cbuf.scala 265:72:@2961.4]
  assign _T_88643 = _T_88529 == 4'he; // @[NV_NVDLA_cbuf.scala 265:151:@2968.4]
  assign _T_88644 = io_sc2buf_wt_rd_addr_valid & _T_88643; // @[NV_NVDLA_cbuf.scala 265:72:@2969.4]
  assign _T_88651 = _T_88529 == 4'hf; // @[NV_NVDLA_cbuf.scala 265:151:@2976.4]
  assign _T_88652 = io_sc2buf_wt_rd_addr_valid & _T_88651; // @[NV_NVDLA_cbuf.scala 265:72:@2977.4]
  assign _T_88939 = _T_88532 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2985.4]
  assign _T_88940 = io_sc2buf_wt_rd_addr_bits[8:0]; // @[NV_NVDLA_cbuf.scala 285:128:@2986.4]
  assign _T_88941 = _T_88939 & _T_88940; // @[NV_NVDLA_cbuf.scala 285:101:@2987.4]
  assign _T_88951 = _T_88540 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@2995.4]
  assign _T_88953 = _T_88951 & _T_88940; // @[NV_NVDLA_cbuf.scala 285:101:@2997.4]
  assign _T_88963 = _T_88548 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@3005.4]
  assign _T_88965 = _T_88963 & _T_88940; // @[NV_NVDLA_cbuf.scala 285:101:@3007.4]
  assign _T_88975 = _T_88556 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@3015.4]
  assign _T_88977 = _T_88975 & _T_88940; // @[NV_NVDLA_cbuf.scala 285:101:@3017.4]
  assign _T_88987 = _T_88564 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@3025.4]
  assign _T_88989 = _T_88987 & _T_88940; // @[NV_NVDLA_cbuf.scala 285:101:@3027.4]
  assign _T_88999 = _T_88572 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@3035.4]
  assign _T_89001 = _T_88999 & _T_88940; // @[NV_NVDLA_cbuf.scala 285:101:@3037.4]
  assign _T_89011 = _T_88580 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@3045.4]
  assign _T_89013 = _T_89011 & _T_88940; // @[NV_NVDLA_cbuf.scala 285:101:@3047.4]
  assign _T_89023 = _T_88588 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@3055.4]
  assign _T_89025 = _T_89023 & _T_88940; // @[NV_NVDLA_cbuf.scala 285:101:@3057.4]
  assign _T_89035 = _T_88596 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@3065.4]
  assign _T_89037 = _T_89035 & _T_88940; // @[NV_NVDLA_cbuf.scala 285:101:@3067.4]
  assign _T_89047 = _T_88604 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@3075.4]
  assign _T_89049 = _T_89047 & _T_88940; // @[NV_NVDLA_cbuf.scala 285:101:@3077.4]
  assign _T_89059 = _T_88612 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@3085.4]
  assign _T_89061 = _T_89059 & _T_88940; // @[NV_NVDLA_cbuf.scala 285:101:@3087.4]
  assign _T_89071 = _T_88620 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@3095.4]
  assign _T_89073 = _T_89071 & _T_88940; // @[NV_NVDLA_cbuf.scala 285:101:@3097.4]
  assign _T_89083 = _T_88628 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@3105.4]
  assign _T_89085 = _T_89083 & _T_88940; // @[NV_NVDLA_cbuf.scala 285:101:@3107.4]
  assign _T_89095 = _T_88636 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@3115.4]
  assign _T_89097 = _T_89095 & _T_88940; // @[NV_NVDLA_cbuf.scala 285:101:@3117.4]
  assign _T_89107 = _T_88644 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@3125.4]
  assign _T_89109 = _T_89107 & _T_88940; // @[NV_NVDLA_cbuf.scala 285:101:@3127.4]
  assign _T_89119 = _T_88652 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@3135.4]
  assign _T_89121 = _T_89119 & _T_88940; // @[NV_NVDLA_cbuf.scala 285:101:@3137.4]
  assign _T_92339 = {_T_91073_3_1,_T_91073_3_0,_T_91073_2_1,_T_91073_2_0,_T_91073_1_1,_T_91073_1_0,_T_91073_0_1,_T_91073_0_0}; // @[NV_NVDLA_cbuf.scala 298:70:@3220.4]
  assign _T_92347 = {_T_91073_7_1,_T_91073_7_0,_T_91073_6_1,_T_91073_6_0,_T_91073_5_1,_T_91073_5_0,_T_91073_4_1,_T_91073_4_0,_T_92339}; // @[NV_NVDLA_cbuf.scala 298:70:@3228.4]
  assign _T_92354 = {_T_91073_11_1,_T_91073_11_0,_T_91073_10_1,_T_91073_10_0,_T_91073_9_1,_T_91073_9_0,_T_91073_8_1,_T_91073_8_0}; // @[NV_NVDLA_cbuf.scala 298:70:@3235.4]
  assign _T_92363 = {_T_91073_15_1,_T_91073_15_0,_T_91073_14_1,_T_91073_14_0,_T_91073_13_1,_T_91073_13_0,_T_91073_12_1,_T_91073_12_0,_T_92354,_T_92347}; // @[NV_NVDLA_cbuf.scala 298:70:@3244.4]
  assign _T_92400 = _T_91073_0_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3265.4]
  assign _T_92401 = _T_86790_0_1 & _T_92400; // @[NV_NVDLA_cbuf.scala 315:63:@3266.4]
  assign _T_92405 = _T_91073_0_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3268.4]
  assign _T_92406 = _T_86790_0_0 & _T_92405; // @[NV_NVDLA_cbuf.scala 316:61:@3269.4]
  assign _T_92411 = _T_91073_1_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3273.4]
  assign _T_92412 = _T_86790_1_1 & _T_92411; // @[NV_NVDLA_cbuf.scala 315:63:@3274.4]
  assign _T_92416 = _T_91073_1_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3276.4]
  assign _T_92417 = _T_86790_1_0 & _T_92416; // @[NV_NVDLA_cbuf.scala 316:61:@3277.4]
  assign _T_92422 = _T_91073_2_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3281.4]
  assign _T_92423 = _T_86790_2_1 & _T_92422; // @[NV_NVDLA_cbuf.scala 315:63:@3282.4]
  assign _T_92427 = _T_91073_2_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3284.4]
  assign _T_92428 = _T_86790_2_0 & _T_92427; // @[NV_NVDLA_cbuf.scala 316:61:@3285.4]
  assign _T_92433 = _T_91073_3_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3289.4]
  assign _T_92434 = _T_86790_3_1 & _T_92433; // @[NV_NVDLA_cbuf.scala 315:63:@3290.4]
  assign _T_92438 = _T_91073_3_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3292.4]
  assign _T_92439 = _T_86790_3_0 & _T_92438; // @[NV_NVDLA_cbuf.scala 316:61:@3293.4]
  assign _T_92444 = _T_91073_4_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3297.4]
  assign _T_92445 = _T_86790_4_1 & _T_92444; // @[NV_NVDLA_cbuf.scala 315:63:@3298.4]
  assign _T_92449 = _T_91073_4_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3300.4]
  assign _T_92450 = _T_86790_4_0 & _T_92449; // @[NV_NVDLA_cbuf.scala 316:61:@3301.4]
  assign _T_92455 = _T_91073_5_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3305.4]
  assign _T_92456 = _T_86790_5_1 & _T_92455; // @[NV_NVDLA_cbuf.scala 315:63:@3306.4]
  assign _T_92460 = _T_91073_5_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3308.4]
  assign _T_92461 = _T_86790_5_0 & _T_92460; // @[NV_NVDLA_cbuf.scala 316:61:@3309.4]
  assign _T_92466 = _T_91073_6_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3313.4]
  assign _T_92467 = _T_86790_6_1 & _T_92466; // @[NV_NVDLA_cbuf.scala 315:63:@3314.4]
  assign _T_92471 = _T_91073_6_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3316.4]
  assign _T_92472 = _T_86790_6_0 & _T_92471; // @[NV_NVDLA_cbuf.scala 316:61:@3317.4]
  assign _T_92477 = _T_91073_7_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3321.4]
  assign _T_92478 = _T_86790_7_1 & _T_92477; // @[NV_NVDLA_cbuf.scala 315:63:@3322.4]
  assign _T_92482 = _T_91073_7_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3324.4]
  assign _T_92483 = _T_86790_7_0 & _T_92482; // @[NV_NVDLA_cbuf.scala 316:61:@3325.4]
  assign _T_92488 = _T_91073_8_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3329.4]
  assign _T_92489 = _T_86790_8_1 & _T_92488; // @[NV_NVDLA_cbuf.scala 315:63:@3330.4]
  assign _T_92493 = _T_91073_8_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3332.4]
  assign _T_92494 = _T_86790_8_0 & _T_92493; // @[NV_NVDLA_cbuf.scala 316:61:@3333.4]
  assign _T_92499 = _T_91073_9_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3337.4]
  assign _T_92500 = _T_86790_9_1 & _T_92499; // @[NV_NVDLA_cbuf.scala 315:63:@3338.4]
  assign _T_92504 = _T_91073_9_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3340.4]
  assign _T_92505 = _T_86790_9_0 & _T_92504; // @[NV_NVDLA_cbuf.scala 316:61:@3341.4]
  assign _T_92510 = _T_91073_10_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3345.4]
  assign _T_92511 = _T_86790_10_1 & _T_92510; // @[NV_NVDLA_cbuf.scala 315:63:@3346.4]
  assign _T_92515 = _T_91073_10_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3348.4]
  assign _T_92516 = _T_86790_10_0 & _T_92515; // @[NV_NVDLA_cbuf.scala 316:61:@3349.4]
  assign _T_92521 = _T_91073_11_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3353.4]
  assign _T_92522 = _T_86790_11_1 & _T_92521; // @[NV_NVDLA_cbuf.scala 315:63:@3354.4]
  assign _T_92526 = _T_91073_11_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3356.4]
  assign _T_92527 = _T_86790_11_0 & _T_92526; // @[NV_NVDLA_cbuf.scala 316:61:@3357.4]
  assign _T_92532 = _T_91073_12_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3361.4]
  assign _T_92533 = _T_86790_12_1 & _T_92532; // @[NV_NVDLA_cbuf.scala 315:63:@3362.4]
  assign _T_92537 = _T_91073_12_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3364.4]
  assign _T_92538 = _T_86790_12_0 & _T_92537; // @[NV_NVDLA_cbuf.scala 316:61:@3365.4]
  assign _T_92543 = _T_91073_13_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3369.4]
  assign _T_92544 = _T_86790_13_1 & _T_92543; // @[NV_NVDLA_cbuf.scala 315:63:@3370.4]
  assign _T_92548 = _T_91073_13_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3372.4]
  assign _T_92549 = _T_86790_13_0 & _T_92548; // @[NV_NVDLA_cbuf.scala 316:61:@3373.4]
  assign _T_92554 = _T_91073_14_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3377.4]
  assign _T_92555 = _T_86790_14_1 & _T_92554; // @[NV_NVDLA_cbuf.scala 315:63:@3378.4]
  assign _T_92559 = _T_91073_14_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3380.4]
  assign _T_92560 = _T_86790_14_0 & _T_92559; // @[NV_NVDLA_cbuf.scala 316:61:@3381.4]
  assign _T_92565 = _T_91073_15_1 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3385.4]
  assign _T_92566 = _T_86790_15_1 & _T_92565; // @[NV_NVDLA_cbuf.scala 315:63:@3386.4]
  assign _T_92570 = _T_91073_15_0 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@3388.4]
  assign _T_92571 = _T_86790_15_0 & _T_92570; // @[NV_NVDLA_cbuf.scala 316:61:@3389.4]
  assign _T_92672 = _T_92609_0 | _T_92609_1; // @[NV_NVDLA_cbuf.scala 354:57:@3410.4]
  assign _T_92673 = _T_92672 | _T_92609_2; // @[NV_NVDLA_cbuf.scala 354:83:@3411.4]
  assign _T_92675 = _T_92609_4 | _T_92609_5; // @[NV_NVDLA_cbuf.scala 354:57:@3414.4]
  assign _T_92676 = _T_92675 | _T_92609_6; // @[NV_NVDLA_cbuf.scala 354:83:@3415.4]
  assign _T_92678 = _T_92609_8 | _T_92609_9; // @[NV_NVDLA_cbuf.scala 354:57:@3418.4]
  assign _T_92679 = _T_92678 | _T_92609_10; // @[NV_NVDLA_cbuf.scala 354:83:@3419.4]
  assign _T_92681 = _T_92609_12 | _T_92609_13; // @[NV_NVDLA_cbuf.scala 354:57:@3422.4]
  assign _T_92682 = _T_92681 | _T_92609_14; // @[NV_NVDLA_cbuf.scala 354:83:@3423.4]
  assign _T_92691 = _T_92665_0 | _T_92665_1; // @[NV_NVDLA_cbuf.scala 359:57:@3427.4]
  assign _T_92692 = _T_92691 | _T_92665_2; // @[NV_NVDLA_cbuf.scala 359:83:@3428.4]
  assign _T_95463 = _T_19413 | _T_88532; // @[NV_NVDLA_cbuf.scala 382:68:@3517.4]
  assign _T_95468 = _T_21412 & _T_21414; // @[NV_NVDLA_cbuf.scala 383:103:@3521.4]
  assign _T_95473 = _T_88939 & _T_88941; // @[NV_NVDLA_cbuf.scala 384:98:@3524.4]
  assign _T_95487 = _T_19421 | _T_88540; // @[NV_NVDLA_cbuf.scala 382:68:@3537.4]
  assign _T_95492 = _T_21424 & _T_21426; // @[NV_NVDLA_cbuf.scala 383:103:@3541.4]
  assign _T_95497 = _T_88951 & _T_88953; // @[NV_NVDLA_cbuf.scala 384:98:@3544.4]
  assign _T_95511 = _T_19429 | _T_88548; // @[NV_NVDLA_cbuf.scala 382:68:@3557.4]
  assign _T_95516 = _T_21436 & _T_21438; // @[NV_NVDLA_cbuf.scala 383:103:@3561.4]
  assign _T_95521 = _T_88963 & _T_88965; // @[NV_NVDLA_cbuf.scala 384:98:@3564.4]
  assign _T_95535 = _T_19437 | _T_88556; // @[NV_NVDLA_cbuf.scala 382:68:@3577.4]
  assign _T_95540 = _T_21448 & _T_21450; // @[NV_NVDLA_cbuf.scala 383:103:@3581.4]
  assign _T_95545 = _T_88975 & _T_88977; // @[NV_NVDLA_cbuf.scala 384:98:@3584.4]
  assign _T_95559 = _T_19445 | _T_88564; // @[NV_NVDLA_cbuf.scala 382:68:@3597.4]
  assign _T_95564 = _T_21460 & _T_21462; // @[NV_NVDLA_cbuf.scala 383:103:@3601.4]
  assign _T_95569 = _T_88987 & _T_88989; // @[NV_NVDLA_cbuf.scala 384:98:@3604.4]
  assign _T_95583 = _T_19453 | _T_88572; // @[NV_NVDLA_cbuf.scala 382:68:@3617.4]
  assign _T_95588 = _T_21472 & _T_21474; // @[NV_NVDLA_cbuf.scala 383:103:@3621.4]
  assign _T_95593 = _T_88999 & _T_89001; // @[NV_NVDLA_cbuf.scala 384:98:@3624.4]
  assign _T_95607 = _T_19461 | _T_88580; // @[NV_NVDLA_cbuf.scala 382:68:@3637.4]
  assign _T_95612 = _T_21484 & _T_21486; // @[NV_NVDLA_cbuf.scala 383:103:@3641.4]
  assign _T_95617 = _T_89011 & _T_89013; // @[NV_NVDLA_cbuf.scala 384:98:@3644.4]
  assign _T_95631 = _T_19469 | _T_88588; // @[NV_NVDLA_cbuf.scala 382:68:@3657.4]
  assign _T_95636 = _T_21496 & _T_21498; // @[NV_NVDLA_cbuf.scala 383:103:@3661.4]
  assign _T_95641 = _T_89023 & _T_89025; // @[NV_NVDLA_cbuf.scala 384:98:@3664.4]
  assign _T_95655 = _T_19477 | _T_88596; // @[NV_NVDLA_cbuf.scala 382:68:@3677.4]
  assign _T_95660 = _T_21508 & _T_21510; // @[NV_NVDLA_cbuf.scala 383:103:@3681.4]
  assign _T_95665 = _T_89035 & _T_89037; // @[NV_NVDLA_cbuf.scala 384:98:@3684.4]
  assign _T_95679 = _T_19485 | _T_88604; // @[NV_NVDLA_cbuf.scala 382:68:@3697.4]
  assign _T_95684 = _T_21520 & _T_21522; // @[NV_NVDLA_cbuf.scala 383:103:@3701.4]
  assign _T_95689 = _T_89047 & _T_89049; // @[NV_NVDLA_cbuf.scala 384:98:@3704.4]
  assign _T_95703 = _T_19493 | _T_88612; // @[NV_NVDLA_cbuf.scala 382:68:@3717.4]
  assign _T_95708 = _T_21532 & _T_21534; // @[NV_NVDLA_cbuf.scala 383:103:@3721.4]
  assign _T_95713 = _T_89059 & _T_89061; // @[NV_NVDLA_cbuf.scala 384:98:@3724.4]
  assign _T_95727 = _T_19501 | _T_88620; // @[NV_NVDLA_cbuf.scala 382:68:@3737.4]
  assign _T_95732 = _T_21544 & _T_21546; // @[NV_NVDLA_cbuf.scala 383:103:@3741.4]
  assign _T_95737 = _T_89071 & _T_89073; // @[NV_NVDLA_cbuf.scala 384:98:@3744.4]
  assign _T_95751 = _T_19509 | _T_88628; // @[NV_NVDLA_cbuf.scala 382:68:@3757.4]
  assign _T_95756 = _T_21556 & _T_21558; // @[NV_NVDLA_cbuf.scala 383:103:@3761.4]
  assign _T_95761 = _T_89083 & _T_89085; // @[NV_NVDLA_cbuf.scala 384:98:@3764.4]
  assign _T_95775 = _T_19517 | _T_88636; // @[NV_NVDLA_cbuf.scala 382:68:@3777.4]
  assign _T_95780 = _T_21568 & _T_21570; // @[NV_NVDLA_cbuf.scala 383:103:@3781.4]
  assign _T_95785 = _T_89095 & _T_89097; // @[NV_NVDLA_cbuf.scala 384:98:@3784.4]
  assign _T_95799 = _T_19525 | _T_88644; // @[NV_NVDLA_cbuf.scala 382:68:@3797.4]
  assign _T_95804 = _T_21580 & _T_21582; // @[NV_NVDLA_cbuf.scala 383:103:@3801.4]
  assign _T_95809 = _T_89107 & _T_89109; // @[NV_NVDLA_cbuf.scala 384:98:@3804.4]
  assign _T_95823 = _T_19533 | _T_88652; // @[NV_NVDLA_cbuf.scala 382:68:@3817.4]
  assign _T_95828 = _T_21592 & _T_21594; // @[NV_NVDLA_cbuf.scala 383:103:@3821.4]
  assign _T_95833 = _T_89119 & _T_89121; // @[NV_NVDLA_cbuf.scala 384:98:@3824.4]
  assign io_sc2buf_dat_rd_data_valid = _T_86716; // @[NV_NVDLA_cbuf.scala 177:33:@2681.4]
  assign io_sc2buf_dat_rd_data_bits = _T_88249; // @[NV_NVDLA_cbuf.scala 254:32:@2853.4]
  assign io_sc2buf_wt_rd_data_valid = _T_92374; // @[NV_NVDLA_cbuf.scala 298:32:@3262.4]
  assign io_sc2buf_wt_rd_data_bits = _T_92695; // @[NV_NVDLA_cbuf.scala 370:31:@3433.4]
  assign nv_ram_rws_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@3933.4]
  assign nv_ram_rws_io_re = _T_94145_0_0; // @[NV_NVDLA_cbuf.scala 394:45:@3934.4]
  assign nv_ram_rws_io_we = _T_16500_0_0; // @[NV_NVDLA_cbuf.scala 396:45:@3937.4]
  assign nv_ram_rws_io_ra = _T_95257_0_0; // @[NV_NVDLA_cbuf.scala 395:45:@3936.4]
  assign nv_ram_rws_io_wa = _T_13733_0_0; // @[NV_NVDLA_cbuf.scala 397:45:@3939.4]
  assign nv_ram_rws_io_di = _T_14845_0_0; // @[NV_NVDLA_cbuf.scala 398:45:@3940.4]
  assign nv_ram_rws_1_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@3942.4]
  assign nv_ram_rws_1_io_re = _T_94145_0_1; // @[NV_NVDLA_cbuf.scala 394:45:@3943.4]
  assign nv_ram_rws_1_io_we = _T_16500_0_1; // @[NV_NVDLA_cbuf.scala 396:45:@3946.4]
  assign nv_ram_rws_1_io_ra = _T_95257_0_1; // @[NV_NVDLA_cbuf.scala 395:45:@3945.4]
  assign nv_ram_rws_1_io_wa = _T_13733_0_1; // @[NV_NVDLA_cbuf.scala 397:45:@3948.4]
  assign nv_ram_rws_1_io_di = _T_14845_0_1; // @[NV_NVDLA_cbuf.scala 398:45:@3949.4]
  assign nv_ram_rws_2_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@3951.4]
  assign nv_ram_rws_2_io_re = _T_94145_1_0; // @[NV_NVDLA_cbuf.scala 394:45:@3952.4]
  assign nv_ram_rws_2_io_we = _T_16500_1_0; // @[NV_NVDLA_cbuf.scala 396:45:@3955.4]
  assign nv_ram_rws_2_io_ra = _T_95257_1_0; // @[NV_NVDLA_cbuf.scala 395:45:@3954.4]
  assign nv_ram_rws_2_io_wa = _T_13733_1_0; // @[NV_NVDLA_cbuf.scala 397:45:@3957.4]
  assign nv_ram_rws_2_io_di = _T_14845_1_0; // @[NV_NVDLA_cbuf.scala 398:45:@3958.4]
  assign nv_ram_rws_3_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@3960.4]
  assign nv_ram_rws_3_io_re = _T_94145_1_1; // @[NV_NVDLA_cbuf.scala 394:45:@3961.4]
  assign nv_ram_rws_3_io_we = _T_16500_1_1; // @[NV_NVDLA_cbuf.scala 396:45:@3964.4]
  assign nv_ram_rws_3_io_ra = _T_95257_1_1; // @[NV_NVDLA_cbuf.scala 395:45:@3963.4]
  assign nv_ram_rws_3_io_wa = _T_13733_1_1; // @[NV_NVDLA_cbuf.scala 397:45:@3966.4]
  assign nv_ram_rws_3_io_di = _T_14845_1_1; // @[NV_NVDLA_cbuf.scala 398:45:@3967.4]
  assign nv_ram_rws_4_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@3969.4]
  assign nv_ram_rws_4_io_re = _T_94145_2_0; // @[NV_NVDLA_cbuf.scala 394:45:@3970.4]
  assign nv_ram_rws_4_io_we = _T_16500_2_0; // @[NV_NVDLA_cbuf.scala 396:45:@3973.4]
  assign nv_ram_rws_4_io_ra = _T_95257_2_0; // @[NV_NVDLA_cbuf.scala 395:45:@3972.4]
  assign nv_ram_rws_4_io_wa = _T_13733_2_0; // @[NV_NVDLA_cbuf.scala 397:45:@3975.4]
  assign nv_ram_rws_4_io_di = _T_14845_2_0; // @[NV_NVDLA_cbuf.scala 398:45:@3976.4]
  assign nv_ram_rws_5_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@3978.4]
  assign nv_ram_rws_5_io_re = _T_94145_2_1; // @[NV_NVDLA_cbuf.scala 394:45:@3979.4]
  assign nv_ram_rws_5_io_we = _T_16500_2_1; // @[NV_NVDLA_cbuf.scala 396:45:@3982.4]
  assign nv_ram_rws_5_io_ra = _T_95257_2_1; // @[NV_NVDLA_cbuf.scala 395:45:@3981.4]
  assign nv_ram_rws_5_io_wa = _T_13733_2_1; // @[NV_NVDLA_cbuf.scala 397:45:@3984.4]
  assign nv_ram_rws_5_io_di = _T_14845_2_1; // @[NV_NVDLA_cbuf.scala 398:45:@3985.4]
  assign nv_ram_rws_6_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@3987.4]
  assign nv_ram_rws_6_io_re = _T_94145_3_0; // @[NV_NVDLA_cbuf.scala 394:45:@3988.4]
  assign nv_ram_rws_6_io_we = _T_16500_3_0; // @[NV_NVDLA_cbuf.scala 396:45:@3991.4]
  assign nv_ram_rws_6_io_ra = _T_95257_3_0; // @[NV_NVDLA_cbuf.scala 395:45:@3990.4]
  assign nv_ram_rws_6_io_wa = _T_13733_3_0; // @[NV_NVDLA_cbuf.scala 397:45:@3993.4]
  assign nv_ram_rws_6_io_di = _T_14845_3_0; // @[NV_NVDLA_cbuf.scala 398:45:@3994.4]
  assign nv_ram_rws_7_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@3996.4]
  assign nv_ram_rws_7_io_re = _T_94145_3_1; // @[NV_NVDLA_cbuf.scala 394:45:@3997.4]
  assign nv_ram_rws_7_io_we = _T_16500_3_1; // @[NV_NVDLA_cbuf.scala 396:45:@4000.4]
  assign nv_ram_rws_7_io_ra = _T_95257_3_1; // @[NV_NVDLA_cbuf.scala 395:45:@3999.4]
  assign nv_ram_rws_7_io_wa = _T_13733_3_1; // @[NV_NVDLA_cbuf.scala 397:45:@4002.4]
  assign nv_ram_rws_7_io_di = _T_14845_3_1; // @[NV_NVDLA_cbuf.scala 398:45:@4003.4]
  assign nv_ram_rws_8_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4005.4]
  assign nv_ram_rws_8_io_re = _T_94145_4_0; // @[NV_NVDLA_cbuf.scala 394:45:@4006.4]
  assign nv_ram_rws_8_io_we = _T_16500_4_0; // @[NV_NVDLA_cbuf.scala 396:45:@4009.4]
  assign nv_ram_rws_8_io_ra = _T_95257_4_0; // @[NV_NVDLA_cbuf.scala 395:45:@4008.4]
  assign nv_ram_rws_8_io_wa = _T_13733_4_0; // @[NV_NVDLA_cbuf.scala 397:45:@4011.4]
  assign nv_ram_rws_8_io_di = _T_14845_4_0; // @[NV_NVDLA_cbuf.scala 398:45:@4012.4]
  assign nv_ram_rws_9_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4014.4]
  assign nv_ram_rws_9_io_re = _T_94145_4_1; // @[NV_NVDLA_cbuf.scala 394:45:@4015.4]
  assign nv_ram_rws_9_io_we = _T_16500_4_1; // @[NV_NVDLA_cbuf.scala 396:45:@4018.4]
  assign nv_ram_rws_9_io_ra = _T_95257_4_1; // @[NV_NVDLA_cbuf.scala 395:45:@4017.4]
  assign nv_ram_rws_9_io_wa = _T_13733_4_1; // @[NV_NVDLA_cbuf.scala 397:45:@4020.4]
  assign nv_ram_rws_9_io_di = _T_14845_4_1; // @[NV_NVDLA_cbuf.scala 398:45:@4021.4]
  assign nv_ram_rws_10_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4023.4]
  assign nv_ram_rws_10_io_re = _T_94145_5_0; // @[NV_NVDLA_cbuf.scala 394:45:@4024.4]
  assign nv_ram_rws_10_io_we = _T_16500_5_0; // @[NV_NVDLA_cbuf.scala 396:45:@4027.4]
  assign nv_ram_rws_10_io_ra = _T_95257_5_0; // @[NV_NVDLA_cbuf.scala 395:45:@4026.4]
  assign nv_ram_rws_10_io_wa = _T_13733_5_0; // @[NV_NVDLA_cbuf.scala 397:45:@4029.4]
  assign nv_ram_rws_10_io_di = _T_14845_5_0; // @[NV_NVDLA_cbuf.scala 398:45:@4030.4]
  assign nv_ram_rws_11_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4032.4]
  assign nv_ram_rws_11_io_re = _T_94145_5_1; // @[NV_NVDLA_cbuf.scala 394:45:@4033.4]
  assign nv_ram_rws_11_io_we = _T_16500_5_1; // @[NV_NVDLA_cbuf.scala 396:45:@4036.4]
  assign nv_ram_rws_11_io_ra = _T_95257_5_1; // @[NV_NVDLA_cbuf.scala 395:45:@4035.4]
  assign nv_ram_rws_11_io_wa = _T_13733_5_1; // @[NV_NVDLA_cbuf.scala 397:45:@4038.4]
  assign nv_ram_rws_11_io_di = _T_14845_5_1; // @[NV_NVDLA_cbuf.scala 398:45:@4039.4]
  assign nv_ram_rws_12_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4041.4]
  assign nv_ram_rws_12_io_re = _T_94145_6_0; // @[NV_NVDLA_cbuf.scala 394:45:@4042.4]
  assign nv_ram_rws_12_io_we = _T_16500_6_0; // @[NV_NVDLA_cbuf.scala 396:45:@4045.4]
  assign nv_ram_rws_12_io_ra = _T_95257_6_0; // @[NV_NVDLA_cbuf.scala 395:45:@4044.4]
  assign nv_ram_rws_12_io_wa = _T_13733_6_0; // @[NV_NVDLA_cbuf.scala 397:45:@4047.4]
  assign nv_ram_rws_12_io_di = _T_14845_6_0; // @[NV_NVDLA_cbuf.scala 398:45:@4048.4]
  assign nv_ram_rws_13_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4050.4]
  assign nv_ram_rws_13_io_re = _T_94145_6_1; // @[NV_NVDLA_cbuf.scala 394:45:@4051.4]
  assign nv_ram_rws_13_io_we = _T_16500_6_1; // @[NV_NVDLA_cbuf.scala 396:45:@4054.4]
  assign nv_ram_rws_13_io_ra = _T_95257_6_1; // @[NV_NVDLA_cbuf.scala 395:45:@4053.4]
  assign nv_ram_rws_13_io_wa = _T_13733_6_1; // @[NV_NVDLA_cbuf.scala 397:45:@4056.4]
  assign nv_ram_rws_13_io_di = _T_14845_6_1; // @[NV_NVDLA_cbuf.scala 398:45:@4057.4]
  assign nv_ram_rws_14_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4059.4]
  assign nv_ram_rws_14_io_re = _T_94145_7_0; // @[NV_NVDLA_cbuf.scala 394:45:@4060.4]
  assign nv_ram_rws_14_io_we = _T_16500_7_0; // @[NV_NVDLA_cbuf.scala 396:45:@4063.4]
  assign nv_ram_rws_14_io_ra = _T_95257_7_0; // @[NV_NVDLA_cbuf.scala 395:45:@4062.4]
  assign nv_ram_rws_14_io_wa = _T_13733_7_0; // @[NV_NVDLA_cbuf.scala 397:45:@4065.4]
  assign nv_ram_rws_14_io_di = _T_14845_7_0; // @[NV_NVDLA_cbuf.scala 398:45:@4066.4]
  assign nv_ram_rws_15_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4068.4]
  assign nv_ram_rws_15_io_re = _T_94145_7_1; // @[NV_NVDLA_cbuf.scala 394:45:@4069.4]
  assign nv_ram_rws_15_io_we = _T_16500_7_1; // @[NV_NVDLA_cbuf.scala 396:45:@4072.4]
  assign nv_ram_rws_15_io_ra = _T_95257_7_1; // @[NV_NVDLA_cbuf.scala 395:45:@4071.4]
  assign nv_ram_rws_15_io_wa = _T_13733_7_1; // @[NV_NVDLA_cbuf.scala 397:45:@4074.4]
  assign nv_ram_rws_15_io_di = _T_14845_7_1; // @[NV_NVDLA_cbuf.scala 398:45:@4075.4]
  assign nv_ram_rws_16_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4077.4]
  assign nv_ram_rws_16_io_re = _T_94145_8_0; // @[NV_NVDLA_cbuf.scala 394:45:@4078.4]
  assign nv_ram_rws_16_io_we = _T_16500_8_0; // @[NV_NVDLA_cbuf.scala 396:45:@4081.4]
  assign nv_ram_rws_16_io_ra = _T_95257_8_0; // @[NV_NVDLA_cbuf.scala 395:45:@4080.4]
  assign nv_ram_rws_16_io_wa = _T_13733_8_0; // @[NV_NVDLA_cbuf.scala 397:45:@4083.4]
  assign nv_ram_rws_16_io_di = _T_14845_8_0; // @[NV_NVDLA_cbuf.scala 398:45:@4084.4]
  assign nv_ram_rws_17_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4086.4]
  assign nv_ram_rws_17_io_re = _T_94145_8_1; // @[NV_NVDLA_cbuf.scala 394:45:@4087.4]
  assign nv_ram_rws_17_io_we = _T_16500_8_1; // @[NV_NVDLA_cbuf.scala 396:45:@4090.4]
  assign nv_ram_rws_17_io_ra = _T_95257_8_1; // @[NV_NVDLA_cbuf.scala 395:45:@4089.4]
  assign nv_ram_rws_17_io_wa = _T_13733_8_1; // @[NV_NVDLA_cbuf.scala 397:45:@4092.4]
  assign nv_ram_rws_17_io_di = _T_14845_8_1; // @[NV_NVDLA_cbuf.scala 398:45:@4093.4]
  assign nv_ram_rws_18_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4095.4]
  assign nv_ram_rws_18_io_re = _T_94145_9_0; // @[NV_NVDLA_cbuf.scala 394:45:@4096.4]
  assign nv_ram_rws_18_io_we = _T_16500_9_0; // @[NV_NVDLA_cbuf.scala 396:45:@4099.4]
  assign nv_ram_rws_18_io_ra = _T_95257_9_0; // @[NV_NVDLA_cbuf.scala 395:45:@4098.4]
  assign nv_ram_rws_18_io_wa = _T_13733_9_0; // @[NV_NVDLA_cbuf.scala 397:45:@4101.4]
  assign nv_ram_rws_18_io_di = _T_14845_9_0; // @[NV_NVDLA_cbuf.scala 398:45:@4102.4]
  assign nv_ram_rws_19_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4104.4]
  assign nv_ram_rws_19_io_re = _T_94145_9_1; // @[NV_NVDLA_cbuf.scala 394:45:@4105.4]
  assign nv_ram_rws_19_io_we = _T_16500_9_1; // @[NV_NVDLA_cbuf.scala 396:45:@4108.4]
  assign nv_ram_rws_19_io_ra = _T_95257_9_1; // @[NV_NVDLA_cbuf.scala 395:45:@4107.4]
  assign nv_ram_rws_19_io_wa = _T_13733_9_1; // @[NV_NVDLA_cbuf.scala 397:45:@4110.4]
  assign nv_ram_rws_19_io_di = _T_14845_9_1; // @[NV_NVDLA_cbuf.scala 398:45:@4111.4]
  assign nv_ram_rws_20_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4113.4]
  assign nv_ram_rws_20_io_re = _T_94145_10_0; // @[NV_NVDLA_cbuf.scala 394:45:@4114.4]
  assign nv_ram_rws_20_io_we = _T_16500_10_0; // @[NV_NVDLA_cbuf.scala 396:45:@4117.4]
  assign nv_ram_rws_20_io_ra = _T_95257_10_0; // @[NV_NVDLA_cbuf.scala 395:45:@4116.4]
  assign nv_ram_rws_20_io_wa = _T_13733_10_0; // @[NV_NVDLA_cbuf.scala 397:45:@4119.4]
  assign nv_ram_rws_20_io_di = _T_14845_10_0; // @[NV_NVDLA_cbuf.scala 398:45:@4120.4]
  assign nv_ram_rws_21_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4122.4]
  assign nv_ram_rws_21_io_re = _T_94145_10_1; // @[NV_NVDLA_cbuf.scala 394:45:@4123.4]
  assign nv_ram_rws_21_io_we = _T_16500_10_1; // @[NV_NVDLA_cbuf.scala 396:45:@4126.4]
  assign nv_ram_rws_21_io_ra = _T_95257_10_1; // @[NV_NVDLA_cbuf.scala 395:45:@4125.4]
  assign nv_ram_rws_21_io_wa = _T_13733_10_1; // @[NV_NVDLA_cbuf.scala 397:45:@4128.4]
  assign nv_ram_rws_21_io_di = _T_14845_10_1; // @[NV_NVDLA_cbuf.scala 398:45:@4129.4]
  assign nv_ram_rws_22_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4131.4]
  assign nv_ram_rws_22_io_re = _T_94145_11_0; // @[NV_NVDLA_cbuf.scala 394:45:@4132.4]
  assign nv_ram_rws_22_io_we = _T_16500_11_0; // @[NV_NVDLA_cbuf.scala 396:45:@4135.4]
  assign nv_ram_rws_22_io_ra = _T_95257_11_0; // @[NV_NVDLA_cbuf.scala 395:45:@4134.4]
  assign nv_ram_rws_22_io_wa = _T_13733_11_0; // @[NV_NVDLA_cbuf.scala 397:45:@4137.4]
  assign nv_ram_rws_22_io_di = _T_14845_11_0; // @[NV_NVDLA_cbuf.scala 398:45:@4138.4]
  assign nv_ram_rws_23_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4140.4]
  assign nv_ram_rws_23_io_re = _T_94145_11_1; // @[NV_NVDLA_cbuf.scala 394:45:@4141.4]
  assign nv_ram_rws_23_io_we = _T_16500_11_1; // @[NV_NVDLA_cbuf.scala 396:45:@4144.4]
  assign nv_ram_rws_23_io_ra = _T_95257_11_1; // @[NV_NVDLA_cbuf.scala 395:45:@4143.4]
  assign nv_ram_rws_23_io_wa = _T_13733_11_1; // @[NV_NVDLA_cbuf.scala 397:45:@4146.4]
  assign nv_ram_rws_23_io_di = _T_14845_11_1; // @[NV_NVDLA_cbuf.scala 398:45:@4147.4]
  assign nv_ram_rws_24_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4149.4]
  assign nv_ram_rws_24_io_re = _T_94145_12_0; // @[NV_NVDLA_cbuf.scala 394:45:@4150.4]
  assign nv_ram_rws_24_io_we = _T_16500_12_0; // @[NV_NVDLA_cbuf.scala 396:45:@4153.4]
  assign nv_ram_rws_24_io_ra = _T_95257_12_0; // @[NV_NVDLA_cbuf.scala 395:45:@4152.4]
  assign nv_ram_rws_24_io_wa = _T_13733_12_0; // @[NV_NVDLA_cbuf.scala 397:45:@4155.4]
  assign nv_ram_rws_24_io_di = _T_14845_12_0; // @[NV_NVDLA_cbuf.scala 398:45:@4156.4]
  assign nv_ram_rws_25_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4158.4]
  assign nv_ram_rws_25_io_re = _T_94145_12_1; // @[NV_NVDLA_cbuf.scala 394:45:@4159.4]
  assign nv_ram_rws_25_io_we = _T_16500_12_1; // @[NV_NVDLA_cbuf.scala 396:45:@4162.4]
  assign nv_ram_rws_25_io_ra = _T_95257_12_1; // @[NV_NVDLA_cbuf.scala 395:45:@4161.4]
  assign nv_ram_rws_25_io_wa = _T_13733_12_1; // @[NV_NVDLA_cbuf.scala 397:45:@4164.4]
  assign nv_ram_rws_25_io_di = _T_14845_12_1; // @[NV_NVDLA_cbuf.scala 398:45:@4165.4]
  assign nv_ram_rws_26_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4167.4]
  assign nv_ram_rws_26_io_re = _T_94145_13_0; // @[NV_NVDLA_cbuf.scala 394:45:@4168.4]
  assign nv_ram_rws_26_io_we = _T_16500_13_0; // @[NV_NVDLA_cbuf.scala 396:45:@4171.4]
  assign nv_ram_rws_26_io_ra = _T_95257_13_0; // @[NV_NVDLA_cbuf.scala 395:45:@4170.4]
  assign nv_ram_rws_26_io_wa = _T_13733_13_0; // @[NV_NVDLA_cbuf.scala 397:45:@4173.4]
  assign nv_ram_rws_26_io_di = _T_14845_13_0; // @[NV_NVDLA_cbuf.scala 398:45:@4174.4]
  assign nv_ram_rws_27_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4176.4]
  assign nv_ram_rws_27_io_re = _T_94145_13_1; // @[NV_NVDLA_cbuf.scala 394:45:@4177.4]
  assign nv_ram_rws_27_io_we = _T_16500_13_1; // @[NV_NVDLA_cbuf.scala 396:45:@4180.4]
  assign nv_ram_rws_27_io_ra = _T_95257_13_1; // @[NV_NVDLA_cbuf.scala 395:45:@4179.4]
  assign nv_ram_rws_27_io_wa = _T_13733_13_1; // @[NV_NVDLA_cbuf.scala 397:45:@4182.4]
  assign nv_ram_rws_27_io_di = _T_14845_13_1; // @[NV_NVDLA_cbuf.scala 398:45:@4183.4]
  assign nv_ram_rws_28_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4185.4]
  assign nv_ram_rws_28_io_re = _T_94145_14_0; // @[NV_NVDLA_cbuf.scala 394:45:@4186.4]
  assign nv_ram_rws_28_io_we = _T_16500_14_0; // @[NV_NVDLA_cbuf.scala 396:45:@4189.4]
  assign nv_ram_rws_28_io_ra = _T_95257_14_0; // @[NV_NVDLA_cbuf.scala 395:45:@4188.4]
  assign nv_ram_rws_28_io_wa = _T_13733_14_0; // @[NV_NVDLA_cbuf.scala 397:45:@4191.4]
  assign nv_ram_rws_28_io_di = _T_14845_14_0; // @[NV_NVDLA_cbuf.scala 398:45:@4192.4]
  assign nv_ram_rws_29_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4194.4]
  assign nv_ram_rws_29_io_re = _T_94145_14_1; // @[NV_NVDLA_cbuf.scala 394:45:@4195.4]
  assign nv_ram_rws_29_io_we = _T_16500_14_1; // @[NV_NVDLA_cbuf.scala 396:45:@4198.4]
  assign nv_ram_rws_29_io_ra = _T_95257_14_1; // @[NV_NVDLA_cbuf.scala 395:45:@4197.4]
  assign nv_ram_rws_29_io_wa = _T_13733_14_1; // @[NV_NVDLA_cbuf.scala 397:45:@4200.4]
  assign nv_ram_rws_29_io_di = _T_14845_14_1; // @[NV_NVDLA_cbuf.scala 398:45:@4201.4]
  assign nv_ram_rws_30_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4203.4]
  assign nv_ram_rws_30_io_re = _T_94145_15_0; // @[NV_NVDLA_cbuf.scala 394:45:@4204.4]
  assign nv_ram_rws_30_io_we = _T_16500_15_0; // @[NV_NVDLA_cbuf.scala 396:45:@4207.4]
  assign nv_ram_rws_30_io_ra = _T_95257_15_0; // @[NV_NVDLA_cbuf.scala 395:45:@4206.4]
  assign nv_ram_rws_30_io_wa = _T_13733_15_0; // @[NV_NVDLA_cbuf.scala 397:45:@4209.4]
  assign nv_ram_rws_30_io_di = _T_14845_15_0; // @[NV_NVDLA_cbuf.scala 398:45:@4210.4]
  assign nv_ram_rws_31_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_cbuf.scala 393:46:@4212.4]
  assign nv_ram_rws_31_io_re = _T_94145_15_1; // @[NV_NVDLA_cbuf.scala 394:45:@4213.4]
  assign nv_ram_rws_31_io_we = _T_16500_15_1; // @[NV_NVDLA_cbuf.scala 396:45:@4216.4]
  assign nv_ram_rws_31_io_ra = _T_95257_15_1; // @[NV_NVDLA_cbuf.scala 395:45:@4215.4]
  assign nv_ram_rws_31_io_wa = _T_13733_15_1; // @[NV_NVDLA_cbuf.scala 397:45:@4218.4]
  assign nv_ram_rws_31_io_di = _T_14845_15_1; // @[NV_NVDLA_cbuf.scala 398:45:@4219.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_7112_0_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_7112_0_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_7112_1_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_7112_1_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_7112_2_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_7112_2_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_7112_3_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_7112_3_1 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_7112_4_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_7112_4_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_7112_5_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_7112_5_1 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_7112_6_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_7112_6_1 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_7112_7_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_7112_7_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_7112_8_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_7112_8_1 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_7112_9_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_7112_9_1 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_7112_10_0 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_7112_10_1 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_7112_11_0 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_7112_11_1 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_7112_12_0 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_7112_12_1 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_7112_13_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_7112_13_1 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_7112_14_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_7112_14_1 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_7112_15_0 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_7112_15_1 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_8201_0 = _RAND_32[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_8201_1 = _RAND_33[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {8{`RANDOM}};
  _T_8215_0 = _RAND_34[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {8{`RANDOM}};
  _T_8215_1 = _RAND_35[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_9669_0_0 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_9669_0_1 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_9669_1_0 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_9669_1_1 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_9669_2_0 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_9669_2_1 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_9669_3_0 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_9669_3_1 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_9669_4_0 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_9669_4_1 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_9669_5_0 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_9669_5_1 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_9669_6_0 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_9669_6_1 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_9669_7_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_9669_7_1 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_9669_8_0 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_9669_8_1 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_9669_9_0 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_9669_9_1 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_9669_10_0 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_9669_10_1 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_9669_11_0 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_9669_11_1 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_9669_12_0 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_9669_12_1 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_9669_13_0 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_9669_13_1 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_9669_14_0 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_9669_14_1 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_9669_15_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_9669_15_1 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_13733_0_0 = _RAND_68[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_13733_0_1 = _RAND_69[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_13733_1_0 = _RAND_70[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_13733_1_1 = _RAND_71[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_13733_2_0 = _RAND_72[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_13733_2_1 = _RAND_73[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_13733_3_0 = _RAND_74[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_13733_3_1 = _RAND_75[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_13733_4_0 = _RAND_76[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_13733_4_1 = _RAND_77[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_13733_5_0 = _RAND_78[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_13733_5_1 = _RAND_79[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_13733_6_0 = _RAND_80[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_13733_6_1 = _RAND_81[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_13733_7_0 = _RAND_82[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_13733_7_1 = _RAND_83[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_13733_8_0 = _RAND_84[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_13733_8_1 = _RAND_85[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_13733_9_0 = _RAND_86[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_13733_9_1 = _RAND_87[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_13733_10_0 = _RAND_88[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_13733_10_1 = _RAND_89[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_13733_11_0 = _RAND_90[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_13733_11_1 = _RAND_91[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_13733_12_0 = _RAND_92[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_13733_12_1 = _RAND_93[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_13733_13_0 = _RAND_94[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_13733_13_1 = _RAND_95[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_13733_14_0 = _RAND_96[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_13733_14_1 = _RAND_97[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_13733_15_0 = _RAND_98[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_13733_15_1 = _RAND_99[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {8{`RANDOM}};
  _T_14845_0_0 = _RAND_100[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {8{`RANDOM}};
  _T_14845_0_1 = _RAND_101[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {8{`RANDOM}};
  _T_14845_1_0 = _RAND_102[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {8{`RANDOM}};
  _T_14845_1_1 = _RAND_103[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {8{`RANDOM}};
  _T_14845_2_0 = _RAND_104[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {8{`RANDOM}};
  _T_14845_2_1 = _RAND_105[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {8{`RANDOM}};
  _T_14845_3_0 = _RAND_106[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {8{`RANDOM}};
  _T_14845_3_1 = _RAND_107[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {8{`RANDOM}};
  _T_14845_4_0 = _RAND_108[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {8{`RANDOM}};
  _T_14845_4_1 = _RAND_109[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {8{`RANDOM}};
  _T_14845_5_0 = _RAND_110[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {8{`RANDOM}};
  _T_14845_5_1 = _RAND_111[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {8{`RANDOM}};
  _T_14845_6_0 = _RAND_112[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {8{`RANDOM}};
  _T_14845_6_1 = _RAND_113[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {8{`RANDOM}};
  _T_14845_7_0 = _RAND_114[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {8{`RANDOM}};
  _T_14845_7_1 = _RAND_115[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {8{`RANDOM}};
  _T_14845_8_0 = _RAND_116[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {8{`RANDOM}};
  _T_14845_8_1 = _RAND_117[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {8{`RANDOM}};
  _T_14845_9_0 = _RAND_118[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {8{`RANDOM}};
  _T_14845_9_1 = _RAND_119[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {8{`RANDOM}};
  _T_14845_10_0 = _RAND_120[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {8{`RANDOM}};
  _T_14845_10_1 = _RAND_121[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {8{`RANDOM}};
  _T_14845_11_0 = _RAND_122[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {8{`RANDOM}};
  _T_14845_11_1 = _RAND_123[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {8{`RANDOM}};
  _T_14845_12_0 = _RAND_124[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {8{`RANDOM}};
  _T_14845_12_1 = _RAND_125[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {8{`RANDOM}};
  _T_14845_13_0 = _RAND_126[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {8{`RANDOM}};
  _T_14845_13_1 = _RAND_127[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {8{`RANDOM}};
  _T_14845_14_0 = _RAND_128[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {8{`RANDOM}};
  _T_14845_14_1 = _RAND_129[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {8{`RANDOM}};
  _T_14845_15_0 = _RAND_130[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {8{`RANDOM}};
  _T_14845_15_1 = _RAND_131[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_16500_0_0 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_16500_0_1 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_16500_1_0 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_16500_1_1 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_16500_2_0 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_16500_2_1 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_16500_3_0 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_16500_3_1 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_16500_4_0 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_16500_4_1 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_16500_5_0 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_16500_5_1 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_16500_6_0 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_16500_6_1 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_16500_7_0 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_16500_7_1 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_16500_8_0 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_16500_8_1 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_16500_9_0 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_16500_9_1 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_16500_10_0 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_16500_10_1 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_16500_11_0 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_16500_11_1 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_16500_12_0 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_16500_12_1 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_16500_13_0 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_16500_13_1 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_16500_14_0 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_16500_14_1 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_16500_15_0 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_16500_15_1 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_39941_0_0_0 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_39941_0_1_0 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_39941_1_0_0 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_39941_1_1_0 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_39941_2_0_0 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_39941_2_1_0 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_39941_3_0_0 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_39941_3_1_0 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_39941_4_0_0 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_39941_4_1_0 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_39941_5_0_0 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_39941_5_1_0 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_39941_6_0_0 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_39941_6_1_0 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_39941_7_0_0 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_39941_7_1_0 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_39941_8_0_0 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_39941_8_1_0 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_39941_9_0_0 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_39941_9_1_0 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_39941_10_0_0 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_39941_10_1_0 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_39941_11_0_0 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_39941_11_1_0 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_39941_12_0_0 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_39941_12_1_0 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_39941_13_0_0 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_39941_13_1_0 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_39941_14_0_0 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_39941_14_1_0 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_39941_15_0_0 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_39941_15_1_0 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_72478_0_0_0 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_72478_0_1_0 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_72478_1_0_0 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_72478_1_1_0 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_72478_2_0_0 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_72478_2_1_0 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_72478_3_0_0 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_72478_3_1_0 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_72478_4_0_0 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_72478_4_1_0 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_72478_5_0_0 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_72478_5_1_0 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_72478_6_0_0 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_72478_6_1_0 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_72478_7_0_0 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_72478_7_1_0 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_72478_8_0_0 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_72478_8_1_0 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_72478_9_0_0 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_72478_9_1_0 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_72478_10_0_0 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_72478_10_1_0 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_72478_11_0_0 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_72478_11_1_0 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_72478_12_0_0 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_72478_12_1_0 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_72478_13_0_0 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_72478_13_1_0 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_72478_14_0_0 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_72478_14_1_0 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_72478_15_0_0 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_72478_15_1_0 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_86710 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_86712 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_86714 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_86716 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {16{`RANDOM}};
  _T_87674_0_0 = _RAND_232[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {16{`RANDOM}};
  _T_87674_1_0 = _RAND_233[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {16{`RANDOM}};
  _T_87674_2_0 = _RAND_234[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {16{`RANDOM}};
  _T_87674_3_0 = _RAND_235[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {16{`RANDOM}};
  _T_87674_4_0 = _RAND_236[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {16{`RANDOM}};
  _T_87674_5_0 = _RAND_237[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {16{`RANDOM}};
  _T_87674_6_0 = _RAND_238[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {16{`RANDOM}};
  _T_87674_7_0 = _RAND_239[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {16{`RANDOM}};
  _T_87674_8_0 = _RAND_240[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {16{`RANDOM}};
  _T_87674_9_0 = _RAND_241[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {16{`RANDOM}};
  _T_87674_10_0 = _RAND_242[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {16{`RANDOM}};
  _T_87674_11_0 = _RAND_243[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {16{`RANDOM}};
  _T_87674_12_0 = _RAND_244[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {16{`RANDOM}};
  _T_87674_13_0 = _RAND_245[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {16{`RANDOM}};
  _T_87674_14_0 = _RAND_246[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {16{`RANDOM}};
  _T_87674_15_0 = _RAND_247[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {16{`RANDOM}};
  _T_88155_0_0 = _RAND_248[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {16{`RANDOM}};
  _T_88155_1_0 = _RAND_249[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {16{`RANDOM}};
  _T_88155_2_0 = _RAND_250[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {16{`RANDOM}};
  _T_88155_3_0 = _RAND_251[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {16{`RANDOM}};
  _T_88225_0_0 = _RAND_252[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {16{`RANDOM}};
  _T_88249 = _RAND_253[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_89522_0_0 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_89522_0_1 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_89522_1_0 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_89522_1_1 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_89522_2_0 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_89522_2_1 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_89522_3_0 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_89522_3_1 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_89522_4_0 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_89522_4_1 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_89522_5_0 = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_89522_5_1 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_89522_6_0 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_89522_6_1 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_89522_7_0 = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_89522_7_1 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_89522_8_0 = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_89522_8_1 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_89522_9_0 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_89522_9_1 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_89522_10_0 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_89522_10_1 = _RAND_275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_89522_11_0 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_89522_11_1 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_89522_12_0 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_89522_12_1 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_89522_13_0 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_89522_13_1 = _RAND_281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_89522_14_0 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_89522_14_1 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_89522_15_0 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_89522_15_1 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_91073_0_0 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_91073_0_1 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_91073_1_0 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_91073_1_1 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_91073_2_0 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_91073_2_1 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_91073_3_0 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_91073_3_1 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_91073_4_0 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_91073_4_1 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_91073_5_0 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_91073_5_1 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_91073_6_0 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_91073_6_1 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_91073_7_0 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_91073_7_1 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_91073_8_0 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_91073_8_1 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_91073_9_0 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_91073_9_1 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_91073_10_0 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_91073_10_1 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_91073_11_0 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_91073_11_1 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_91073_12_0 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_91073_12_1 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_91073_13_0 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_91073_13_1 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_91073_14_0 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_91073_14_1 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_91073_15_0 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_91073_15_1 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_92368 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_92370 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_92372 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_92374 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {16{`RANDOM}};
  _T_92609_0 = _RAND_322[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {16{`RANDOM}};
  _T_92609_1 = _RAND_323[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {16{`RANDOM}};
  _T_92609_2 = _RAND_324[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {16{`RANDOM}};
  _T_92609_3 = _RAND_325[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {16{`RANDOM}};
  _T_92609_4 = _RAND_326[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {16{`RANDOM}};
  _T_92609_5 = _RAND_327[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {16{`RANDOM}};
  _T_92609_6 = _RAND_328[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {16{`RANDOM}};
  _T_92609_7 = _RAND_329[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {16{`RANDOM}};
  _T_92609_8 = _RAND_330[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {16{`RANDOM}};
  _T_92609_9 = _RAND_331[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {16{`RANDOM}};
  _T_92609_10 = _RAND_332[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {16{`RANDOM}};
  _T_92609_11 = _RAND_333[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {16{`RANDOM}};
  _T_92609_12 = _RAND_334[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {16{`RANDOM}};
  _T_92609_13 = _RAND_335[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {16{`RANDOM}};
  _T_92609_14 = _RAND_336[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {16{`RANDOM}};
  _T_92609_15 = _RAND_337[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {16{`RANDOM}};
  _T_92665_0 = _RAND_338[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {16{`RANDOM}};
  _T_92665_1 = _RAND_339[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {16{`RANDOM}};
  _T_92665_2 = _RAND_340[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {16{`RANDOM}};
  _T_92665_3 = _RAND_341[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {16{`RANDOM}};
  _T_92687_0 = _RAND_342[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {16{`RANDOM}};
  _T_92695 = _RAND_343[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_94145_0_0 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_94145_0_1 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_94145_1_0 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_94145_1_1 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_94145_2_0 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_94145_2_1 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_94145_3_0 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_94145_3_1 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_94145_4_0 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_94145_4_1 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_94145_5_0 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_94145_5_1 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_94145_6_0 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_94145_6_1 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_94145_7_0 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_94145_7_1 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_94145_8_0 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_94145_8_1 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_94145_9_0 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_94145_9_1 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_94145_10_0 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_94145_10_1 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_94145_11_0 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_94145_11_1 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_94145_12_0 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_94145_12_1 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_94145_13_0 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_94145_13_1 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_94145_14_0 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_94145_14_1 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_94145_15_0 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_94145_15_1 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_95257_0_0 = _RAND_376[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_95257_0_1 = _RAND_377[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_95257_1_0 = _RAND_378[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_95257_1_1 = _RAND_379[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_95257_2_0 = _RAND_380[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_95257_2_1 = _RAND_381[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_95257_3_0 = _RAND_382[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_95257_3_1 = _RAND_383[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_95257_4_0 = _RAND_384[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_95257_4_1 = _RAND_385[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_95257_5_0 = _RAND_386[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_95257_5_1 = _RAND_387[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_95257_6_0 = _RAND_388[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_95257_6_1 = _RAND_389[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_95257_7_0 = _RAND_390[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_95257_7_1 = _RAND_391[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_95257_8_0 = _RAND_392[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_95257_8_1 = _RAND_393[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_95257_9_0 = _RAND_394[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_95257_9_1 = _RAND_395[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_95257_10_0 = _RAND_396[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_95257_10_1 = _RAND_397[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_95257_11_0 = _RAND_398[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_95257_11_1 = _RAND_399[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_95257_12_0 = _RAND_400[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_95257_12_1 = _RAND_401[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_95257_13_0 = _RAND_402[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_95257_13_1 = _RAND_403[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_95257_14_0 = _RAND_404[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_95257_14_1 = _RAND_405[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_95257_15_0 = _RAND_406[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_95257_15_1 = _RAND_407[8:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (_T_178) begin
      _T_7112_0_0 <= 1'h0;
    end else begin
      _T_7112_0_0 <= _T_8151;
    end
    if (_T_178) begin
      _T_7112_0_1 <= 1'h0;
    end else begin
      _T_7112_0_1 <= _T_8152;
    end
    if (_T_178) begin
      _T_7112_1_0 <= 1'h0;
    end else begin
      _T_7112_1_0 <= _T_8153;
    end
    if (_T_178) begin
      _T_7112_1_1 <= 1'h0;
    end else begin
      _T_7112_1_1 <= _T_8154;
    end
    if (_T_178) begin
      _T_7112_2_0 <= 1'h0;
    end else begin
      _T_7112_2_0 <= _T_8155;
    end
    if (_T_178) begin
      _T_7112_2_1 <= 1'h0;
    end else begin
      _T_7112_2_1 <= _T_8156;
    end
    if (_T_178) begin
      _T_7112_3_0 <= 1'h0;
    end else begin
      _T_7112_3_0 <= _T_8157;
    end
    if (_T_178) begin
      _T_7112_3_1 <= 1'h0;
    end else begin
      _T_7112_3_1 <= _T_8158;
    end
    if (_T_178) begin
      _T_7112_4_0 <= 1'h0;
    end else begin
      _T_7112_4_0 <= _T_8159;
    end
    if (_T_178) begin
      _T_7112_4_1 <= 1'h0;
    end else begin
      _T_7112_4_1 <= _T_8160;
    end
    if (_T_178) begin
      _T_7112_5_0 <= 1'h0;
    end else begin
      _T_7112_5_0 <= _T_8161;
    end
    if (_T_178) begin
      _T_7112_5_1 <= 1'h0;
    end else begin
      _T_7112_5_1 <= _T_8162;
    end
    if (_T_178) begin
      _T_7112_6_0 <= 1'h0;
    end else begin
      _T_7112_6_0 <= _T_8163;
    end
    if (_T_178) begin
      _T_7112_6_1 <= 1'h0;
    end else begin
      _T_7112_6_1 <= _T_8164;
    end
    if (_T_178) begin
      _T_7112_7_0 <= 1'h0;
    end else begin
      _T_7112_7_0 <= _T_8165;
    end
    if (_T_178) begin
      _T_7112_7_1 <= 1'h0;
    end else begin
      _T_7112_7_1 <= _T_8166;
    end
    if (_T_178) begin
      _T_7112_8_0 <= 1'h0;
    end else begin
      _T_7112_8_0 <= _T_8167;
    end
    if (_T_178) begin
      _T_7112_8_1 <= 1'h0;
    end else begin
      _T_7112_8_1 <= _T_8168;
    end
    if (_T_178) begin
      _T_7112_9_0 <= 1'h0;
    end else begin
      _T_7112_9_0 <= _T_8169;
    end
    if (_T_178) begin
      _T_7112_9_1 <= 1'h0;
    end else begin
      _T_7112_9_1 <= _T_8170;
    end
    if (_T_178) begin
      _T_7112_10_0 <= 1'h0;
    end else begin
      _T_7112_10_0 <= _T_8171;
    end
    if (_T_178) begin
      _T_7112_10_1 <= 1'h0;
    end else begin
      _T_7112_10_1 <= _T_8172;
    end
    if (_T_178) begin
      _T_7112_11_0 <= 1'h0;
    end else begin
      _T_7112_11_0 <= _T_8173;
    end
    if (_T_178) begin
      _T_7112_11_1 <= 1'h0;
    end else begin
      _T_7112_11_1 <= _T_8174;
    end
    if (_T_178) begin
      _T_7112_12_0 <= 1'h0;
    end else begin
      _T_7112_12_0 <= _T_8175;
    end
    if (_T_178) begin
      _T_7112_12_1 <= 1'h0;
    end else begin
      _T_7112_12_1 <= _T_8176;
    end
    if (_T_178) begin
      _T_7112_13_0 <= 1'h0;
    end else begin
      _T_7112_13_0 <= _T_8177;
    end
    if (_T_178) begin
      _T_7112_13_1 <= 1'h0;
    end else begin
      _T_7112_13_1 <= _T_8178;
    end
    if (_T_178) begin
      _T_7112_14_0 <= 1'h0;
    end else begin
      _T_7112_14_0 <= _T_8179;
    end
    if (_T_178) begin
      _T_7112_14_1 <= 1'h0;
    end else begin
      _T_7112_14_1 <= _T_8180;
    end
    if (_T_178) begin
      _T_7112_15_0 <= 1'h0;
    end else begin
      _T_7112_15_0 <= _T_8181;
    end
    if (_T_178) begin
      _T_7112_15_1 <= 1'h0;
    end else begin
      _T_7112_15_1 <= _T_8182;
    end
    if (_T_178) begin
      _T_8201_0 <= 13'h0;
    end else begin
      _T_8201_0 <= io_cdma2buf_wr_addr_0;
    end
    if (_T_178) begin
      _T_8201_1 <= 13'h0;
    end else begin
      _T_8201_1 <= io_cdma2buf_wr_addr_1;
    end
    _T_8215_0 <= io_cdma2buf_wr_data_0;
    _T_8215_1 <= io_cdma2buf_wr_data_1;
    if (_T_178) begin
      _T_9669_0_0 <= 1'h0;
    end else begin
      _T_9669_0_0 <= _T_10708;
    end
    if (_T_178) begin
      _T_9669_0_1 <= 1'h0;
    end else begin
      _T_9669_0_1 <= _T_10724;
    end
    if (_T_178) begin
      _T_9669_1_0 <= 1'h0;
    end else begin
      _T_9669_1_0 <= _T_10709;
    end
    if (_T_178) begin
      _T_9669_1_1 <= 1'h0;
    end else begin
      _T_9669_1_1 <= _T_10725;
    end
    if (_T_178) begin
      _T_9669_2_0 <= 1'h0;
    end else begin
      _T_9669_2_0 <= _T_10710;
    end
    if (_T_178) begin
      _T_9669_2_1 <= 1'h0;
    end else begin
      _T_9669_2_1 <= _T_10726;
    end
    if (_T_178) begin
      _T_9669_3_0 <= 1'h0;
    end else begin
      _T_9669_3_0 <= _T_10711;
    end
    if (_T_178) begin
      _T_9669_3_1 <= 1'h0;
    end else begin
      _T_9669_3_1 <= _T_10727;
    end
    if (_T_178) begin
      _T_9669_4_0 <= 1'h0;
    end else begin
      _T_9669_4_0 <= _T_10712;
    end
    if (_T_178) begin
      _T_9669_4_1 <= 1'h0;
    end else begin
      _T_9669_4_1 <= _T_10728;
    end
    if (_T_178) begin
      _T_9669_5_0 <= 1'h0;
    end else begin
      _T_9669_5_0 <= _T_10713;
    end
    if (_T_178) begin
      _T_9669_5_1 <= 1'h0;
    end else begin
      _T_9669_5_1 <= _T_10729;
    end
    if (_T_178) begin
      _T_9669_6_0 <= 1'h0;
    end else begin
      _T_9669_6_0 <= _T_10714;
    end
    if (_T_178) begin
      _T_9669_6_1 <= 1'h0;
    end else begin
      _T_9669_6_1 <= _T_10730;
    end
    if (_T_178) begin
      _T_9669_7_0 <= 1'h0;
    end else begin
      _T_9669_7_0 <= _T_10715;
    end
    if (_T_178) begin
      _T_9669_7_1 <= 1'h0;
    end else begin
      _T_9669_7_1 <= _T_10731;
    end
    if (_T_178) begin
      _T_9669_8_0 <= 1'h0;
    end else begin
      _T_9669_8_0 <= _T_10716;
    end
    if (_T_178) begin
      _T_9669_8_1 <= 1'h0;
    end else begin
      _T_9669_8_1 <= _T_10732;
    end
    if (_T_178) begin
      _T_9669_9_0 <= 1'h0;
    end else begin
      _T_9669_9_0 <= _T_10717;
    end
    if (_T_178) begin
      _T_9669_9_1 <= 1'h0;
    end else begin
      _T_9669_9_1 <= _T_10733;
    end
    if (_T_178) begin
      _T_9669_10_0 <= 1'h0;
    end else begin
      _T_9669_10_0 <= _T_10718;
    end
    if (_T_178) begin
      _T_9669_10_1 <= 1'h0;
    end else begin
      _T_9669_10_1 <= _T_10734;
    end
    if (_T_178) begin
      _T_9669_11_0 <= 1'h0;
    end else begin
      _T_9669_11_0 <= _T_10719;
    end
    if (_T_178) begin
      _T_9669_11_1 <= 1'h0;
    end else begin
      _T_9669_11_1 <= _T_10735;
    end
    if (_T_178) begin
      _T_9669_12_0 <= 1'h0;
    end else begin
      _T_9669_12_0 <= _T_10720;
    end
    if (_T_178) begin
      _T_9669_12_1 <= 1'h0;
    end else begin
      _T_9669_12_1 <= _T_10736;
    end
    if (_T_178) begin
      _T_9669_13_0 <= 1'h0;
    end else begin
      _T_9669_13_0 <= _T_10721;
    end
    if (_T_178) begin
      _T_9669_13_1 <= 1'h0;
    end else begin
      _T_9669_13_1 <= _T_10737;
    end
    if (_T_178) begin
      _T_9669_14_0 <= 1'h0;
    end else begin
      _T_9669_14_0 <= _T_10722;
    end
    if (_T_178) begin
      _T_9669_14_1 <= 1'h0;
    end else begin
      _T_9669_14_1 <= _T_10738;
    end
    if (_T_178) begin
      _T_9669_15_0 <= 1'h0;
    end else begin
      _T_9669_15_0 <= _T_10723;
    end
    if (_T_178) begin
      _T_9669_15_1 <= 1'h0;
    end else begin
      _T_9669_15_1 <= _T_10739;
    end
    if (_T_178) begin
      _T_13733_0_0 <= 9'h0;
    end else begin
      _T_13733_0_0 <= _T_12252;
    end
    if (_T_178) begin
      _T_13733_0_1 <= 9'h0;
    end else begin
      _T_13733_0_1 <= _T_12252;
    end
    if (_T_178) begin
      _T_13733_1_0 <= 9'h0;
    end else begin
      _T_13733_1_0 <= _T_12254;
    end
    if (_T_178) begin
      _T_13733_1_1 <= 9'h0;
    end else begin
      _T_13733_1_1 <= _T_12254;
    end
    if (_T_178) begin
      _T_13733_2_0 <= 9'h0;
    end else begin
      _T_13733_2_0 <= _T_12256;
    end
    if (_T_178) begin
      _T_13733_2_1 <= 9'h0;
    end else begin
      _T_13733_2_1 <= _T_12256;
    end
    if (_T_178) begin
      _T_13733_3_0 <= 9'h0;
    end else begin
      _T_13733_3_0 <= _T_12258;
    end
    if (_T_178) begin
      _T_13733_3_1 <= 9'h0;
    end else begin
      _T_13733_3_1 <= _T_12258;
    end
    if (_T_178) begin
      _T_13733_4_0 <= 9'h0;
    end else begin
      _T_13733_4_0 <= _T_12260;
    end
    if (_T_178) begin
      _T_13733_4_1 <= 9'h0;
    end else begin
      _T_13733_4_1 <= _T_12260;
    end
    if (_T_178) begin
      _T_13733_5_0 <= 9'h0;
    end else begin
      _T_13733_5_0 <= _T_12262;
    end
    if (_T_178) begin
      _T_13733_5_1 <= 9'h0;
    end else begin
      _T_13733_5_1 <= _T_12262;
    end
    if (_T_178) begin
      _T_13733_6_0 <= 9'h0;
    end else begin
      _T_13733_6_0 <= _T_12264;
    end
    if (_T_178) begin
      _T_13733_6_1 <= 9'h0;
    end else begin
      _T_13733_6_1 <= _T_12264;
    end
    if (_T_178) begin
      _T_13733_7_0 <= 9'h0;
    end else begin
      _T_13733_7_0 <= _T_12266;
    end
    if (_T_178) begin
      _T_13733_7_1 <= 9'h0;
    end else begin
      _T_13733_7_1 <= _T_12266;
    end
    if (_T_178) begin
      _T_13733_8_0 <= 9'h0;
    end else begin
      _T_13733_8_0 <= _T_12268;
    end
    if (_T_178) begin
      _T_13733_8_1 <= 9'h0;
    end else begin
      _T_13733_8_1 <= _T_12268;
    end
    if (_T_178) begin
      _T_13733_9_0 <= 9'h0;
    end else begin
      _T_13733_9_0 <= _T_12270;
    end
    if (_T_178) begin
      _T_13733_9_1 <= 9'h0;
    end else begin
      _T_13733_9_1 <= _T_12270;
    end
    if (_T_178) begin
      _T_13733_10_0 <= 9'h0;
    end else begin
      _T_13733_10_0 <= _T_12272;
    end
    if (_T_178) begin
      _T_13733_10_1 <= 9'h0;
    end else begin
      _T_13733_10_1 <= _T_12272;
    end
    if (_T_178) begin
      _T_13733_11_0 <= 9'h0;
    end else begin
      _T_13733_11_0 <= _T_12274;
    end
    if (_T_178) begin
      _T_13733_11_1 <= 9'h0;
    end else begin
      _T_13733_11_1 <= _T_12274;
    end
    if (_T_178) begin
      _T_13733_12_0 <= 9'h0;
    end else begin
      _T_13733_12_0 <= _T_12276;
    end
    if (_T_178) begin
      _T_13733_12_1 <= 9'h0;
    end else begin
      _T_13733_12_1 <= _T_12276;
    end
    if (_T_178) begin
      _T_13733_13_0 <= 9'h0;
    end else begin
      _T_13733_13_0 <= _T_12278;
    end
    if (_T_178) begin
      _T_13733_13_1 <= 9'h0;
    end else begin
      _T_13733_13_1 <= _T_12278;
    end
    if (_T_178) begin
      _T_13733_14_0 <= 9'h0;
    end else begin
      _T_13733_14_0 <= _T_12280;
    end
    if (_T_178) begin
      _T_13733_14_1 <= 9'h0;
    end else begin
      _T_13733_14_1 <= _T_12280;
    end
    if (_T_178) begin
      _T_13733_15_0 <= 9'h0;
    end else begin
      _T_13733_15_0 <= _T_12282;
    end
    if (_T_178) begin
      _T_13733_15_1 <= 9'h0;
    end else begin
      _T_13733_15_1 <= _T_12282;
    end
    _T_14845_0_0 <= _T_11351 | _T_11361;
    _T_14845_0_1 <= _T_11351 | _T_11361;
    _T_14845_1_0 <= _T_11373 | _T_11383;
    _T_14845_1_1 <= _T_11373 | _T_11383;
    _T_14845_2_0 <= _T_11395 | _T_11405;
    _T_14845_2_1 <= _T_11395 | _T_11405;
    _T_14845_3_0 <= _T_11417 | _T_11427;
    _T_14845_3_1 <= _T_11417 | _T_11427;
    _T_14845_4_0 <= _T_11439 | _T_11449;
    _T_14845_4_1 <= _T_11439 | _T_11449;
    _T_14845_5_0 <= _T_11461 | _T_11471;
    _T_14845_5_1 <= _T_11461 | _T_11471;
    _T_14845_6_0 <= _T_11483 | _T_11493;
    _T_14845_6_1 <= _T_11483 | _T_11493;
    _T_14845_7_0 <= _T_11505 | _T_11515;
    _T_14845_7_1 <= _T_11505 | _T_11515;
    _T_14845_8_0 <= _T_11527 | _T_11537;
    _T_14845_8_1 <= _T_11527 | _T_11537;
    _T_14845_9_0 <= _T_11549 | _T_11559;
    _T_14845_9_1 <= _T_11549 | _T_11559;
    _T_14845_10_0 <= _T_11571 | _T_11581;
    _T_14845_10_1 <= _T_11571 | _T_11581;
    _T_14845_11_0 <= _T_11593 | _T_11603;
    _T_14845_11_1 <= _T_11593 | _T_11603;
    _T_14845_12_0 <= _T_11615 | _T_11625;
    _T_14845_12_1 <= _T_11615 | _T_11625;
    _T_14845_13_0 <= _T_11637 | _T_11647;
    _T_14845_13_1 <= _T_11637 | _T_11647;
    _T_14845_14_0 <= _T_11659 | _T_11669;
    _T_14845_14_1 <= _T_11659 | _T_11669;
    _T_14845_15_0 <= _T_11681 | _T_11691;
    _T_14845_15_1 <= _T_11681 | _T_11691;
    if (_T_178) begin
      _T_16500_0_0 <= 1'h0;
    end else begin
      _T_16500_0_0 <= _T_7112_0_0;
    end
    if (_T_178) begin
      _T_16500_0_1 <= 1'h0;
    end else begin
      _T_16500_0_1 <= _T_7112_0_1;
    end
    if (_T_178) begin
      _T_16500_1_0 <= 1'h0;
    end else begin
      _T_16500_1_0 <= _T_7112_1_0;
    end
    if (_T_178) begin
      _T_16500_1_1 <= 1'h0;
    end else begin
      _T_16500_1_1 <= _T_7112_1_1;
    end
    if (_T_178) begin
      _T_16500_2_0 <= 1'h0;
    end else begin
      _T_16500_2_0 <= _T_7112_2_0;
    end
    if (_T_178) begin
      _T_16500_2_1 <= 1'h0;
    end else begin
      _T_16500_2_1 <= _T_7112_2_1;
    end
    if (_T_178) begin
      _T_16500_3_0 <= 1'h0;
    end else begin
      _T_16500_3_0 <= _T_7112_3_0;
    end
    if (_T_178) begin
      _T_16500_3_1 <= 1'h0;
    end else begin
      _T_16500_3_1 <= _T_7112_3_1;
    end
    if (_T_178) begin
      _T_16500_4_0 <= 1'h0;
    end else begin
      _T_16500_4_0 <= _T_7112_4_0;
    end
    if (_T_178) begin
      _T_16500_4_1 <= 1'h0;
    end else begin
      _T_16500_4_1 <= _T_7112_4_1;
    end
    if (_T_178) begin
      _T_16500_5_0 <= 1'h0;
    end else begin
      _T_16500_5_0 <= _T_7112_5_0;
    end
    if (_T_178) begin
      _T_16500_5_1 <= 1'h0;
    end else begin
      _T_16500_5_1 <= _T_7112_5_1;
    end
    if (_T_178) begin
      _T_16500_6_0 <= 1'h0;
    end else begin
      _T_16500_6_0 <= _T_7112_6_0;
    end
    if (_T_178) begin
      _T_16500_6_1 <= 1'h0;
    end else begin
      _T_16500_6_1 <= _T_7112_6_1;
    end
    if (_T_178) begin
      _T_16500_7_0 <= 1'h0;
    end else begin
      _T_16500_7_0 <= _T_7112_7_0;
    end
    if (_T_178) begin
      _T_16500_7_1 <= 1'h0;
    end else begin
      _T_16500_7_1 <= _T_7112_7_1;
    end
    if (_T_178) begin
      _T_16500_8_0 <= 1'h0;
    end else begin
      _T_16500_8_0 <= _T_7112_8_0;
    end
    if (_T_178) begin
      _T_16500_8_1 <= 1'h0;
    end else begin
      _T_16500_8_1 <= _T_7112_8_1;
    end
    if (_T_178) begin
      _T_16500_9_0 <= 1'h0;
    end else begin
      _T_16500_9_0 <= _T_7112_9_0;
    end
    if (_T_178) begin
      _T_16500_9_1 <= 1'h0;
    end else begin
      _T_16500_9_1 <= _T_7112_9_1;
    end
    if (_T_178) begin
      _T_16500_10_0 <= 1'h0;
    end else begin
      _T_16500_10_0 <= _T_7112_10_0;
    end
    if (_T_178) begin
      _T_16500_10_1 <= 1'h0;
    end else begin
      _T_16500_10_1 <= _T_7112_10_1;
    end
    if (_T_178) begin
      _T_16500_11_0 <= 1'h0;
    end else begin
      _T_16500_11_0 <= _T_7112_11_0;
    end
    if (_T_178) begin
      _T_16500_11_1 <= 1'h0;
    end else begin
      _T_16500_11_1 <= _T_7112_11_1;
    end
    if (_T_178) begin
      _T_16500_12_0 <= 1'h0;
    end else begin
      _T_16500_12_0 <= _T_7112_12_0;
    end
    if (_T_178) begin
      _T_16500_12_1 <= 1'h0;
    end else begin
      _T_16500_12_1 <= _T_7112_12_1;
    end
    if (_T_178) begin
      _T_16500_13_0 <= 1'h0;
    end else begin
      _T_16500_13_0 <= _T_7112_13_0;
    end
    if (_T_178) begin
      _T_16500_13_1 <= 1'h0;
    end else begin
      _T_16500_13_1 <= _T_7112_13_1;
    end
    if (_T_178) begin
      _T_16500_14_0 <= 1'h0;
    end else begin
      _T_16500_14_0 <= _T_7112_14_0;
    end
    if (_T_178) begin
      _T_16500_14_1 <= 1'h0;
    end else begin
      _T_16500_14_1 <= _T_7112_14_1;
    end
    if (_T_178) begin
      _T_16500_15_0 <= 1'h0;
    end else begin
      _T_16500_15_0 <= _T_7112_15_0;
    end
    if (_T_178) begin
      _T_16500_15_1 <= 1'h0;
    end else begin
      _T_16500_15_1 <= _T_7112_15_1;
    end
    if (_T_178) begin
      _T_39941_0_0_0 <= 1'h0;
    end else begin
      _T_39941_0_0_0 <= _T_19413;
    end
    if (_T_178) begin
      _T_39941_0_1_0 <= 1'h0;
    end else begin
      _T_39941_0_1_0 <= _T_19413;
    end
    if (_T_178) begin
      _T_39941_1_0_0 <= 1'h0;
    end else begin
      _T_39941_1_0_0 <= _T_19421;
    end
    if (_T_178) begin
      _T_39941_1_1_0 <= 1'h0;
    end else begin
      _T_39941_1_1_0 <= _T_19421;
    end
    if (_T_178) begin
      _T_39941_2_0_0 <= 1'h0;
    end else begin
      _T_39941_2_0_0 <= _T_19429;
    end
    if (_T_178) begin
      _T_39941_2_1_0 <= 1'h0;
    end else begin
      _T_39941_2_1_0 <= _T_19429;
    end
    if (_T_178) begin
      _T_39941_3_0_0 <= 1'h0;
    end else begin
      _T_39941_3_0_0 <= _T_19437;
    end
    if (_T_178) begin
      _T_39941_3_1_0 <= 1'h0;
    end else begin
      _T_39941_3_1_0 <= _T_19437;
    end
    if (_T_178) begin
      _T_39941_4_0_0 <= 1'h0;
    end else begin
      _T_39941_4_0_0 <= _T_19445;
    end
    if (_T_178) begin
      _T_39941_4_1_0 <= 1'h0;
    end else begin
      _T_39941_4_1_0 <= _T_19445;
    end
    if (_T_178) begin
      _T_39941_5_0_0 <= 1'h0;
    end else begin
      _T_39941_5_0_0 <= _T_19453;
    end
    if (_T_178) begin
      _T_39941_5_1_0 <= 1'h0;
    end else begin
      _T_39941_5_1_0 <= _T_19453;
    end
    if (_T_178) begin
      _T_39941_6_0_0 <= 1'h0;
    end else begin
      _T_39941_6_0_0 <= _T_19461;
    end
    if (_T_178) begin
      _T_39941_6_1_0 <= 1'h0;
    end else begin
      _T_39941_6_1_0 <= _T_19461;
    end
    if (_T_178) begin
      _T_39941_7_0_0 <= 1'h0;
    end else begin
      _T_39941_7_0_0 <= _T_19469;
    end
    if (_T_178) begin
      _T_39941_7_1_0 <= 1'h0;
    end else begin
      _T_39941_7_1_0 <= _T_19469;
    end
    if (_T_178) begin
      _T_39941_8_0_0 <= 1'h0;
    end else begin
      _T_39941_8_0_0 <= _T_19477;
    end
    if (_T_178) begin
      _T_39941_8_1_0 <= 1'h0;
    end else begin
      _T_39941_8_1_0 <= _T_19477;
    end
    if (_T_178) begin
      _T_39941_9_0_0 <= 1'h0;
    end else begin
      _T_39941_9_0_0 <= _T_19485;
    end
    if (_T_178) begin
      _T_39941_9_1_0 <= 1'h0;
    end else begin
      _T_39941_9_1_0 <= _T_19485;
    end
    if (_T_178) begin
      _T_39941_10_0_0 <= 1'h0;
    end else begin
      _T_39941_10_0_0 <= _T_19493;
    end
    if (_T_178) begin
      _T_39941_10_1_0 <= 1'h0;
    end else begin
      _T_39941_10_1_0 <= _T_19493;
    end
    if (_T_178) begin
      _T_39941_11_0_0 <= 1'h0;
    end else begin
      _T_39941_11_0_0 <= _T_19501;
    end
    if (_T_178) begin
      _T_39941_11_1_0 <= 1'h0;
    end else begin
      _T_39941_11_1_0 <= _T_19501;
    end
    if (_T_178) begin
      _T_39941_12_0_0 <= 1'h0;
    end else begin
      _T_39941_12_0_0 <= _T_19509;
    end
    if (_T_178) begin
      _T_39941_12_1_0 <= 1'h0;
    end else begin
      _T_39941_12_1_0 <= _T_19509;
    end
    if (_T_178) begin
      _T_39941_13_0_0 <= 1'h0;
    end else begin
      _T_39941_13_0_0 <= _T_19517;
    end
    if (_T_178) begin
      _T_39941_13_1_0 <= 1'h0;
    end else begin
      _T_39941_13_1_0 <= _T_19517;
    end
    if (_T_178) begin
      _T_39941_14_0_0 <= 1'h0;
    end else begin
      _T_39941_14_0_0 <= _T_19525;
    end
    if (_T_178) begin
      _T_39941_14_1_0 <= 1'h0;
    end else begin
      _T_39941_14_1_0 <= _T_19525;
    end
    if (_T_178) begin
      _T_39941_15_0_0 <= 1'h0;
    end else begin
      _T_39941_15_0_0 <= _T_19533;
    end
    if (_T_178) begin
      _T_39941_15_1_0 <= 1'h0;
    end else begin
      _T_39941_15_1_0 <= _T_19533;
    end
    if (_T_178) begin
      _T_72478_0_0_0 <= 1'h0;
    end else begin
      _T_72478_0_0_0 <= _T_39941_0_0_0;
    end
    if (_T_178) begin
      _T_72478_0_1_0 <= 1'h0;
    end else begin
      _T_72478_0_1_0 <= _T_39941_0_1_0;
    end
    if (_T_178) begin
      _T_72478_1_0_0 <= 1'h0;
    end else begin
      _T_72478_1_0_0 <= _T_39941_1_0_0;
    end
    if (_T_178) begin
      _T_72478_1_1_0 <= 1'h0;
    end else begin
      _T_72478_1_1_0 <= _T_39941_1_1_0;
    end
    if (_T_178) begin
      _T_72478_2_0_0 <= 1'h0;
    end else begin
      _T_72478_2_0_0 <= _T_39941_2_0_0;
    end
    if (_T_178) begin
      _T_72478_2_1_0 <= 1'h0;
    end else begin
      _T_72478_2_1_0 <= _T_39941_2_1_0;
    end
    if (_T_178) begin
      _T_72478_3_0_0 <= 1'h0;
    end else begin
      _T_72478_3_0_0 <= _T_39941_3_0_0;
    end
    if (_T_178) begin
      _T_72478_3_1_0 <= 1'h0;
    end else begin
      _T_72478_3_1_0 <= _T_39941_3_1_0;
    end
    if (_T_178) begin
      _T_72478_4_0_0 <= 1'h0;
    end else begin
      _T_72478_4_0_0 <= _T_39941_4_0_0;
    end
    if (_T_178) begin
      _T_72478_4_1_0 <= 1'h0;
    end else begin
      _T_72478_4_1_0 <= _T_39941_4_1_0;
    end
    if (_T_178) begin
      _T_72478_5_0_0 <= 1'h0;
    end else begin
      _T_72478_5_0_0 <= _T_39941_5_0_0;
    end
    if (_T_178) begin
      _T_72478_5_1_0 <= 1'h0;
    end else begin
      _T_72478_5_1_0 <= _T_39941_5_1_0;
    end
    if (_T_178) begin
      _T_72478_6_0_0 <= 1'h0;
    end else begin
      _T_72478_6_0_0 <= _T_39941_6_0_0;
    end
    if (_T_178) begin
      _T_72478_6_1_0 <= 1'h0;
    end else begin
      _T_72478_6_1_0 <= _T_39941_6_1_0;
    end
    if (_T_178) begin
      _T_72478_7_0_0 <= 1'h0;
    end else begin
      _T_72478_7_0_0 <= _T_39941_7_0_0;
    end
    if (_T_178) begin
      _T_72478_7_1_0 <= 1'h0;
    end else begin
      _T_72478_7_1_0 <= _T_39941_7_1_0;
    end
    if (_T_178) begin
      _T_72478_8_0_0 <= 1'h0;
    end else begin
      _T_72478_8_0_0 <= _T_39941_8_0_0;
    end
    if (_T_178) begin
      _T_72478_8_1_0 <= 1'h0;
    end else begin
      _T_72478_8_1_0 <= _T_39941_8_1_0;
    end
    if (_T_178) begin
      _T_72478_9_0_0 <= 1'h0;
    end else begin
      _T_72478_9_0_0 <= _T_39941_9_0_0;
    end
    if (_T_178) begin
      _T_72478_9_1_0 <= 1'h0;
    end else begin
      _T_72478_9_1_0 <= _T_39941_9_1_0;
    end
    if (_T_178) begin
      _T_72478_10_0_0 <= 1'h0;
    end else begin
      _T_72478_10_0_0 <= _T_39941_10_0_0;
    end
    if (_T_178) begin
      _T_72478_10_1_0 <= 1'h0;
    end else begin
      _T_72478_10_1_0 <= _T_39941_10_1_0;
    end
    if (_T_178) begin
      _T_72478_11_0_0 <= 1'h0;
    end else begin
      _T_72478_11_0_0 <= _T_39941_11_0_0;
    end
    if (_T_178) begin
      _T_72478_11_1_0 <= 1'h0;
    end else begin
      _T_72478_11_1_0 <= _T_39941_11_1_0;
    end
    if (_T_178) begin
      _T_72478_12_0_0 <= 1'h0;
    end else begin
      _T_72478_12_0_0 <= _T_39941_12_0_0;
    end
    if (_T_178) begin
      _T_72478_12_1_0 <= 1'h0;
    end else begin
      _T_72478_12_1_0 <= _T_39941_12_1_0;
    end
    if (_T_178) begin
      _T_72478_13_0_0 <= 1'h0;
    end else begin
      _T_72478_13_0_0 <= _T_39941_13_0_0;
    end
    if (_T_178) begin
      _T_72478_13_1_0 <= 1'h0;
    end else begin
      _T_72478_13_1_0 <= _T_39941_13_1_0;
    end
    if (_T_178) begin
      _T_72478_14_0_0 <= 1'h0;
    end else begin
      _T_72478_14_0_0 <= _T_39941_14_0_0;
    end
    if (_T_178) begin
      _T_72478_14_1_0 <= 1'h0;
    end else begin
      _T_72478_14_1_0 <= _T_39941_14_1_0;
    end
    if (_T_178) begin
      _T_72478_15_0_0 <= 1'h0;
    end else begin
      _T_72478_15_0_0 <= _T_39941_15_0_0;
    end
    if (_T_178) begin
      _T_72478_15_1_0 <= 1'h0;
    end else begin
      _T_72478_15_1_0 <= _T_39941_15_1_0;
    end
    _T_86710 <= _T_86705 != 32'h0;
    _T_86712 <= _T_86710;
    _T_86714 <= _T_86712;
    _T_86716 <= _T_86714;
    _T_87674_0_0 <= {_T_87211,_T_87216};
    _T_87674_1_0 <= {_T_87222,_T_87227};
    _T_87674_2_0 <= {_T_87233,_T_87238};
    _T_87674_3_0 <= {_T_87244,_T_87249};
    _T_87674_4_0 <= {_T_87255,_T_87260};
    _T_87674_5_0 <= {_T_87266,_T_87271};
    _T_87674_6_0 <= {_T_87277,_T_87282};
    _T_87674_7_0 <= {_T_87288,_T_87293};
    _T_87674_8_0 <= {_T_87299,_T_87304};
    _T_87674_9_0 <= {_T_87310,_T_87315};
    _T_87674_10_0 <= {_T_87321,_T_87326};
    _T_87674_11_0 <= {_T_87332,_T_87337};
    _T_87674_12_0 <= {_T_87343,_T_87348};
    _T_87674_13_0 <= {_T_87354,_T_87359};
    _T_87674_14_0 <= {_T_87365,_T_87370};
    _T_87674_15_0 <= {_T_87376,_T_87381};
    _T_88155_0_0 <= _T_88203 | _T_87674_3_0;
    _T_88155_1_0 <= _T_88206 | _T_87674_7_0;
    _T_88155_2_0 <= _T_88209 | _T_87674_11_0;
    _T_88155_3_0 <= _T_88212 | _T_87674_15_0;
    _T_88225_0_0 <= _T_88246 | _T_88155_3_0;
    _T_88249 <= _T_88225_0_0;
    _T_89522_0_0 <= io_sc2buf_wt_rd_addr_valid & _T_88531;
    _T_89522_0_1 <= io_sc2buf_wt_rd_addr_valid & _T_88531;
    _T_89522_1_0 <= io_sc2buf_wt_rd_addr_valid & _T_88539;
    _T_89522_1_1 <= io_sc2buf_wt_rd_addr_valid & _T_88539;
    _T_89522_2_0 <= io_sc2buf_wt_rd_addr_valid & _T_88547;
    _T_89522_2_1 <= io_sc2buf_wt_rd_addr_valid & _T_88547;
    _T_89522_3_0 <= io_sc2buf_wt_rd_addr_valid & _T_88555;
    _T_89522_3_1 <= io_sc2buf_wt_rd_addr_valid & _T_88555;
    _T_89522_4_0 <= io_sc2buf_wt_rd_addr_valid & _T_88563;
    _T_89522_4_1 <= io_sc2buf_wt_rd_addr_valid & _T_88563;
    _T_89522_5_0 <= io_sc2buf_wt_rd_addr_valid & _T_88571;
    _T_89522_5_1 <= io_sc2buf_wt_rd_addr_valid & _T_88571;
    _T_89522_6_0 <= io_sc2buf_wt_rd_addr_valid & _T_88579;
    _T_89522_6_1 <= io_sc2buf_wt_rd_addr_valid & _T_88579;
    _T_89522_7_0 <= io_sc2buf_wt_rd_addr_valid & _T_88587;
    _T_89522_7_1 <= io_sc2buf_wt_rd_addr_valid & _T_88587;
    _T_89522_8_0 <= io_sc2buf_wt_rd_addr_valid & _T_88595;
    _T_89522_8_1 <= io_sc2buf_wt_rd_addr_valid & _T_88595;
    _T_89522_9_0 <= io_sc2buf_wt_rd_addr_valid & _T_88603;
    _T_89522_9_1 <= io_sc2buf_wt_rd_addr_valid & _T_88603;
    _T_89522_10_0 <= io_sc2buf_wt_rd_addr_valid & _T_88611;
    _T_89522_10_1 <= io_sc2buf_wt_rd_addr_valid & _T_88611;
    _T_89522_11_0 <= io_sc2buf_wt_rd_addr_valid & _T_88619;
    _T_89522_11_1 <= io_sc2buf_wt_rd_addr_valid & _T_88619;
    _T_89522_12_0 <= io_sc2buf_wt_rd_addr_valid & _T_88627;
    _T_89522_12_1 <= io_sc2buf_wt_rd_addr_valid & _T_88627;
    _T_89522_13_0 <= io_sc2buf_wt_rd_addr_valid & _T_88635;
    _T_89522_13_1 <= io_sc2buf_wt_rd_addr_valid & _T_88635;
    _T_89522_14_0 <= io_sc2buf_wt_rd_addr_valid & _T_88643;
    _T_89522_14_1 <= io_sc2buf_wt_rd_addr_valid & _T_88643;
    _T_89522_15_0 <= io_sc2buf_wt_rd_addr_valid & _T_88651;
    _T_89522_15_1 <= io_sc2buf_wt_rd_addr_valid & _T_88651;
    _T_91073_0_0 <= _T_89522_0_0;
    _T_91073_0_1 <= _T_89522_0_1;
    _T_91073_1_0 <= _T_89522_1_0;
    _T_91073_1_1 <= _T_89522_1_1;
    _T_91073_2_0 <= _T_89522_2_0;
    _T_91073_2_1 <= _T_89522_2_1;
    _T_91073_3_0 <= _T_89522_3_0;
    _T_91073_3_1 <= _T_89522_3_1;
    _T_91073_4_0 <= _T_89522_4_0;
    _T_91073_4_1 <= _T_89522_4_1;
    _T_91073_5_0 <= _T_89522_5_0;
    _T_91073_5_1 <= _T_89522_5_1;
    _T_91073_6_0 <= _T_89522_6_0;
    _T_91073_6_1 <= _T_89522_6_1;
    _T_91073_7_0 <= _T_89522_7_0;
    _T_91073_7_1 <= _T_89522_7_1;
    _T_91073_8_0 <= _T_89522_8_0;
    _T_91073_8_1 <= _T_89522_8_1;
    _T_91073_9_0 <= _T_89522_9_0;
    _T_91073_9_1 <= _T_89522_9_1;
    _T_91073_10_0 <= _T_89522_10_0;
    _T_91073_10_1 <= _T_89522_10_1;
    _T_91073_11_0 <= _T_89522_11_0;
    _T_91073_11_1 <= _T_89522_11_1;
    _T_91073_12_0 <= _T_89522_12_0;
    _T_91073_12_1 <= _T_89522_12_1;
    _T_91073_13_0 <= _T_89522_13_0;
    _T_91073_13_1 <= _T_89522_13_1;
    _T_91073_14_0 <= _T_89522_14_0;
    _T_91073_14_1 <= _T_89522_14_1;
    _T_91073_15_0 <= _T_89522_15_0;
    _T_91073_15_1 <= _T_89522_15_1;
    _T_92368 <= _T_92363 != 32'h0;
    _T_92370 <= _T_92368;
    _T_92372 <= _T_92370;
    _T_92374 <= _T_92372;
    _T_92609_0 <= {_T_92401,_T_92406};
    _T_92609_1 <= {_T_92412,_T_92417};
    _T_92609_2 <= {_T_92423,_T_92428};
    _T_92609_3 <= {_T_92434,_T_92439};
    _T_92609_4 <= {_T_92445,_T_92450};
    _T_92609_5 <= {_T_92456,_T_92461};
    _T_92609_6 <= {_T_92467,_T_92472};
    _T_92609_7 <= {_T_92478,_T_92483};
    _T_92609_8 <= {_T_92489,_T_92494};
    _T_92609_9 <= {_T_92500,_T_92505};
    _T_92609_10 <= {_T_92511,_T_92516};
    _T_92609_11 <= {_T_92522,_T_92527};
    _T_92609_12 <= {_T_92533,_T_92538};
    _T_92609_13 <= {_T_92544,_T_92549};
    _T_92609_14 <= {_T_92555,_T_92560};
    _T_92609_15 <= {_T_92566,_T_92571};
    _T_92665_0 <= _T_92673 | _T_92609_3;
    _T_92665_1 <= _T_92676 | _T_92609_7;
    _T_92665_2 <= _T_92679 | _T_92609_11;
    _T_92665_3 <= _T_92682 | _T_92609_15;
    _T_92687_0 <= _T_92692 | _T_92665_3;
    _T_92695 <= _T_92687_0;
    if (_T_178) begin
      _T_94145_0_0 <= 1'h0;
    end else begin
      _T_94145_0_0 <= _T_95463;
    end
    if (_T_178) begin
      _T_94145_0_1 <= 1'h0;
    end else begin
      _T_94145_0_1 <= _T_95463;
    end
    if (_T_178) begin
      _T_94145_1_0 <= 1'h0;
    end else begin
      _T_94145_1_0 <= _T_95487;
    end
    if (_T_178) begin
      _T_94145_1_1 <= 1'h0;
    end else begin
      _T_94145_1_1 <= _T_95487;
    end
    if (_T_178) begin
      _T_94145_2_0 <= 1'h0;
    end else begin
      _T_94145_2_0 <= _T_95511;
    end
    if (_T_178) begin
      _T_94145_2_1 <= 1'h0;
    end else begin
      _T_94145_2_1 <= _T_95511;
    end
    if (_T_178) begin
      _T_94145_3_0 <= 1'h0;
    end else begin
      _T_94145_3_0 <= _T_95535;
    end
    if (_T_178) begin
      _T_94145_3_1 <= 1'h0;
    end else begin
      _T_94145_3_1 <= _T_95535;
    end
    if (_T_178) begin
      _T_94145_4_0 <= 1'h0;
    end else begin
      _T_94145_4_0 <= _T_95559;
    end
    if (_T_178) begin
      _T_94145_4_1 <= 1'h0;
    end else begin
      _T_94145_4_1 <= _T_95559;
    end
    if (_T_178) begin
      _T_94145_5_0 <= 1'h0;
    end else begin
      _T_94145_5_0 <= _T_95583;
    end
    if (_T_178) begin
      _T_94145_5_1 <= 1'h0;
    end else begin
      _T_94145_5_1 <= _T_95583;
    end
    if (_T_178) begin
      _T_94145_6_0 <= 1'h0;
    end else begin
      _T_94145_6_0 <= _T_95607;
    end
    if (_T_178) begin
      _T_94145_6_1 <= 1'h0;
    end else begin
      _T_94145_6_1 <= _T_95607;
    end
    if (_T_178) begin
      _T_94145_7_0 <= 1'h0;
    end else begin
      _T_94145_7_0 <= _T_95631;
    end
    if (_T_178) begin
      _T_94145_7_1 <= 1'h0;
    end else begin
      _T_94145_7_1 <= _T_95631;
    end
    if (_T_178) begin
      _T_94145_8_0 <= 1'h0;
    end else begin
      _T_94145_8_0 <= _T_95655;
    end
    if (_T_178) begin
      _T_94145_8_1 <= 1'h0;
    end else begin
      _T_94145_8_1 <= _T_95655;
    end
    if (_T_178) begin
      _T_94145_9_0 <= 1'h0;
    end else begin
      _T_94145_9_0 <= _T_95679;
    end
    if (_T_178) begin
      _T_94145_9_1 <= 1'h0;
    end else begin
      _T_94145_9_1 <= _T_95679;
    end
    if (_T_178) begin
      _T_94145_10_0 <= 1'h0;
    end else begin
      _T_94145_10_0 <= _T_95703;
    end
    if (_T_178) begin
      _T_94145_10_1 <= 1'h0;
    end else begin
      _T_94145_10_1 <= _T_95703;
    end
    if (_T_178) begin
      _T_94145_11_0 <= 1'h0;
    end else begin
      _T_94145_11_0 <= _T_95727;
    end
    if (_T_178) begin
      _T_94145_11_1 <= 1'h0;
    end else begin
      _T_94145_11_1 <= _T_95727;
    end
    if (_T_178) begin
      _T_94145_12_0 <= 1'h0;
    end else begin
      _T_94145_12_0 <= _T_95751;
    end
    if (_T_178) begin
      _T_94145_12_1 <= 1'h0;
    end else begin
      _T_94145_12_1 <= _T_95751;
    end
    if (_T_178) begin
      _T_94145_13_0 <= 1'h0;
    end else begin
      _T_94145_13_0 <= _T_95775;
    end
    if (_T_178) begin
      _T_94145_13_1 <= 1'h0;
    end else begin
      _T_94145_13_1 <= _T_95775;
    end
    if (_T_178) begin
      _T_94145_14_0 <= 1'h0;
    end else begin
      _T_94145_14_0 <= _T_95799;
    end
    if (_T_178) begin
      _T_94145_14_1 <= 1'h0;
    end else begin
      _T_94145_14_1 <= _T_95799;
    end
    if (_T_178) begin
      _T_94145_15_0 <= 1'h0;
    end else begin
      _T_94145_15_0 <= _T_95823;
    end
    if (_T_178) begin
      _T_94145_15_1 <= 1'h0;
    end else begin
      _T_94145_15_1 <= _T_95823;
    end
    _T_95257_0_0 <= _T_95468 | _T_95473;
    _T_95257_0_1 <= _T_95468 | _T_95473;
    _T_95257_1_0 <= _T_95492 | _T_95497;
    _T_95257_1_1 <= _T_95492 | _T_95497;
    _T_95257_2_0 <= _T_95516 | _T_95521;
    _T_95257_2_1 <= _T_95516 | _T_95521;
    _T_95257_3_0 <= _T_95540 | _T_95545;
    _T_95257_3_1 <= _T_95540 | _T_95545;
    _T_95257_4_0 <= _T_95564 | _T_95569;
    _T_95257_4_1 <= _T_95564 | _T_95569;
    _T_95257_5_0 <= _T_95588 | _T_95593;
    _T_95257_5_1 <= _T_95588 | _T_95593;
    _T_95257_6_0 <= _T_95612 | _T_95617;
    _T_95257_6_1 <= _T_95612 | _T_95617;
    _T_95257_7_0 <= _T_95636 | _T_95641;
    _T_95257_7_1 <= _T_95636 | _T_95641;
    _T_95257_8_0 <= _T_95660 | _T_95665;
    _T_95257_8_1 <= _T_95660 | _T_95665;
    _T_95257_9_0 <= _T_95684 | _T_95689;
    _T_95257_9_1 <= _T_95684 | _T_95689;
    _T_95257_10_0 <= _T_95708 | _T_95713;
    _T_95257_10_1 <= _T_95708 | _T_95713;
    _T_95257_11_0 <= _T_95732 | _T_95737;
    _T_95257_11_1 <= _T_95732 | _T_95737;
    _T_95257_12_0 <= _T_95756 | _T_95761;
    _T_95257_12_1 <= _T_95756 | _T_95761;
    _T_95257_13_0 <= _T_95780 | _T_95785;
    _T_95257_13_1 <= _T_95780 | _T_95785;
    _T_95257_14_0 <= _T_95804 | _T_95809;
    _T_95257_14_1 <= _T_95804 | _T_95809;
    _T_95257_15_0 <= _T_95828 | _T_95833;
    _T_95257_15_1 <= _T_95828 | _T_95833;
  end
endmodule
