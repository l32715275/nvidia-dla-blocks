module NV_NVDLA_CMAC_CORE_rt_in_dft( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input        io_nvdla_core_clk, // @[:@6.4]
  input        io_nvdla_core_rstn, // @[:@6.4]
  input        io_sc2mac_dat_valid, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_0, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_1, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_2, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_3, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_4, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_5, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_6, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_7, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_8, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_9, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_10, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_11, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_12, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_13, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_14, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_15, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_16, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_17, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_18, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_19, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_20, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_21, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_22, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_23, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_24, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_25, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_26, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_27, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_28, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_29, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_30, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_31, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_32, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_33, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_34, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_35, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_36, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_37, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_38, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_39, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_40, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_41, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_42, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_43, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_44, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_45, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_46, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_47, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_48, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_49, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_50, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_51, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_52, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_53, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_54, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_55, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_56, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_57, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_58, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_59, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_60, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_61, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_62, // @[:@6.4]
  input        io_sc2mac_dat_bits_mask_63, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_0, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_1, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_2, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_3, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_4, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_5, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_6, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_7, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_8, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_9, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_10, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_11, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_12, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_13, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_14, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_15, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_16, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_17, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_18, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_19, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_20, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_21, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_22, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_23, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_24, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_25, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_26, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_27, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_28, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_29, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_30, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_31, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_32, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_33, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_34, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_35, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_36, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_37, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_38, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_39, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_40, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_41, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_42, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_43, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_44, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_45, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_46, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_47, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_48, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_49, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_50, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_51, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_52, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_53, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_54, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_55, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_56, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_57, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_58, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_59, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_60, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_61, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_62, // @[:@6.4]
  input  [7:0] io_sc2mac_dat_bits_data_63, // @[:@6.4]
  input  [8:0] io_sc2mac_dat_bits_pd, // @[:@6.4]
  input        io_sc2mac_wt_valid, // @[:@6.4]
  input        io_sc2mac_wt_bits_sel_0, // @[:@6.4]
  input        io_sc2mac_wt_bits_sel_1, // @[:@6.4]
  input        io_sc2mac_wt_bits_sel_2, // @[:@6.4]
  input        io_sc2mac_wt_bits_sel_3, // @[:@6.4]
  input        io_sc2mac_wt_bits_sel_4, // @[:@6.4]
  input        io_sc2mac_wt_bits_sel_5, // @[:@6.4]
  input        io_sc2mac_wt_bits_sel_6, // @[:@6.4]
  input        io_sc2mac_wt_bits_sel_7, // @[:@6.4]
  input        io_sc2mac_wt_bits_sel_8, // @[:@6.4]
  input        io_sc2mac_wt_bits_sel_9, // @[:@6.4]
  input        io_sc2mac_wt_bits_sel_10, // @[:@6.4]
  input        io_sc2mac_wt_bits_sel_11, // @[:@6.4]
  input        io_sc2mac_wt_bits_sel_12, // @[:@6.4]
  input        io_sc2mac_wt_bits_sel_13, // @[:@6.4]
  input        io_sc2mac_wt_bits_sel_14, // @[:@6.4]
  input        io_sc2mac_wt_bits_sel_15, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_0, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_1, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_2, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_3, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_4, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_5, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_6, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_7, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_8, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_9, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_10, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_11, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_12, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_13, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_14, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_15, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_16, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_17, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_18, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_19, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_20, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_21, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_22, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_23, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_24, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_25, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_26, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_27, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_28, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_29, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_30, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_31, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_32, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_33, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_34, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_35, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_36, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_37, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_38, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_39, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_40, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_41, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_42, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_43, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_44, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_45, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_46, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_47, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_48, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_49, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_50, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_51, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_52, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_53, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_54, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_55, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_56, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_57, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_58, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_59, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_60, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_61, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_62, // @[:@6.4]
  input        io_sc2mac_wt_bits_mask_63, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_0, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_1, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_2, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_3, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_4, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_5, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_6, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_7, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_8, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_9, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_10, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_11, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_12, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_13, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_14, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_15, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_16, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_17, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_18, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_19, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_20, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_21, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_22, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_23, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_24, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_25, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_26, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_27, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_28, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_29, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_30, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_31, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_32, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_33, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_34, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_35, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_36, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_37, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_38, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_39, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_40, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_41, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_42, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_43, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_44, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_45, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_46, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_47, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_48, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_49, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_50, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_51, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_52, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_53, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_54, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_55, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_56, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_57, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_58, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_59, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_60, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_61, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_62, // @[:@6.4]
  input  [7:0] io_sc2mac_wt_bits_data_63, // @[:@6.4]
  output       io_in_dat_valid, // @[:@6.4]
  output       io_in_dat_bits_mask_0, // @[:@6.4]
  output       io_in_dat_bits_mask_1, // @[:@6.4]
  output       io_in_dat_bits_mask_2, // @[:@6.4]
  output       io_in_dat_bits_mask_3, // @[:@6.4]
  output       io_in_dat_bits_mask_4, // @[:@6.4]
  output       io_in_dat_bits_mask_5, // @[:@6.4]
  output       io_in_dat_bits_mask_6, // @[:@6.4]
  output       io_in_dat_bits_mask_7, // @[:@6.4]
  output       io_in_dat_bits_mask_8, // @[:@6.4]
  output       io_in_dat_bits_mask_9, // @[:@6.4]
  output       io_in_dat_bits_mask_10, // @[:@6.4]
  output       io_in_dat_bits_mask_11, // @[:@6.4]
  output       io_in_dat_bits_mask_12, // @[:@6.4]
  output       io_in_dat_bits_mask_13, // @[:@6.4]
  output       io_in_dat_bits_mask_14, // @[:@6.4]
  output       io_in_dat_bits_mask_15, // @[:@6.4]
  output       io_in_dat_bits_mask_16, // @[:@6.4]
  output       io_in_dat_bits_mask_17, // @[:@6.4]
  output       io_in_dat_bits_mask_18, // @[:@6.4]
  output       io_in_dat_bits_mask_19, // @[:@6.4]
  output       io_in_dat_bits_mask_20, // @[:@6.4]
  output       io_in_dat_bits_mask_21, // @[:@6.4]
  output       io_in_dat_bits_mask_22, // @[:@6.4]
  output       io_in_dat_bits_mask_23, // @[:@6.4]
  output       io_in_dat_bits_mask_24, // @[:@6.4]
  output       io_in_dat_bits_mask_25, // @[:@6.4]
  output       io_in_dat_bits_mask_26, // @[:@6.4]
  output       io_in_dat_bits_mask_27, // @[:@6.4]
  output       io_in_dat_bits_mask_28, // @[:@6.4]
  output       io_in_dat_bits_mask_29, // @[:@6.4]
  output       io_in_dat_bits_mask_30, // @[:@6.4]
  output       io_in_dat_bits_mask_31, // @[:@6.4]
  output       io_in_dat_bits_mask_32, // @[:@6.4]
  output       io_in_dat_bits_mask_33, // @[:@6.4]
  output       io_in_dat_bits_mask_34, // @[:@6.4]
  output       io_in_dat_bits_mask_35, // @[:@6.4]
  output       io_in_dat_bits_mask_36, // @[:@6.4]
  output       io_in_dat_bits_mask_37, // @[:@6.4]
  output       io_in_dat_bits_mask_38, // @[:@6.4]
  output       io_in_dat_bits_mask_39, // @[:@6.4]
  output       io_in_dat_bits_mask_40, // @[:@6.4]
  output       io_in_dat_bits_mask_41, // @[:@6.4]
  output       io_in_dat_bits_mask_42, // @[:@6.4]
  output       io_in_dat_bits_mask_43, // @[:@6.4]
  output       io_in_dat_bits_mask_44, // @[:@6.4]
  output       io_in_dat_bits_mask_45, // @[:@6.4]
  output       io_in_dat_bits_mask_46, // @[:@6.4]
  output       io_in_dat_bits_mask_47, // @[:@6.4]
  output       io_in_dat_bits_mask_48, // @[:@6.4]
  output       io_in_dat_bits_mask_49, // @[:@6.4]
  output       io_in_dat_bits_mask_50, // @[:@6.4]
  output       io_in_dat_bits_mask_51, // @[:@6.4]
  output       io_in_dat_bits_mask_52, // @[:@6.4]
  output       io_in_dat_bits_mask_53, // @[:@6.4]
  output       io_in_dat_bits_mask_54, // @[:@6.4]
  output       io_in_dat_bits_mask_55, // @[:@6.4]
  output       io_in_dat_bits_mask_56, // @[:@6.4]
  output       io_in_dat_bits_mask_57, // @[:@6.4]
  output       io_in_dat_bits_mask_58, // @[:@6.4]
  output       io_in_dat_bits_mask_59, // @[:@6.4]
  output       io_in_dat_bits_mask_60, // @[:@6.4]
  output       io_in_dat_bits_mask_61, // @[:@6.4]
  output       io_in_dat_bits_mask_62, // @[:@6.4]
  output       io_in_dat_bits_mask_63, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_0, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_1, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_2, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_3, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_4, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_5, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_6, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_7, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_8, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_9, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_10, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_11, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_12, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_13, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_14, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_15, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_16, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_17, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_18, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_19, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_20, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_21, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_22, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_23, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_24, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_25, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_26, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_27, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_28, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_29, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_30, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_31, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_32, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_33, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_34, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_35, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_36, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_37, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_38, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_39, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_40, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_41, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_42, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_43, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_44, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_45, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_46, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_47, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_48, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_49, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_50, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_51, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_52, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_53, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_54, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_55, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_56, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_57, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_58, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_59, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_60, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_61, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_62, // @[:@6.4]
  output [7:0] io_in_dat_bits_data_63, // @[:@6.4]
  output [8:0] io_in_dat_bits_pd, // @[:@6.4]
  output       io_in_wt_valid, // @[:@6.4]
  output       io_in_wt_bits_sel_0, // @[:@6.4]
  output       io_in_wt_bits_sel_1, // @[:@6.4]
  output       io_in_wt_bits_sel_2, // @[:@6.4]
  output       io_in_wt_bits_sel_3, // @[:@6.4]
  output       io_in_wt_bits_sel_4, // @[:@6.4]
  output       io_in_wt_bits_sel_5, // @[:@6.4]
  output       io_in_wt_bits_sel_6, // @[:@6.4]
  output       io_in_wt_bits_sel_7, // @[:@6.4]
  output       io_in_wt_bits_sel_8, // @[:@6.4]
  output       io_in_wt_bits_sel_9, // @[:@6.4]
  output       io_in_wt_bits_sel_10, // @[:@6.4]
  output       io_in_wt_bits_sel_11, // @[:@6.4]
  output       io_in_wt_bits_sel_12, // @[:@6.4]
  output       io_in_wt_bits_sel_13, // @[:@6.4]
  output       io_in_wt_bits_sel_14, // @[:@6.4]
  output       io_in_wt_bits_sel_15, // @[:@6.4]
  output       io_in_wt_bits_mask_0, // @[:@6.4]
  output       io_in_wt_bits_mask_1, // @[:@6.4]
  output       io_in_wt_bits_mask_2, // @[:@6.4]
  output       io_in_wt_bits_mask_3, // @[:@6.4]
  output       io_in_wt_bits_mask_4, // @[:@6.4]
  output       io_in_wt_bits_mask_5, // @[:@6.4]
  output       io_in_wt_bits_mask_6, // @[:@6.4]
  output       io_in_wt_bits_mask_7, // @[:@6.4]
  output       io_in_wt_bits_mask_8, // @[:@6.4]
  output       io_in_wt_bits_mask_9, // @[:@6.4]
  output       io_in_wt_bits_mask_10, // @[:@6.4]
  output       io_in_wt_bits_mask_11, // @[:@6.4]
  output       io_in_wt_bits_mask_12, // @[:@6.4]
  output       io_in_wt_bits_mask_13, // @[:@6.4]
  output       io_in_wt_bits_mask_14, // @[:@6.4]
  output       io_in_wt_bits_mask_15, // @[:@6.4]
  output       io_in_wt_bits_mask_16, // @[:@6.4]
  output       io_in_wt_bits_mask_17, // @[:@6.4]
  output       io_in_wt_bits_mask_18, // @[:@6.4]
  output       io_in_wt_bits_mask_19, // @[:@6.4]
  output       io_in_wt_bits_mask_20, // @[:@6.4]
  output       io_in_wt_bits_mask_21, // @[:@6.4]
  output       io_in_wt_bits_mask_22, // @[:@6.4]
  output       io_in_wt_bits_mask_23, // @[:@6.4]
  output       io_in_wt_bits_mask_24, // @[:@6.4]
  output       io_in_wt_bits_mask_25, // @[:@6.4]
  output       io_in_wt_bits_mask_26, // @[:@6.4]
  output       io_in_wt_bits_mask_27, // @[:@6.4]
  output       io_in_wt_bits_mask_28, // @[:@6.4]
  output       io_in_wt_bits_mask_29, // @[:@6.4]
  output       io_in_wt_bits_mask_30, // @[:@6.4]
  output       io_in_wt_bits_mask_31, // @[:@6.4]
  output       io_in_wt_bits_mask_32, // @[:@6.4]
  output       io_in_wt_bits_mask_33, // @[:@6.4]
  output       io_in_wt_bits_mask_34, // @[:@6.4]
  output       io_in_wt_bits_mask_35, // @[:@6.4]
  output       io_in_wt_bits_mask_36, // @[:@6.4]
  output       io_in_wt_bits_mask_37, // @[:@6.4]
  output       io_in_wt_bits_mask_38, // @[:@6.4]
  output       io_in_wt_bits_mask_39, // @[:@6.4]
  output       io_in_wt_bits_mask_40, // @[:@6.4]
  output       io_in_wt_bits_mask_41, // @[:@6.4]
  output       io_in_wt_bits_mask_42, // @[:@6.4]
  output       io_in_wt_bits_mask_43, // @[:@6.4]
  output       io_in_wt_bits_mask_44, // @[:@6.4]
  output       io_in_wt_bits_mask_45, // @[:@6.4]
  output       io_in_wt_bits_mask_46, // @[:@6.4]
  output       io_in_wt_bits_mask_47, // @[:@6.4]
  output       io_in_wt_bits_mask_48, // @[:@6.4]
  output       io_in_wt_bits_mask_49, // @[:@6.4]
  output       io_in_wt_bits_mask_50, // @[:@6.4]
  output       io_in_wt_bits_mask_51, // @[:@6.4]
  output       io_in_wt_bits_mask_52, // @[:@6.4]
  output       io_in_wt_bits_mask_53, // @[:@6.4]
  output       io_in_wt_bits_mask_54, // @[:@6.4]
  output       io_in_wt_bits_mask_55, // @[:@6.4]
  output       io_in_wt_bits_mask_56, // @[:@6.4]
  output       io_in_wt_bits_mask_57, // @[:@6.4]
  output       io_in_wt_bits_mask_58, // @[:@6.4]
  output       io_in_wt_bits_mask_59, // @[:@6.4]
  output       io_in_wt_bits_mask_60, // @[:@6.4]
  output       io_in_wt_bits_mask_61, // @[:@6.4]
  output       io_in_wt_bits_mask_62, // @[:@6.4]
  output       io_in_wt_bits_mask_63, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_0, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_1, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_2, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_3, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_4, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_5, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_6, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_7, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_8, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_9, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_10, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_11, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_12, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_13, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_14, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_15, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_16, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_17, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_18, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_19, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_20, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_21, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_22, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_23, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_24, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_25, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_26, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_27, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_28, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_29, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_30, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_31, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_32, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_33, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_34, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_35, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_36, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_37, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_38, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_39, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_40, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_41, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_42, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_43, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_44, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_45, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_46, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_47, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_48, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_49, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_50, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_51, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_52, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_53, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_54, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_55, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_56, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_57, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_58, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_59, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_60, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_61, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_62, // @[:@6.4]
  output [7:0] io_in_wt_bits_data_63 // @[:@6.4]
);
  wire  _T_3014; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 45:38:@8.4]
  reg [7:0] _T_3085_0; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_0;
  reg [7:0] _T_3085_1; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_1;
  reg [7:0] _T_3085_2; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_2;
  reg [7:0] _T_3085_3; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_3;
  reg [7:0] _T_3085_4; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_4;
  reg [7:0] _T_3085_5; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_5;
  reg [7:0] _T_3085_6; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_6;
  reg [7:0] _T_3085_7; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_7;
  reg [7:0] _T_3085_8; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_8;
  reg [7:0] _T_3085_9; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_9;
  reg [7:0] _T_3085_10; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_10;
  reg [7:0] _T_3085_11; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_11;
  reg [7:0] _T_3085_12; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_12;
  reg [7:0] _T_3085_13; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_13;
  reg [7:0] _T_3085_14; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_14;
  reg [7:0] _T_3085_15; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_15;
  reg [7:0] _T_3085_16; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_16;
  reg [7:0] _T_3085_17; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_17;
  reg [7:0] _T_3085_18; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_18;
  reg [7:0] _T_3085_19; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_19;
  reg [7:0] _T_3085_20; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_20;
  reg [7:0] _T_3085_21; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_21;
  reg [7:0] _T_3085_22; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_22;
  reg [7:0] _T_3085_23; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_23;
  reg [7:0] _T_3085_24; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_24;
  reg [7:0] _T_3085_25; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_25;
  reg [7:0] _T_3085_26; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_26;
  reg [7:0] _T_3085_27; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_27;
  reg [7:0] _T_3085_28; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_28;
  reg [7:0] _T_3085_29; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_29;
  reg [7:0] _T_3085_30; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_30;
  reg [7:0] _T_3085_31; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_31;
  reg [7:0] _T_3085_32; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_32;
  reg [7:0] _T_3085_33; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_33;
  reg [7:0] _T_3085_34; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_34;
  reg [7:0] _T_3085_35; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_35;
  reg [7:0] _T_3085_36; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_36;
  reg [7:0] _T_3085_37; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_37;
  reg [7:0] _T_3085_38; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_38;
  reg [7:0] _T_3085_39; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_39;
  reg [7:0] _T_3085_40; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_40;
  reg [7:0] _T_3085_41; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_41;
  reg [7:0] _T_3085_42; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_42;
  reg [7:0] _T_3085_43; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_43;
  reg [7:0] _T_3085_44; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_44;
  reg [7:0] _T_3085_45; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_45;
  reg [7:0] _T_3085_46; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_46;
  reg [7:0] _T_3085_47; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_47;
  reg [7:0] _T_3085_48; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_48;
  reg [7:0] _T_3085_49; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_49;
  reg [7:0] _T_3085_50; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_50;
  reg [7:0] _T_3085_51; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_51;
  reg [7:0] _T_3085_52; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_52;
  reg [7:0] _T_3085_53; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_53;
  reg [7:0] _T_3085_54; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_54;
  reg [7:0] _T_3085_55; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_55;
  reg [7:0] _T_3085_56; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_56;
  reg [7:0] _T_3085_57; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_57;
  reg [7:0] _T_3085_58; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_58;
  reg [7:0] _T_3085_59; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_59;
  reg [7:0] _T_3085_60; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_60;
  reg [7:0] _T_3085_61; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_61;
  reg [7:0] _T_3085_62; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_62;
  reg [7:0] _T_3085_63; // @[retiming.scala 9:92:@10.4]
  reg [31:0] _RAND_63;
  reg [7:0] _T_3152_0; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_64;
  reg [7:0] _T_3152_1; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_65;
  reg [7:0] _T_3152_2; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_66;
  reg [7:0] _T_3152_3; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_67;
  reg [7:0] _T_3152_4; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_68;
  reg [7:0] _T_3152_5; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_69;
  reg [7:0] _T_3152_6; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_70;
  reg [7:0] _T_3152_7; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_71;
  reg [7:0] _T_3152_8; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_72;
  reg [7:0] _T_3152_9; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_73;
  reg [7:0] _T_3152_10; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_74;
  reg [7:0] _T_3152_11; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_75;
  reg [7:0] _T_3152_12; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_76;
  reg [7:0] _T_3152_13; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_77;
  reg [7:0] _T_3152_14; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_78;
  reg [7:0] _T_3152_15; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_79;
  reg [7:0] _T_3152_16; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_80;
  reg [7:0] _T_3152_17; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_81;
  reg [7:0] _T_3152_18; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_82;
  reg [7:0] _T_3152_19; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_83;
  reg [7:0] _T_3152_20; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_84;
  reg [7:0] _T_3152_21; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_85;
  reg [7:0] _T_3152_22; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_86;
  reg [7:0] _T_3152_23; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_87;
  reg [7:0] _T_3152_24; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_88;
  reg [7:0] _T_3152_25; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_89;
  reg [7:0] _T_3152_26; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_90;
  reg [7:0] _T_3152_27; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_91;
  reg [7:0] _T_3152_28; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_92;
  reg [7:0] _T_3152_29; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_93;
  reg [7:0] _T_3152_30; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_94;
  reg [7:0] _T_3152_31; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_95;
  reg [7:0] _T_3152_32; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_96;
  reg [7:0] _T_3152_33; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_97;
  reg [7:0] _T_3152_34; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_98;
  reg [7:0] _T_3152_35; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_99;
  reg [7:0] _T_3152_36; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_100;
  reg [7:0] _T_3152_37; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_101;
  reg [7:0] _T_3152_38; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_102;
  reg [7:0] _T_3152_39; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_103;
  reg [7:0] _T_3152_40; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_104;
  reg [7:0] _T_3152_41; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_105;
  reg [7:0] _T_3152_42; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_106;
  reg [7:0] _T_3152_43; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_107;
  reg [7:0] _T_3152_44; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_108;
  reg [7:0] _T_3152_45; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_109;
  reg [7:0] _T_3152_46; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_110;
  reg [7:0] _T_3152_47; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_111;
  reg [7:0] _T_3152_48; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_112;
  reg [7:0] _T_3152_49; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_113;
  reg [7:0] _T_3152_50; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_114;
  reg [7:0] _T_3152_51; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_115;
  reg [7:0] _T_3152_52; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_116;
  reg [7:0] _T_3152_53; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_117;
  reg [7:0] _T_3152_54; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_118;
  reg [7:0] _T_3152_55; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_119;
  reg [7:0] _T_3152_56; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_120;
  reg [7:0] _T_3152_57; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_121;
  reg [7:0] _T_3152_58; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_122;
  reg [7:0] _T_3152_59; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_123;
  reg [7:0] _T_3152_60; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_124;
  reg [7:0] _T_3152_61; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_125;
  reg [7:0] _T_3152_62; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_126;
  reg [7:0] _T_3152_63; // @[retiming.scala 9:92:@11.4]
  reg [31:0] _RAND_127;
  reg  _T_3555_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_128;
  reg  _T_3555_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_129;
  reg  _T_3555_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_130;
  reg  _T_3555_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_131;
  reg  _T_3555_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_132;
  reg  _T_3555_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_133;
  reg  _T_3555_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_134;
  reg  _T_3555_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_135;
  reg  _T_3555_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_136;
  reg  _T_3555_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_137;
  reg  _T_3555_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_138;
  reg  _T_3555_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_139;
  reg  _T_3555_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_140;
  reg  _T_3555_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_141;
  reg  _T_3555_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_142;
  reg  _T_3555_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_143;
  reg  _T_3555_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_144;
  reg  _T_3555_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_145;
  reg  _T_3555_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_146;
  reg  _T_3555_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_147;
  reg  _T_3555_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_148;
  reg  _T_3555_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_149;
  reg  _T_3555_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_150;
  reg  _T_3555_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_151;
  reg  _T_3555_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_152;
  reg  _T_3555_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_153;
  reg  _T_3555_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_154;
  reg  _T_3555_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_155;
  reg  _T_3555_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_156;
  reg  _T_3555_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_157;
  reg  _T_3555_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_158;
  reg  _T_3555_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_159;
  reg  _T_3555_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_160;
  reg  _T_3555_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_161;
  reg  _T_3555_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_162;
  reg  _T_3555_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_163;
  reg  _T_3555_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_164;
  reg  _T_3555_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_165;
  reg  _T_3555_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_166;
  reg  _T_3555_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_167;
  reg  _T_3555_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_168;
  reg  _T_3555_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_169;
  reg  _T_3555_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_170;
  reg  _T_3555_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_171;
  reg  _T_3555_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_172;
  reg  _T_3555_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_173;
  reg  _T_3555_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_174;
  reg  _T_3555_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_175;
  reg  _T_3555_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_176;
  reg  _T_3555_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_177;
  reg  _T_3555_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_178;
  reg  _T_3555_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_179;
  reg  _T_3555_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_180;
  reg  _T_3555_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_181;
  reg  _T_3555_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_182;
  reg  _T_3555_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_183;
  reg  _T_3555_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_184;
  reg  _T_3555_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_185;
  reg  _T_3555_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_186;
  reg  _T_3555_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_187;
  reg  _T_3555_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_188;
  reg  _T_3555_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_189;
  reg  _T_3555_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_190;
  reg  _T_3555_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@78.4]
  reg [31:0] _RAND_191;
  reg  _T_4018_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_192;
  reg  _T_4018_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_193;
  reg  _T_4018_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_194;
  reg  _T_4018_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_195;
  reg  _T_4018_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_196;
  reg  _T_4018_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_197;
  reg  _T_4018_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_198;
  reg  _T_4018_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_199;
  reg  _T_4018_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_200;
  reg  _T_4018_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_201;
  reg  _T_4018_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_202;
  reg  _T_4018_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_203;
  reg  _T_4018_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_204;
  reg  _T_4018_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_205;
  reg  _T_4018_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_206;
  reg  _T_4018_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_207;
  reg  _T_4018_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_208;
  reg  _T_4018_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_209;
  reg  _T_4018_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_210;
  reg  _T_4018_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_211;
  reg  _T_4018_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_212;
  reg  _T_4018_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_213;
  reg  _T_4018_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_214;
  reg  _T_4018_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_215;
  reg  _T_4018_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_216;
  reg  _T_4018_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_217;
  reg  _T_4018_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_218;
  reg  _T_4018_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_219;
  reg  _T_4018_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_220;
  reg  _T_4018_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_221;
  reg  _T_4018_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_222;
  reg  _T_4018_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_223;
  reg  _T_4018_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_224;
  reg  _T_4018_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_225;
  reg  _T_4018_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_226;
  reg  _T_4018_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_227;
  reg  _T_4018_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_228;
  reg  _T_4018_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_229;
  reg  _T_4018_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_230;
  reg  _T_4018_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_231;
  reg  _T_4018_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_232;
  reg  _T_4018_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_233;
  reg  _T_4018_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_234;
  reg  _T_4018_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_235;
  reg  _T_4018_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_236;
  reg  _T_4018_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_237;
  reg  _T_4018_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_238;
  reg  _T_4018_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_239;
  reg  _T_4018_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_240;
  reg  _T_4018_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_241;
  reg  _T_4018_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_242;
  reg  _T_4018_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_243;
  reg  _T_4018_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_244;
  reg  _T_4018_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_245;
  reg  _T_4018_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_246;
  reg  _T_4018_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_247;
  reg  _T_4018_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_248;
  reg  _T_4018_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_249;
  reg  _T_4018_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_250;
  reg  _T_4018_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_251;
  reg  _T_4018_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_252;
  reg  _T_4018_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_253;
  reg  _T_4018_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_254;
  reg  _T_4018_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 50:70:@144.4]
  reg [31:0] _RAND_255;
  reg  _T_4219; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 52:70:@146.4]
  reg [31:0] _RAND_256;
  reg  _T_4222; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 52:70:@147.4]
  reg [31:0] _RAND_257;
  reg [8:0] _T_4227; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 54:70:@149.4]
  reg [31:0] _RAND_258;
  reg [8:0] _T_4230; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 54:70:@150.4]
  reg [31:0] _RAND_259;
  reg [7:0] _T_4301_0; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_260;
  reg [7:0] _T_4301_1; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_261;
  reg [7:0] _T_4301_2; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_262;
  reg [7:0] _T_4301_3; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_263;
  reg [7:0] _T_4301_4; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_264;
  reg [7:0] _T_4301_5; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_265;
  reg [7:0] _T_4301_6; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_266;
  reg [7:0] _T_4301_7; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_267;
  reg [7:0] _T_4301_8; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_268;
  reg [7:0] _T_4301_9; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_269;
  reg [7:0] _T_4301_10; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_270;
  reg [7:0] _T_4301_11; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_271;
  reg [7:0] _T_4301_12; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_272;
  reg [7:0] _T_4301_13; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_273;
  reg [7:0] _T_4301_14; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_274;
  reg [7:0] _T_4301_15; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_275;
  reg [7:0] _T_4301_16; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_276;
  reg [7:0] _T_4301_17; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_277;
  reg [7:0] _T_4301_18; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_278;
  reg [7:0] _T_4301_19; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_279;
  reg [7:0] _T_4301_20; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_280;
  reg [7:0] _T_4301_21; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_281;
  reg [7:0] _T_4301_22; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_282;
  reg [7:0] _T_4301_23; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_283;
  reg [7:0] _T_4301_24; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_284;
  reg [7:0] _T_4301_25; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_285;
  reg [7:0] _T_4301_26; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_286;
  reg [7:0] _T_4301_27; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_287;
  reg [7:0] _T_4301_28; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_288;
  reg [7:0] _T_4301_29; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_289;
  reg [7:0] _T_4301_30; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_290;
  reg [7:0] _T_4301_31; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_291;
  reg [7:0] _T_4301_32; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_292;
  reg [7:0] _T_4301_33; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_293;
  reg [7:0] _T_4301_34; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_294;
  reg [7:0] _T_4301_35; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_295;
  reg [7:0] _T_4301_36; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_296;
  reg [7:0] _T_4301_37; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_297;
  reg [7:0] _T_4301_38; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_298;
  reg [7:0] _T_4301_39; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_299;
  reg [7:0] _T_4301_40; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_300;
  reg [7:0] _T_4301_41; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_301;
  reg [7:0] _T_4301_42; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_302;
  reg [7:0] _T_4301_43; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_303;
  reg [7:0] _T_4301_44; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_304;
  reg [7:0] _T_4301_45; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_305;
  reg [7:0] _T_4301_46; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_306;
  reg [7:0] _T_4301_47; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_307;
  reg [7:0] _T_4301_48; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_308;
  reg [7:0] _T_4301_49; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_309;
  reg [7:0] _T_4301_50; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_310;
  reg [7:0] _T_4301_51; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_311;
  reg [7:0] _T_4301_52; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_312;
  reg [7:0] _T_4301_53; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_313;
  reg [7:0] _T_4301_54; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_314;
  reg [7:0] _T_4301_55; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_315;
  reg [7:0] _T_4301_56; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_316;
  reg [7:0] _T_4301_57; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_317;
  reg [7:0] _T_4301_58; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_318;
  reg [7:0] _T_4301_59; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_319;
  reg [7:0] _T_4301_60; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_320;
  reg [7:0] _T_4301_61; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_321;
  reg [7:0] _T_4301_62; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_322;
  reg [7:0] _T_4301_63; // @[retiming.scala 9:92:@152.4]
  reg [31:0] _RAND_323;
  reg [7:0] _T_4368_0; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_324;
  reg [7:0] _T_4368_1; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_325;
  reg [7:0] _T_4368_2; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_326;
  reg [7:0] _T_4368_3; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_327;
  reg [7:0] _T_4368_4; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_328;
  reg [7:0] _T_4368_5; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_329;
  reg [7:0] _T_4368_6; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_330;
  reg [7:0] _T_4368_7; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_331;
  reg [7:0] _T_4368_8; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_332;
  reg [7:0] _T_4368_9; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_333;
  reg [7:0] _T_4368_10; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_334;
  reg [7:0] _T_4368_11; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_335;
  reg [7:0] _T_4368_12; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_336;
  reg [7:0] _T_4368_13; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_337;
  reg [7:0] _T_4368_14; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_338;
  reg [7:0] _T_4368_15; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_339;
  reg [7:0] _T_4368_16; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_340;
  reg [7:0] _T_4368_17; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_341;
  reg [7:0] _T_4368_18; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_342;
  reg [7:0] _T_4368_19; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_343;
  reg [7:0] _T_4368_20; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_344;
  reg [7:0] _T_4368_21; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_345;
  reg [7:0] _T_4368_22; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_346;
  reg [7:0] _T_4368_23; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_347;
  reg [7:0] _T_4368_24; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_348;
  reg [7:0] _T_4368_25; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_349;
  reg [7:0] _T_4368_26; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_350;
  reg [7:0] _T_4368_27; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_351;
  reg [7:0] _T_4368_28; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_352;
  reg [7:0] _T_4368_29; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_353;
  reg [7:0] _T_4368_30; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_354;
  reg [7:0] _T_4368_31; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_355;
  reg [7:0] _T_4368_32; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_356;
  reg [7:0] _T_4368_33; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_357;
  reg [7:0] _T_4368_34; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_358;
  reg [7:0] _T_4368_35; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_359;
  reg [7:0] _T_4368_36; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_360;
  reg [7:0] _T_4368_37; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_361;
  reg [7:0] _T_4368_38; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_362;
  reg [7:0] _T_4368_39; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_363;
  reg [7:0] _T_4368_40; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_364;
  reg [7:0] _T_4368_41; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_365;
  reg [7:0] _T_4368_42; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_366;
  reg [7:0] _T_4368_43; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_367;
  reg [7:0] _T_4368_44; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_368;
  reg [7:0] _T_4368_45; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_369;
  reg [7:0] _T_4368_46; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_370;
  reg [7:0] _T_4368_47; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_371;
  reg [7:0] _T_4368_48; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_372;
  reg [7:0] _T_4368_49; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_373;
  reg [7:0] _T_4368_50; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_374;
  reg [7:0] _T_4368_51; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_375;
  reg [7:0] _T_4368_52; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_376;
  reg [7:0] _T_4368_53; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_377;
  reg [7:0] _T_4368_54; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_378;
  reg [7:0] _T_4368_55; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_379;
  reg [7:0] _T_4368_56; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_380;
  reg [7:0] _T_4368_57; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_381;
  reg [7:0] _T_4368_58; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_382;
  reg [7:0] _T_4368_59; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_383;
  reg [7:0] _T_4368_60; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_384;
  reg [7:0] _T_4368_61; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_385;
  reg [7:0] _T_4368_62; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_386;
  reg [7:0] _T_4368_63; // @[retiming.scala 9:92:@153.4]
  reg [31:0] _RAND_387;
  reg  _T_4771_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_388;
  reg  _T_4771_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_389;
  reg  _T_4771_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_390;
  reg  _T_4771_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_391;
  reg  _T_4771_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_392;
  reg  _T_4771_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_393;
  reg  _T_4771_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_394;
  reg  _T_4771_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_395;
  reg  _T_4771_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_396;
  reg  _T_4771_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_397;
  reg  _T_4771_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_398;
  reg  _T_4771_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_399;
  reg  _T_4771_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_400;
  reg  _T_4771_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_401;
  reg  _T_4771_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_402;
  reg  _T_4771_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_403;
  reg  _T_4771_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_404;
  reg  _T_4771_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_405;
  reg  _T_4771_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_406;
  reg  _T_4771_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_407;
  reg  _T_4771_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_408;
  reg  _T_4771_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_409;
  reg  _T_4771_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_410;
  reg  _T_4771_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_411;
  reg  _T_4771_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_412;
  reg  _T_4771_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_413;
  reg  _T_4771_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_414;
  reg  _T_4771_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_415;
  reg  _T_4771_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_416;
  reg  _T_4771_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_417;
  reg  _T_4771_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_418;
  reg  _T_4771_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_419;
  reg  _T_4771_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_420;
  reg  _T_4771_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_421;
  reg  _T_4771_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_422;
  reg  _T_4771_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_423;
  reg  _T_4771_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_424;
  reg  _T_4771_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_425;
  reg  _T_4771_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_426;
  reg  _T_4771_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_427;
  reg  _T_4771_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_428;
  reg  _T_4771_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_429;
  reg  _T_4771_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_430;
  reg  _T_4771_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_431;
  reg  _T_4771_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_432;
  reg  _T_4771_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_433;
  reg  _T_4771_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_434;
  reg  _T_4771_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_435;
  reg  _T_4771_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_436;
  reg  _T_4771_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_437;
  reg  _T_4771_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_438;
  reg  _T_4771_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_439;
  reg  _T_4771_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_440;
  reg  _T_4771_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_441;
  reg  _T_4771_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_442;
  reg  _T_4771_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_443;
  reg  _T_4771_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_444;
  reg  _T_4771_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_445;
  reg  _T_4771_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_446;
  reg  _T_4771_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_447;
  reg  _T_4771_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_448;
  reg  _T_4771_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_449;
  reg  _T_4771_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_450;
  reg  _T_4771_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@220.4]
  reg [31:0] _RAND_451;
  reg  _T_5234_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_452;
  reg  _T_5234_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_453;
  reg  _T_5234_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_454;
  reg  _T_5234_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_455;
  reg  _T_5234_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_456;
  reg  _T_5234_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_457;
  reg  _T_5234_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_458;
  reg  _T_5234_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_459;
  reg  _T_5234_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_460;
  reg  _T_5234_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_461;
  reg  _T_5234_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_462;
  reg  _T_5234_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_463;
  reg  _T_5234_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_464;
  reg  _T_5234_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_465;
  reg  _T_5234_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_466;
  reg  _T_5234_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_467;
  reg  _T_5234_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_468;
  reg  _T_5234_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_469;
  reg  _T_5234_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_470;
  reg  _T_5234_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_471;
  reg  _T_5234_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_472;
  reg  _T_5234_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_473;
  reg  _T_5234_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_474;
  reg  _T_5234_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_475;
  reg  _T_5234_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_476;
  reg  _T_5234_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_477;
  reg  _T_5234_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_478;
  reg  _T_5234_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_479;
  reg  _T_5234_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_480;
  reg  _T_5234_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_481;
  reg  _T_5234_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_482;
  reg  _T_5234_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_483;
  reg  _T_5234_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_484;
  reg  _T_5234_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_485;
  reg  _T_5234_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_486;
  reg  _T_5234_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_487;
  reg  _T_5234_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_488;
  reg  _T_5234_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_489;
  reg  _T_5234_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_490;
  reg  _T_5234_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_491;
  reg  _T_5234_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_492;
  reg  _T_5234_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_493;
  reg  _T_5234_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_494;
  reg  _T_5234_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_495;
  reg  _T_5234_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_496;
  reg  _T_5234_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_497;
  reg  _T_5234_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_498;
  reg  _T_5234_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_499;
  reg  _T_5234_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_500;
  reg  _T_5234_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_501;
  reg  _T_5234_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_502;
  reg  _T_5234_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_503;
  reg  _T_5234_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_504;
  reg  _T_5234_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_505;
  reg  _T_5234_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_506;
  reg  _T_5234_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_507;
  reg  _T_5234_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_508;
  reg  _T_5234_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_509;
  reg  _T_5234_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_510;
  reg  _T_5234_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_511;
  reg  _T_5234_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_512;
  reg  _T_5234_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_513;
  reg  _T_5234_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_514;
  reg  _T_5234_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 59:70:@286.4]
  reg [31:0] _RAND_515;
  reg  _T_5435; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 61:70:@288.4]
  reg [31:0] _RAND_516;
  reg  _T_5438; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 61:70:@289.4]
  reg [31:0] _RAND_517;
  reg  _T_5535_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@308.4]
  reg [31:0] _RAND_518;
  reg  _T_5535_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@308.4]
  reg [31:0] _RAND_519;
  reg  _T_5535_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@308.4]
  reg [31:0] _RAND_520;
  reg  _T_5535_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@308.4]
  reg [31:0] _RAND_521;
  reg  _T_5535_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@308.4]
  reg [31:0] _RAND_522;
  reg  _T_5535_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@308.4]
  reg [31:0] _RAND_523;
  reg  _T_5535_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@308.4]
  reg [31:0] _RAND_524;
  reg  _T_5535_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@308.4]
  reg [31:0] _RAND_525;
  reg  _T_5535_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@308.4]
  reg [31:0] _RAND_526;
  reg  _T_5535_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@308.4]
  reg [31:0] _RAND_527;
  reg  _T_5535_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@308.4]
  reg [31:0] _RAND_528;
  reg  _T_5535_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@308.4]
  reg [31:0] _RAND_529;
  reg  _T_5535_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@308.4]
  reg [31:0] _RAND_530;
  reg  _T_5535_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@308.4]
  reg [31:0] _RAND_531;
  reg  _T_5535_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@308.4]
  reg [31:0] _RAND_532;
  reg  _T_5535_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@308.4]
  reg [31:0] _RAND_533;
  reg  _T_5662_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@326.4]
  reg [31:0] _RAND_534;
  reg  _T_5662_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@326.4]
  reg [31:0] _RAND_535;
  reg  _T_5662_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@326.4]
  reg [31:0] _RAND_536;
  reg  _T_5662_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@326.4]
  reg [31:0] _RAND_537;
  reg  _T_5662_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@326.4]
  reg [31:0] _RAND_538;
  reg  _T_5662_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@326.4]
  reg [31:0] _RAND_539;
  reg  _T_5662_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@326.4]
  reg [31:0] _RAND_540;
  reg  _T_5662_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@326.4]
  reg [31:0] _RAND_541;
  reg  _T_5662_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@326.4]
  reg [31:0] _RAND_542;
  reg  _T_5662_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@326.4]
  reg [31:0] _RAND_543;
  reg  _T_5662_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@326.4]
  reg [31:0] _RAND_544;
  reg  _T_5662_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@326.4]
  reg [31:0] _RAND_545;
  reg  _T_5662_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@326.4]
  reg [31:0] _RAND_546;
  reg  _T_5662_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@326.4]
  reg [31:0] _RAND_547;
  reg  _T_5662_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@326.4]
  reg [31:0] _RAND_548;
  reg  _T_5662_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 63:70:@326.4]
  reg [31:0] _RAND_549;
  wire  _T_5715; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:33:@603.4]
  wire  _GEN_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _GEN_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire [8:0] _GEN_64; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  wire  _T_5716; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:32:@672.4]
  wire  _GEN_65; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_66; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_67; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_68; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_69; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_70; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_71; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_72; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_73; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_74; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_75; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_76; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_77; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_78; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_79; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_80; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_81; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_82; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_83; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_84; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_85; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_86; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_87; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_88; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_89; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_90; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_91; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_92; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_93; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_94; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_95; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_96; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_97; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_98; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_99; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_100; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_101; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_102; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_103; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_104; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_105; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_106; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_107; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_108; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_109; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_110; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_111; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_112; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_113; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_114; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_115; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_116; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_117; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_118; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_119; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_120; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_121; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_122; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_123; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_124; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_125; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_126; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_127; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_128; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_129; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_130; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_131; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_132; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_133; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_134; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_135; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_136; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_137; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_138; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_139; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_140; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_141; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_142; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_143; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _GEN_144; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  wire  _T_5717; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:33:@1140.4]
  wire  _GEN_273; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_274; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_275; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_276; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_277; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_278; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_279; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_280; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_281; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_282; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_283; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_284; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_285; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_286; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_287; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_288; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_289; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_290; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_291; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_292; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_293; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_294; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_295; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_296; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_297; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_298; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_299; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_300; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_301; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_302; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_303; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_304; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_305; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_306; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_307; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_308; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_309; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_310; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_311; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_312; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_313; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_314; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_315; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_316; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_317; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_318; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_319; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_320; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_321; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_322; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_323; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_324; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_325; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_326; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_327; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_328; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_329; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_330; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_331; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_332; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_333; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_334; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_335; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _GEN_336; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire [8:0] _GEN_337; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  wire  _T_5718; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:32:@1209.4]
  wire  _GEN_338; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_339; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_340; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_341; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_342; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_343; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_344; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_345; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_346; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_347; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_348; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_349; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_350; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_351; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_352; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_353; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_354; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_355; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_356; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_357; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_358; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_359; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_360; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_361; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_362; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_363; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_364; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_365; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_366; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_367; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_368; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_369; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_370; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_371; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_372; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_373; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_374; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_375; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_376; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_377; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_378; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_379; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_380; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_381; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_382; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_383; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_384; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_385; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_386; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_387; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_388; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_389; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_390; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_391; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_392; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_393; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_394; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_395; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_396; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_397; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_398; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_399; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_400; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_401; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_402; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_403; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_404; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_405; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_406; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_407; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_408; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_409; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_410; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_411; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_412; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_413; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_414; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_415; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_416; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  wire  _GEN_417; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _T_3014 = io_nvdla_core_rstn == 1'h0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 45:38:@8.4]
  assign _T_5715 = io_sc2mac_dat_valid | _T_4219; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:33:@603.4]
  assign _GEN_0 = _T_5715 ? io_sc2mac_dat_bits_mask_0 : _T_3555_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_1 = _T_5715 ? io_sc2mac_dat_bits_mask_1 : _T_3555_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_2 = _T_5715 ? io_sc2mac_dat_bits_mask_2 : _T_3555_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_3 = _T_5715 ? io_sc2mac_dat_bits_mask_3 : _T_3555_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_4 = _T_5715 ? io_sc2mac_dat_bits_mask_4 : _T_3555_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_5 = _T_5715 ? io_sc2mac_dat_bits_mask_5 : _T_3555_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_6 = _T_5715 ? io_sc2mac_dat_bits_mask_6 : _T_3555_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_7 = _T_5715 ? io_sc2mac_dat_bits_mask_7 : _T_3555_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_8 = _T_5715 ? io_sc2mac_dat_bits_mask_8 : _T_3555_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_9 = _T_5715 ? io_sc2mac_dat_bits_mask_9 : _T_3555_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_10 = _T_5715 ? io_sc2mac_dat_bits_mask_10 : _T_3555_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_11 = _T_5715 ? io_sc2mac_dat_bits_mask_11 : _T_3555_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_12 = _T_5715 ? io_sc2mac_dat_bits_mask_12 : _T_3555_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_13 = _T_5715 ? io_sc2mac_dat_bits_mask_13 : _T_3555_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_14 = _T_5715 ? io_sc2mac_dat_bits_mask_14 : _T_3555_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_15 = _T_5715 ? io_sc2mac_dat_bits_mask_15 : _T_3555_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_16 = _T_5715 ? io_sc2mac_dat_bits_mask_16 : _T_3555_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_17 = _T_5715 ? io_sc2mac_dat_bits_mask_17 : _T_3555_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_18 = _T_5715 ? io_sc2mac_dat_bits_mask_18 : _T_3555_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_19 = _T_5715 ? io_sc2mac_dat_bits_mask_19 : _T_3555_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_20 = _T_5715 ? io_sc2mac_dat_bits_mask_20 : _T_3555_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_21 = _T_5715 ? io_sc2mac_dat_bits_mask_21 : _T_3555_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_22 = _T_5715 ? io_sc2mac_dat_bits_mask_22 : _T_3555_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_23 = _T_5715 ? io_sc2mac_dat_bits_mask_23 : _T_3555_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_24 = _T_5715 ? io_sc2mac_dat_bits_mask_24 : _T_3555_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_25 = _T_5715 ? io_sc2mac_dat_bits_mask_25 : _T_3555_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_26 = _T_5715 ? io_sc2mac_dat_bits_mask_26 : _T_3555_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_27 = _T_5715 ? io_sc2mac_dat_bits_mask_27 : _T_3555_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_28 = _T_5715 ? io_sc2mac_dat_bits_mask_28 : _T_3555_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_29 = _T_5715 ? io_sc2mac_dat_bits_mask_29 : _T_3555_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_30 = _T_5715 ? io_sc2mac_dat_bits_mask_30 : _T_3555_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_31 = _T_5715 ? io_sc2mac_dat_bits_mask_31 : _T_3555_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_32 = _T_5715 ? io_sc2mac_dat_bits_mask_32 : _T_3555_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_33 = _T_5715 ? io_sc2mac_dat_bits_mask_33 : _T_3555_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_34 = _T_5715 ? io_sc2mac_dat_bits_mask_34 : _T_3555_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_35 = _T_5715 ? io_sc2mac_dat_bits_mask_35 : _T_3555_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_36 = _T_5715 ? io_sc2mac_dat_bits_mask_36 : _T_3555_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_37 = _T_5715 ? io_sc2mac_dat_bits_mask_37 : _T_3555_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_38 = _T_5715 ? io_sc2mac_dat_bits_mask_38 : _T_3555_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_39 = _T_5715 ? io_sc2mac_dat_bits_mask_39 : _T_3555_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_40 = _T_5715 ? io_sc2mac_dat_bits_mask_40 : _T_3555_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_41 = _T_5715 ? io_sc2mac_dat_bits_mask_41 : _T_3555_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_42 = _T_5715 ? io_sc2mac_dat_bits_mask_42 : _T_3555_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_43 = _T_5715 ? io_sc2mac_dat_bits_mask_43 : _T_3555_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_44 = _T_5715 ? io_sc2mac_dat_bits_mask_44 : _T_3555_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_45 = _T_5715 ? io_sc2mac_dat_bits_mask_45 : _T_3555_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_46 = _T_5715 ? io_sc2mac_dat_bits_mask_46 : _T_3555_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_47 = _T_5715 ? io_sc2mac_dat_bits_mask_47 : _T_3555_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_48 = _T_5715 ? io_sc2mac_dat_bits_mask_48 : _T_3555_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_49 = _T_5715 ? io_sc2mac_dat_bits_mask_49 : _T_3555_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_50 = _T_5715 ? io_sc2mac_dat_bits_mask_50 : _T_3555_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_51 = _T_5715 ? io_sc2mac_dat_bits_mask_51 : _T_3555_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_52 = _T_5715 ? io_sc2mac_dat_bits_mask_52 : _T_3555_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_53 = _T_5715 ? io_sc2mac_dat_bits_mask_53 : _T_3555_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_54 = _T_5715 ? io_sc2mac_dat_bits_mask_54 : _T_3555_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_55 = _T_5715 ? io_sc2mac_dat_bits_mask_55 : _T_3555_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_56 = _T_5715 ? io_sc2mac_dat_bits_mask_56 : _T_3555_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_57 = _T_5715 ? io_sc2mac_dat_bits_mask_57 : _T_3555_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_58 = _T_5715 ? io_sc2mac_dat_bits_mask_58 : _T_3555_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_59 = _T_5715 ? io_sc2mac_dat_bits_mask_59 : _T_3555_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_60 = _T_5715 ? io_sc2mac_dat_bits_mask_60 : _T_3555_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_61 = _T_5715 ? io_sc2mac_dat_bits_mask_61 : _T_3555_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_62 = _T_5715 ? io_sc2mac_dat_bits_mask_62 : _T_3555_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_63 = _T_5715 ? io_sc2mac_dat_bits_mask_63 : _T_3555_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _GEN_64 = _T_5715 ? io_sc2mac_dat_bits_pd : _T_4227; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@604.4]
  assign _T_5716 = io_sc2mac_wt_valid | _T_5435; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:32:@672.4]
  assign _GEN_65 = _T_5716 ? io_sc2mac_wt_bits_mask_0 : _T_4771_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_66 = _T_5716 ? io_sc2mac_wt_bits_mask_1 : _T_4771_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_67 = _T_5716 ? io_sc2mac_wt_bits_mask_2 : _T_4771_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_68 = _T_5716 ? io_sc2mac_wt_bits_mask_3 : _T_4771_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_69 = _T_5716 ? io_sc2mac_wt_bits_mask_4 : _T_4771_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_70 = _T_5716 ? io_sc2mac_wt_bits_mask_5 : _T_4771_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_71 = _T_5716 ? io_sc2mac_wt_bits_mask_6 : _T_4771_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_72 = _T_5716 ? io_sc2mac_wt_bits_mask_7 : _T_4771_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_73 = _T_5716 ? io_sc2mac_wt_bits_mask_8 : _T_4771_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_74 = _T_5716 ? io_sc2mac_wt_bits_mask_9 : _T_4771_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_75 = _T_5716 ? io_sc2mac_wt_bits_mask_10 : _T_4771_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_76 = _T_5716 ? io_sc2mac_wt_bits_mask_11 : _T_4771_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_77 = _T_5716 ? io_sc2mac_wt_bits_mask_12 : _T_4771_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_78 = _T_5716 ? io_sc2mac_wt_bits_mask_13 : _T_4771_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_79 = _T_5716 ? io_sc2mac_wt_bits_mask_14 : _T_4771_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_80 = _T_5716 ? io_sc2mac_wt_bits_mask_15 : _T_4771_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_81 = _T_5716 ? io_sc2mac_wt_bits_mask_16 : _T_4771_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_82 = _T_5716 ? io_sc2mac_wt_bits_mask_17 : _T_4771_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_83 = _T_5716 ? io_sc2mac_wt_bits_mask_18 : _T_4771_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_84 = _T_5716 ? io_sc2mac_wt_bits_mask_19 : _T_4771_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_85 = _T_5716 ? io_sc2mac_wt_bits_mask_20 : _T_4771_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_86 = _T_5716 ? io_sc2mac_wt_bits_mask_21 : _T_4771_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_87 = _T_5716 ? io_sc2mac_wt_bits_mask_22 : _T_4771_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_88 = _T_5716 ? io_sc2mac_wt_bits_mask_23 : _T_4771_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_89 = _T_5716 ? io_sc2mac_wt_bits_mask_24 : _T_4771_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_90 = _T_5716 ? io_sc2mac_wt_bits_mask_25 : _T_4771_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_91 = _T_5716 ? io_sc2mac_wt_bits_mask_26 : _T_4771_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_92 = _T_5716 ? io_sc2mac_wt_bits_mask_27 : _T_4771_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_93 = _T_5716 ? io_sc2mac_wt_bits_mask_28 : _T_4771_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_94 = _T_5716 ? io_sc2mac_wt_bits_mask_29 : _T_4771_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_95 = _T_5716 ? io_sc2mac_wt_bits_mask_30 : _T_4771_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_96 = _T_5716 ? io_sc2mac_wt_bits_mask_31 : _T_4771_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_97 = _T_5716 ? io_sc2mac_wt_bits_mask_32 : _T_4771_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_98 = _T_5716 ? io_sc2mac_wt_bits_mask_33 : _T_4771_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_99 = _T_5716 ? io_sc2mac_wt_bits_mask_34 : _T_4771_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_100 = _T_5716 ? io_sc2mac_wt_bits_mask_35 : _T_4771_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_101 = _T_5716 ? io_sc2mac_wt_bits_mask_36 : _T_4771_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_102 = _T_5716 ? io_sc2mac_wt_bits_mask_37 : _T_4771_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_103 = _T_5716 ? io_sc2mac_wt_bits_mask_38 : _T_4771_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_104 = _T_5716 ? io_sc2mac_wt_bits_mask_39 : _T_4771_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_105 = _T_5716 ? io_sc2mac_wt_bits_mask_40 : _T_4771_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_106 = _T_5716 ? io_sc2mac_wt_bits_mask_41 : _T_4771_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_107 = _T_5716 ? io_sc2mac_wt_bits_mask_42 : _T_4771_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_108 = _T_5716 ? io_sc2mac_wt_bits_mask_43 : _T_4771_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_109 = _T_5716 ? io_sc2mac_wt_bits_mask_44 : _T_4771_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_110 = _T_5716 ? io_sc2mac_wt_bits_mask_45 : _T_4771_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_111 = _T_5716 ? io_sc2mac_wt_bits_mask_46 : _T_4771_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_112 = _T_5716 ? io_sc2mac_wt_bits_mask_47 : _T_4771_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_113 = _T_5716 ? io_sc2mac_wt_bits_mask_48 : _T_4771_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_114 = _T_5716 ? io_sc2mac_wt_bits_mask_49 : _T_4771_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_115 = _T_5716 ? io_sc2mac_wt_bits_mask_50 : _T_4771_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_116 = _T_5716 ? io_sc2mac_wt_bits_mask_51 : _T_4771_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_117 = _T_5716 ? io_sc2mac_wt_bits_mask_52 : _T_4771_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_118 = _T_5716 ? io_sc2mac_wt_bits_mask_53 : _T_4771_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_119 = _T_5716 ? io_sc2mac_wt_bits_mask_54 : _T_4771_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_120 = _T_5716 ? io_sc2mac_wt_bits_mask_55 : _T_4771_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_121 = _T_5716 ? io_sc2mac_wt_bits_mask_56 : _T_4771_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_122 = _T_5716 ? io_sc2mac_wt_bits_mask_57 : _T_4771_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_123 = _T_5716 ? io_sc2mac_wt_bits_mask_58 : _T_4771_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_124 = _T_5716 ? io_sc2mac_wt_bits_mask_59 : _T_4771_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_125 = _T_5716 ? io_sc2mac_wt_bits_mask_60 : _T_4771_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_126 = _T_5716 ? io_sc2mac_wt_bits_mask_61 : _T_4771_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_127 = _T_5716 ? io_sc2mac_wt_bits_mask_62 : _T_4771_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_128 = _T_5716 ? io_sc2mac_wt_bits_mask_63 : _T_4771_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_129 = _T_5716 ? io_sc2mac_wt_bits_sel_0 : _T_5535_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_130 = _T_5716 ? io_sc2mac_wt_bits_sel_1 : _T_5535_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_131 = _T_5716 ? io_sc2mac_wt_bits_sel_2 : _T_5535_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_132 = _T_5716 ? io_sc2mac_wt_bits_sel_3 : _T_5535_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_133 = _T_5716 ? io_sc2mac_wt_bits_sel_4 : _T_5535_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_134 = _T_5716 ? io_sc2mac_wt_bits_sel_5 : _T_5535_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_135 = _T_5716 ? io_sc2mac_wt_bits_sel_6 : _T_5535_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_136 = _T_5716 ? io_sc2mac_wt_bits_sel_7 : _T_5535_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_137 = _T_5716 ? io_sc2mac_wt_bits_sel_8 : _T_5535_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_138 = _T_5716 ? io_sc2mac_wt_bits_sel_9 : _T_5535_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_139 = _T_5716 ? io_sc2mac_wt_bits_sel_10 : _T_5535_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_140 = _T_5716 ? io_sc2mac_wt_bits_sel_11 : _T_5535_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_141 = _T_5716 ? io_sc2mac_wt_bits_sel_12 : _T_5535_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_142 = _T_5716 ? io_sc2mac_wt_bits_sel_13 : _T_5535_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_143 = _T_5716 ? io_sc2mac_wt_bits_sel_14 : _T_5535_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _GEN_144 = _T_5716 ? io_sc2mac_wt_bits_sel_15 : _T_5535_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@673.4]
  assign _T_5717 = _T_4219 | _T_4222; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:33:@1140.4]
  assign _GEN_273 = _T_5717 ? _T_3555_0 : _T_4018_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_274 = _T_5717 ? _T_3555_1 : _T_4018_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_275 = _T_5717 ? _T_3555_2 : _T_4018_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_276 = _T_5717 ? _T_3555_3 : _T_4018_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_277 = _T_5717 ? _T_3555_4 : _T_4018_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_278 = _T_5717 ? _T_3555_5 : _T_4018_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_279 = _T_5717 ? _T_3555_6 : _T_4018_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_280 = _T_5717 ? _T_3555_7 : _T_4018_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_281 = _T_5717 ? _T_3555_8 : _T_4018_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_282 = _T_5717 ? _T_3555_9 : _T_4018_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_283 = _T_5717 ? _T_3555_10 : _T_4018_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_284 = _T_5717 ? _T_3555_11 : _T_4018_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_285 = _T_5717 ? _T_3555_12 : _T_4018_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_286 = _T_5717 ? _T_3555_13 : _T_4018_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_287 = _T_5717 ? _T_3555_14 : _T_4018_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_288 = _T_5717 ? _T_3555_15 : _T_4018_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_289 = _T_5717 ? _T_3555_16 : _T_4018_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_290 = _T_5717 ? _T_3555_17 : _T_4018_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_291 = _T_5717 ? _T_3555_18 : _T_4018_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_292 = _T_5717 ? _T_3555_19 : _T_4018_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_293 = _T_5717 ? _T_3555_20 : _T_4018_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_294 = _T_5717 ? _T_3555_21 : _T_4018_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_295 = _T_5717 ? _T_3555_22 : _T_4018_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_296 = _T_5717 ? _T_3555_23 : _T_4018_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_297 = _T_5717 ? _T_3555_24 : _T_4018_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_298 = _T_5717 ? _T_3555_25 : _T_4018_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_299 = _T_5717 ? _T_3555_26 : _T_4018_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_300 = _T_5717 ? _T_3555_27 : _T_4018_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_301 = _T_5717 ? _T_3555_28 : _T_4018_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_302 = _T_5717 ? _T_3555_29 : _T_4018_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_303 = _T_5717 ? _T_3555_30 : _T_4018_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_304 = _T_5717 ? _T_3555_31 : _T_4018_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_305 = _T_5717 ? _T_3555_32 : _T_4018_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_306 = _T_5717 ? _T_3555_33 : _T_4018_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_307 = _T_5717 ? _T_3555_34 : _T_4018_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_308 = _T_5717 ? _T_3555_35 : _T_4018_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_309 = _T_5717 ? _T_3555_36 : _T_4018_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_310 = _T_5717 ? _T_3555_37 : _T_4018_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_311 = _T_5717 ? _T_3555_38 : _T_4018_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_312 = _T_5717 ? _T_3555_39 : _T_4018_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_313 = _T_5717 ? _T_3555_40 : _T_4018_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_314 = _T_5717 ? _T_3555_41 : _T_4018_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_315 = _T_5717 ? _T_3555_42 : _T_4018_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_316 = _T_5717 ? _T_3555_43 : _T_4018_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_317 = _T_5717 ? _T_3555_44 : _T_4018_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_318 = _T_5717 ? _T_3555_45 : _T_4018_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_319 = _T_5717 ? _T_3555_46 : _T_4018_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_320 = _T_5717 ? _T_3555_47 : _T_4018_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_321 = _T_5717 ? _T_3555_48 : _T_4018_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_322 = _T_5717 ? _T_3555_49 : _T_4018_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_323 = _T_5717 ? _T_3555_50 : _T_4018_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_324 = _T_5717 ? _T_3555_51 : _T_4018_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_325 = _T_5717 ? _T_3555_52 : _T_4018_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_326 = _T_5717 ? _T_3555_53 : _T_4018_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_327 = _T_5717 ? _T_3555_54 : _T_4018_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_328 = _T_5717 ? _T_3555_55 : _T_4018_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_329 = _T_5717 ? _T_3555_56 : _T_4018_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_330 = _T_5717 ? _T_3555_57 : _T_4018_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_331 = _T_5717 ? _T_3555_58 : _T_4018_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_332 = _T_5717 ? _T_3555_59 : _T_4018_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_333 = _T_5717 ? _T_3555_60 : _T_4018_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_334 = _T_5717 ? _T_3555_61 : _T_4018_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_335 = _T_5717 ? _T_3555_62 : _T_4018_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_336 = _T_5717 ? _T_3555_63 : _T_4018_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _GEN_337 = _T_5717 ? _T_4227 : _T_4230; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 81:56:@1141.4]
  assign _T_5718 = _T_5435 | _T_5438; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:32:@1209.4]
  assign _GEN_338 = _T_5718 ? _T_4771_0 : _T_5234_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_339 = _T_5718 ? _T_4771_1 : _T_5234_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_340 = _T_5718 ? _T_4771_2 : _T_5234_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_341 = _T_5718 ? _T_4771_3 : _T_5234_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_342 = _T_5718 ? _T_4771_4 : _T_5234_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_343 = _T_5718 ? _T_4771_5 : _T_5234_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_344 = _T_5718 ? _T_4771_6 : _T_5234_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_345 = _T_5718 ? _T_4771_7 : _T_5234_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_346 = _T_5718 ? _T_4771_8 : _T_5234_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_347 = _T_5718 ? _T_4771_9 : _T_5234_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_348 = _T_5718 ? _T_4771_10 : _T_5234_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_349 = _T_5718 ? _T_4771_11 : _T_5234_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_350 = _T_5718 ? _T_4771_12 : _T_5234_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_351 = _T_5718 ? _T_4771_13 : _T_5234_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_352 = _T_5718 ? _T_4771_14 : _T_5234_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_353 = _T_5718 ? _T_4771_15 : _T_5234_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_354 = _T_5718 ? _T_4771_16 : _T_5234_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_355 = _T_5718 ? _T_4771_17 : _T_5234_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_356 = _T_5718 ? _T_4771_18 : _T_5234_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_357 = _T_5718 ? _T_4771_19 : _T_5234_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_358 = _T_5718 ? _T_4771_20 : _T_5234_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_359 = _T_5718 ? _T_4771_21 : _T_5234_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_360 = _T_5718 ? _T_4771_22 : _T_5234_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_361 = _T_5718 ? _T_4771_23 : _T_5234_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_362 = _T_5718 ? _T_4771_24 : _T_5234_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_363 = _T_5718 ? _T_4771_25 : _T_5234_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_364 = _T_5718 ? _T_4771_26 : _T_5234_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_365 = _T_5718 ? _T_4771_27 : _T_5234_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_366 = _T_5718 ? _T_4771_28 : _T_5234_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_367 = _T_5718 ? _T_4771_29 : _T_5234_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_368 = _T_5718 ? _T_4771_30 : _T_5234_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_369 = _T_5718 ? _T_4771_31 : _T_5234_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_370 = _T_5718 ? _T_4771_32 : _T_5234_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_371 = _T_5718 ? _T_4771_33 : _T_5234_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_372 = _T_5718 ? _T_4771_34 : _T_5234_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_373 = _T_5718 ? _T_4771_35 : _T_5234_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_374 = _T_5718 ? _T_4771_36 : _T_5234_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_375 = _T_5718 ? _T_4771_37 : _T_5234_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_376 = _T_5718 ? _T_4771_38 : _T_5234_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_377 = _T_5718 ? _T_4771_39 : _T_5234_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_378 = _T_5718 ? _T_4771_40 : _T_5234_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_379 = _T_5718 ? _T_4771_41 : _T_5234_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_380 = _T_5718 ? _T_4771_42 : _T_5234_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_381 = _T_5718 ? _T_4771_43 : _T_5234_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_382 = _T_5718 ? _T_4771_44 : _T_5234_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_383 = _T_5718 ? _T_4771_45 : _T_5234_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_384 = _T_5718 ? _T_4771_46 : _T_5234_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_385 = _T_5718 ? _T_4771_47 : _T_5234_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_386 = _T_5718 ? _T_4771_48 : _T_5234_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_387 = _T_5718 ? _T_4771_49 : _T_5234_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_388 = _T_5718 ? _T_4771_50 : _T_5234_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_389 = _T_5718 ? _T_4771_51 : _T_5234_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_390 = _T_5718 ? _T_4771_52 : _T_5234_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_391 = _T_5718 ? _T_4771_53 : _T_5234_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_392 = _T_5718 ? _T_4771_54 : _T_5234_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_393 = _T_5718 ? _T_4771_55 : _T_5234_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_394 = _T_5718 ? _T_4771_56 : _T_5234_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_395 = _T_5718 ? _T_4771_57 : _T_5234_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_396 = _T_5718 ? _T_4771_58 : _T_5234_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_397 = _T_5718 ? _T_4771_59 : _T_5234_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_398 = _T_5718 ? _T_4771_60 : _T_5234_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_399 = _T_5718 ? _T_4771_61 : _T_5234_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_400 = _T_5718 ? _T_4771_62 : _T_5234_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_401 = _T_5718 ? _T_4771_63 : _T_5234_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_402 = _T_5718 ? _T_5535_0 : _T_5662_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_403 = _T_5718 ? _T_5535_1 : _T_5662_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_404 = _T_5718 ? _T_5535_2 : _T_5662_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_405 = _T_5718 ? _T_5535_3 : _T_5662_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_406 = _T_5718 ? _T_5535_4 : _T_5662_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_407 = _T_5718 ? _T_5535_5 : _T_5662_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_408 = _T_5718 ? _T_5535_6 : _T_5662_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_409 = _T_5718 ? _T_5535_7 : _T_5662_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_410 = _T_5718 ? _T_5535_8 : _T_5662_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_411 = _T_5718 ? _T_5535_9 : _T_5662_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_412 = _T_5718 ? _T_5535_10 : _T_5662_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_413 = _T_5718 ? _T_5535_11 : _T_5662_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_414 = _T_5718 ? _T_5535_12 : _T_5662_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_415 = _T_5718 ? _T_5535_13 : _T_5662_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_416 = _T_5718 ? _T_5535_14 : _T_5662_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign _GEN_417 = _T_5718 ? _T_5535_15 : _T_5662_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 87:54:@1210.4]
  assign io_in_dat_valid = _T_4222; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 103:21:@1676.4]
  assign io_in_dat_bits_mask_0 = _T_4018_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1677.4]
  assign io_in_dat_bits_mask_1 = _T_4018_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1678.4]
  assign io_in_dat_bits_mask_2 = _T_4018_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1679.4]
  assign io_in_dat_bits_mask_3 = _T_4018_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1680.4]
  assign io_in_dat_bits_mask_4 = _T_4018_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1681.4]
  assign io_in_dat_bits_mask_5 = _T_4018_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1682.4]
  assign io_in_dat_bits_mask_6 = _T_4018_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1683.4]
  assign io_in_dat_bits_mask_7 = _T_4018_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1684.4]
  assign io_in_dat_bits_mask_8 = _T_4018_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1685.4]
  assign io_in_dat_bits_mask_9 = _T_4018_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1686.4]
  assign io_in_dat_bits_mask_10 = _T_4018_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1687.4]
  assign io_in_dat_bits_mask_11 = _T_4018_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1688.4]
  assign io_in_dat_bits_mask_12 = _T_4018_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1689.4]
  assign io_in_dat_bits_mask_13 = _T_4018_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1690.4]
  assign io_in_dat_bits_mask_14 = _T_4018_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1691.4]
  assign io_in_dat_bits_mask_15 = _T_4018_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1692.4]
  assign io_in_dat_bits_mask_16 = _T_4018_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1693.4]
  assign io_in_dat_bits_mask_17 = _T_4018_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1694.4]
  assign io_in_dat_bits_mask_18 = _T_4018_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1695.4]
  assign io_in_dat_bits_mask_19 = _T_4018_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1696.4]
  assign io_in_dat_bits_mask_20 = _T_4018_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1697.4]
  assign io_in_dat_bits_mask_21 = _T_4018_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1698.4]
  assign io_in_dat_bits_mask_22 = _T_4018_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1699.4]
  assign io_in_dat_bits_mask_23 = _T_4018_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1700.4]
  assign io_in_dat_bits_mask_24 = _T_4018_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1701.4]
  assign io_in_dat_bits_mask_25 = _T_4018_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1702.4]
  assign io_in_dat_bits_mask_26 = _T_4018_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1703.4]
  assign io_in_dat_bits_mask_27 = _T_4018_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1704.4]
  assign io_in_dat_bits_mask_28 = _T_4018_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1705.4]
  assign io_in_dat_bits_mask_29 = _T_4018_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1706.4]
  assign io_in_dat_bits_mask_30 = _T_4018_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1707.4]
  assign io_in_dat_bits_mask_31 = _T_4018_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1708.4]
  assign io_in_dat_bits_mask_32 = _T_4018_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1709.4]
  assign io_in_dat_bits_mask_33 = _T_4018_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1710.4]
  assign io_in_dat_bits_mask_34 = _T_4018_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1711.4]
  assign io_in_dat_bits_mask_35 = _T_4018_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1712.4]
  assign io_in_dat_bits_mask_36 = _T_4018_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1713.4]
  assign io_in_dat_bits_mask_37 = _T_4018_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1714.4]
  assign io_in_dat_bits_mask_38 = _T_4018_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1715.4]
  assign io_in_dat_bits_mask_39 = _T_4018_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1716.4]
  assign io_in_dat_bits_mask_40 = _T_4018_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1717.4]
  assign io_in_dat_bits_mask_41 = _T_4018_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1718.4]
  assign io_in_dat_bits_mask_42 = _T_4018_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1719.4]
  assign io_in_dat_bits_mask_43 = _T_4018_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1720.4]
  assign io_in_dat_bits_mask_44 = _T_4018_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1721.4]
  assign io_in_dat_bits_mask_45 = _T_4018_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1722.4]
  assign io_in_dat_bits_mask_46 = _T_4018_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1723.4]
  assign io_in_dat_bits_mask_47 = _T_4018_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1724.4]
  assign io_in_dat_bits_mask_48 = _T_4018_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1725.4]
  assign io_in_dat_bits_mask_49 = _T_4018_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1726.4]
  assign io_in_dat_bits_mask_50 = _T_4018_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1727.4]
  assign io_in_dat_bits_mask_51 = _T_4018_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1728.4]
  assign io_in_dat_bits_mask_52 = _T_4018_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1729.4]
  assign io_in_dat_bits_mask_53 = _T_4018_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1730.4]
  assign io_in_dat_bits_mask_54 = _T_4018_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1731.4]
  assign io_in_dat_bits_mask_55 = _T_4018_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1732.4]
  assign io_in_dat_bits_mask_56 = _T_4018_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1733.4]
  assign io_in_dat_bits_mask_57 = _T_4018_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1734.4]
  assign io_in_dat_bits_mask_58 = _T_4018_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1735.4]
  assign io_in_dat_bits_mask_59 = _T_4018_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1736.4]
  assign io_in_dat_bits_mask_60 = _T_4018_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1737.4]
  assign io_in_dat_bits_mask_61 = _T_4018_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1738.4]
  assign io_in_dat_bits_mask_62 = _T_4018_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1739.4]
  assign io_in_dat_bits_mask_63 = _T_4018_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 104:25:@1740.4]
  assign io_in_dat_bits_data_0 = _T_3152_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1742.4]
  assign io_in_dat_bits_data_1 = _T_3152_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1743.4]
  assign io_in_dat_bits_data_2 = _T_3152_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1744.4]
  assign io_in_dat_bits_data_3 = _T_3152_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1745.4]
  assign io_in_dat_bits_data_4 = _T_3152_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1746.4]
  assign io_in_dat_bits_data_5 = _T_3152_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1747.4]
  assign io_in_dat_bits_data_6 = _T_3152_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1748.4]
  assign io_in_dat_bits_data_7 = _T_3152_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1749.4]
  assign io_in_dat_bits_data_8 = _T_3152_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1750.4]
  assign io_in_dat_bits_data_9 = _T_3152_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1751.4]
  assign io_in_dat_bits_data_10 = _T_3152_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1752.4]
  assign io_in_dat_bits_data_11 = _T_3152_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1753.4]
  assign io_in_dat_bits_data_12 = _T_3152_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1754.4]
  assign io_in_dat_bits_data_13 = _T_3152_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1755.4]
  assign io_in_dat_bits_data_14 = _T_3152_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1756.4]
  assign io_in_dat_bits_data_15 = _T_3152_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1757.4]
  assign io_in_dat_bits_data_16 = _T_3152_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1758.4]
  assign io_in_dat_bits_data_17 = _T_3152_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1759.4]
  assign io_in_dat_bits_data_18 = _T_3152_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1760.4]
  assign io_in_dat_bits_data_19 = _T_3152_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1761.4]
  assign io_in_dat_bits_data_20 = _T_3152_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1762.4]
  assign io_in_dat_bits_data_21 = _T_3152_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1763.4]
  assign io_in_dat_bits_data_22 = _T_3152_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1764.4]
  assign io_in_dat_bits_data_23 = _T_3152_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1765.4]
  assign io_in_dat_bits_data_24 = _T_3152_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1766.4]
  assign io_in_dat_bits_data_25 = _T_3152_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1767.4]
  assign io_in_dat_bits_data_26 = _T_3152_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1768.4]
  assign io_in_dat_bits_data_27 = _T_3152_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1769.4]
  assign io_in_dat_bits_data_28 = _T_3152_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1770.4]
  assign io_in_dat_bits_data_29 = _T_3152_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1771.4]
  assign io_in_dat_bits_data_30 = _T_3152_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1772.4]
  assign io_in_dat_bits_data_31 = _T_3152_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1773.4]
  assign io_in_dat_bits_data_32 = _T_3152_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1774.4]
  assign io_in_dat_bits_data_33 = _T_3152_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1775.4]
  assign io_in_dat_bits_data_34 = _T_3152_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1776.4]
  assign io_in_dat_bits_data_35 = _T_3152_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1777.4]
  assign io_in_dat_bits_data_36 = _T_3152_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1778.4]
  assign io_in_dat_bits_data_37 = _T_3152_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1779.4]
  assign io_in_dat_bits_data_38 = _T_3152_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1780.4]
  assign io_in_dat_bits_data_39 = _T_3152_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1781.4]
  assign io_in_dat_bits_data_40 = _T_3152_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1782.4]
  assign io_in_dat_bits_data_41 = _T_3152_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1783.4]
  assign io_in_dat_bits_data_42 = _T_3152_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1784.4]
  assign io_in_dat_bits_data_43 = _T_3152_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1785.4]
  assign io_in_dat_bits_data_44 = _T_3152_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1786.4]
  assign io_in_dat_bits_data_45 = _T_3152_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1787.4]
  assign io_in_dat_bits_data_46 = _T_3152_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1788.4]
  assign io_in_dat_bits_data_47 = _T_3152_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1789.4]
  assign io_in_dat_bits_data_48 = _T_3152_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1790.4]
  assign io_in_dat_bits_data_49 = _T_3152_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1791.4]
  assign io_in_dat_bits_data_50 = _T_3152_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1792.4]
  assign io_in_dat_bits_data_51 = _T_3152_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1793.4]
  assign io_in_dat_bits_data_52 = _T_3152_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1794.4]
  assign io_in_dat_bits_data_53 = _T_3152_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1795.4]
  assign io_in_dat_bits_data_54 = _T_3152_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1796.4]
  assign io_in_dat_bits_data_55 = _T_3152_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1797.4]
  assign io_in_dat_bits_data_56 = _T_3152_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1798.4]
  assign io_in_dat_bits_data_57 = _T_3152_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1799.4]
  assign io_in_dat_bits_data_58 = _T_3152_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1800.4]
  assign io_in_dat_bits_data_59 = _T_3152_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1801.4]
  assign io_in_dat_bits_data_60 = _T_3152_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1802.4]
  assign io_in_dat_bits_data_61 = _T_3152_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1803.4]
  assign io_in_dat_bits_data_62 = _T_3152_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1804.4]
  assign io_in_dat_bits_data_63 = _T_3152_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 106:25:@1805.4]
  assign io_in_dat_bits_pd = _T_4230; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 105:23:@1741.4]
  assign io_in_wt_valid = _T_5438; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 107:20:@1806.4]
  assign io_in_wt_bits_sel_0 = _T_5662_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 109:23:@1871.4]
  assign io_in_wt_bits_sel_1 = _T_5662_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 109:23:@1872.4]
  assign io_in_wt_bits_sel_2 = _T_5662_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 109:23:@1873.4]
  assign io_in_wt_bits_sel_3 = _T_5662_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 109:23:@1874.4]
  assign io_in_wt_bits_sel_4 = _T_5662_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 109:23:@1875.4]
  assign io_in_wt_bits_sel_5 = _T_5662_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 109:23:@1876.4]
  assign io_in_wt_bits_sel_6 = _T_5662_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 109:23:@1877.4]
  assign io_in_wt_bits_sel_7 = _T_5662_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 109:23:@1878.4]
  assign io_in_wt_bits_sel_8 = _T_5662_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 109:23:@1879.4]
  assign io_in_wt_bits_sel_9 = _T_5662_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 109:23:@1880.4]
  assign io_in_wt_bits_sel_10 = _T_5662_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 109:23:@1881.4]
  assign io_in_wt_bits_sel_11 = _T_5662_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 109:23:@1882.4]
  assign io_in_wt_bits_sel_12 = _T_5662_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 109:23:@1883.4]
  assign io_in_wt_bits_sel_13 = _T_5662_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 109:23:@1884.4]
  assign io_in_wt_bits_sel_14 = _T_5662_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 109:23:@1885.4]
  assign io_in_wt_bits_sel_15 = _T_5662_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 109:23:@1886.4]
  assign io_in_wt_bits_mask_0 = _T_5234_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1807.4]
  assign io_in_wt_bits_mask_1 = _T_5234_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1808.4]
  assign io_in_wt_bits_mask_2 = _T_5234_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1809.4]
  assign io_in_wt_bits_mask_3 = _T_5234_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1810.4]
  assign io_in_wt_bits_mask_4 = _T_5234_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1811.4]
  assign io_in_wt_bits_mask_5 = _T_5234_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1812.4]
  assign io_in_wt_bits_mask_6 = _T_5234_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1813.4]
  assign io_in_wt_bits_mask_7 = _T_5234_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1814.4]
  assign io_in_wt_bits_mask_8 = _T_5234_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1815.4]
  assign io_in_wt_bits_mask_9 = _T_5234_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1816.4]
  assign io_in_wt_bits_mask_10 = _T_5234_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1817.4]
  assign io_in_wt_bits_mask_11 = _T_5234_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1818.4]
  assign io_in_wt_bits_mask_12 = _T_5234_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1819.4]
  assign io_in_wt_bits_mask_13 = _T_5234_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1820.4]
  assign io_in_wt_bits_mask_14 = _T_5234_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1821.4]
  assign io_in_wt_bits_mask_15 = _T_5234_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1822.4]
  assign io_in_wt_bits_mask_16 = _T_5234_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1823.4]
  assign io_in_wt_bits_mask_17 = _T_5234_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1824.4]
  assign io_in_wt_bits_mask_18 = _T_5234_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1825.4]
  assign io_in_wt_bits_mask_19 = _T_5234_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1826.4]
  assign io_in_wt_bits_mask_20 = _T_5234_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1827.4]
  assign io_in_wt_bits_mask_21 = _T_5234_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1828.4]
  assign io_in_wt_bits_mask_22 = _T_5234_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1829.4]
  assign io_in_wt_bits_mask_23 = _T_5234_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1830.4]
  assign io_in_wt_bits_mask_24 = _T_5234_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1831.4]
  assign io_in_wt_bits_mask_25 = _T_5234_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1832.4]
  assign io_in_wt_bits_mask_26 = _T_5234_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1833.4]
  assign io_in_wt_bits_mask_27 = _T_5234_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1834.4]
  assign io_in_wt_bits_mask_28 = _T_5234_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1835.4]
  assign io_in_wt_bits_mask_29 = _T_5234_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1836.4]
  assign io_in_wt_bits_mask_30 = _T_5234_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1837.4]
  assign io_in_wt_bits_mask_31 = _T_5234_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1838.4]
  assign io_in_wt_bits_mask_32 = _T_5234_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1839.4]
  assign io_in_wt_bits_mask_33 = _T_5234_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1840.4]
  assign io_in_wt_bits_mask_34 = _T_5234_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1841.4]
  assign io_in_wt_bits_mask_35 = _T_5234_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1842.4]
  assign io_in_wt_bits_mask_36 = _T_5234_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1843.4]
  assign io_in_wt_bits_mask_37 = _T_5234_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1844.4]
  assign io_in_wt_bits_mask_38 = _T_5234_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1845.4]
  assign io_in_wt_bits_mask_39 = _T_5234_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1846.4]
  assign io_in_wt_bits_mask_40 = _T_5234_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1847.4]
  assign io_in_wt_bits_mask_41 = _T_5234_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1848.4]
  assign io_in_wt_bits_mask_42 = _T_5234_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1849.4]
  assign io_in_wt_bits_mask_43 = _T_5234_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1850.4]
  assign io_in_wt_bits_mask_44 = _T_5234_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1851.4]
  assign io_in_wt_bits_mask_45 = _T_5234_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1852.4]
  assign io_in_wt_bits_mask_46 = _T_5234_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1853.4]
  assign io_in_wt_bits_mask_47 = _T_5234_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1854.4]
  assign io_in_wt_bits_mask_48 = _T_5234_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1855.4]
  assign io_in_wt_bits_mask_49 = _T_5234_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1856.4]
  assign io_in_wt_bits_mask_50 = _T_5234_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1857.4]
  assign io_in_wt_bits_mask_51 = _T_5234_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1858.4]
  assign io_in_wt_bits_mask_52 = _T_5234_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1859.4]
  assign io_in_wt_bits_mask_53 = _T_5234_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1860.4]
  assign io_in_wt_bits_mask_54 = _T_5234_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1861.4]
  assign io_in_wt_bits_mask_55 = _T_5234_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1862.4]
  assign io_in_wt_bits_mask_56 = _T_5234_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1863.4]
  assign io_in_wt_bits_mask_57 = _T_5234_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1864.4]
  assign io_in_wt_bits_mask_58 = _T_5234_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1865.4]
  assign io_in_wt_bits_mask_59 = _T_5234_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1866.4]
  assign io_in_wt_bits_mask_60 = _T_5234_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1867.4]
  assign io_in_wt_bits_mask_61 = _T_5234_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1868.4]
  assign io_in_wt_bits_mask_62 = _T_5234_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1869.4]
  assign io_in_wt_bits_mask_63 = _T_5234_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 108:24:@1870.4]
  assign io_in_wt_bits_data_0 = _T_4368_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1887.4]
  assign io_in_wt_bits_data_1 = _T_4368_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1888.4]
  assign io_in_wt_bits_data_2 = _T_4368_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1889.4]
  assign io_in_wt_bits_data_3 = _T_4368_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1890.4]
  assign io_in_wt_bits_data_4 = _T_4368_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1891.4]
  assign io_in_wt_bits_data_5 = _T_4368_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1892.4]
  assign io_in_wt_bits_data_6 = _T_4368_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1893.4]
  assign io_in_wt_bits_data_7 = _T_4368_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1894.4]
  assign io_in_wt_bits_data_8 = _T_4368_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1895.4]
  assign io_in_wt_bits_data_9 = _T_4368_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1896.4]
  assign io_in_wt_bits_data_10 = _T_4368_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1897.4]
  assign io_in_wt_bits_data_11 = _T_4368_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1898.4]
  assign io_in_wt_bits_data_12 = _T_4368_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1899.4]
  assign io_in_wt_bits_data_13 = _T_4368_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1900.4]
  assign io_in_wt_bits_data_14 = _T_4368_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1901.4]
  assign io_in_wt_bits_data_15 = _T_4368_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1902.4]
  assign io_in_wt_bits_data_16 = _T_4368_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1903.4]
  assign io_in_wt_bits_data_17 = _T_4368_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1904.4]
  assign io_in_wt_bits_data_18 = _T_4368_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1905.4]
  assign io_in_wt_bits_data_19 = _T_4368_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1906.4]
  assign io_in_wt_bits_data_20 = _T_4368_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1907.4]
  assign io_in_wt_bits_data_21 = _T_4368_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1908.4]
  assign io_in_wt_bits_data_22 = _T_4368_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1909.4]
  assign io_in_wt_bits_data_23 = _T_4368_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1910.4]
  assign io_in_wt_bits_data_24 = _T_4368_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1911.4]
  assign io_in_wt_bits_data_25 = _T_4368_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1912.4]
  assign io_in_wt_bits_data_26 = _T_4368_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1913.4]
  assign io_in_wt_bits_data_27 = _T_4368_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1914.4]
  assign io_in_wt_bits_data_28 = _T_4368_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1915.4]
  assign io_in_wt_bits_data_29 = _T_4368_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1916.4]
  assign io_in_wt_bits_data_30 = _T_4368_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1917.4]
  assign io_in_wt_bits_data_31 = _T_4368_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1918.4]
  assign io_in_wt_bits_data_32 = _T_4368_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1919.4]
  assign io_in_wt_bits_data_33 = _T_4368_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1920.4]
  assign io_in_wt_bits_data_34 = _T_4368_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1921.4]
  assign io_in_wt_bits_data_35 = _T_4368_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1922.4]
  assign io_in_wt_bits_data_36 = _T_4368_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1923.4]
  assign io_in_wt_bits_data_37 = _T_4368_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1924.4]
  assign io_in_wt_bits_data_38 = _T_4368_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1925.4]
  assign io_in_wt_bits_data_39 = _T_4368_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1926.4]
  assign io_in_wt_bits_data_40 = _T_4368_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1927.4]
  assign io_in_wt_bits_data_41 = _T_4368_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1928.4]
  assign io_in_wt_bits_data_42 = _T_4368_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1929.4]
  assign io_in_wt_bits_data_43 = _T_4368_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1930.4]
  assign io_in_wt_bits_data_44 = _T_4368_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1931.4]
  assign io_in_wt_bits_data_45 = _T_4368_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1932.4]
  assign io_in_wt_bits_data_46 = _T_4368_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1933.4]
  assign io_in_wt_bits_data_47 = _T_4368_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1934.4]
  assign io_in_wt_bits_data_48 = _T_4368_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1935.4]
  assign io_in_wt_bits_data_49 = _T_4368_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1936.4]
  assign io_in_wt_bits_data_50 = _T_4368_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1937.4]
  assign io_in_wt_bits_data_51 = _T_4368_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1938.4]
  assign io_in_wt_bits_data_52 = _T_4368_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1939.4]
  assign io_in_wt_bits_data_53 = _T_4368_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1940.4]
  assign io_in_wt_bits_data_54 = _T_4368_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1941.4]
  assign io_in_wt_bits_data_55 = _T_4368_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1942.4]
  assign io_in_wt_bits_data_56 = _T_4368_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1943.4]
  assign io_in_wt_bits_data_57 = _T_4368_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1944.4]
  assign io_in_wt_bits_data_58 = _T_4368_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1945.4]
  assign io_in_wt_bits_data_59 = _T_4368_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1946.4]
  assign io_in_wt_bits_data_60 = _T_4368_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1947.4]
  assign io_in_wt_bits_data_61 = _T_4368_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1948.4]
  assign io_in_wt_bits_data_62 = _T_4368_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1949.4]
  assign io_in_wt_bits_data_63 = _T_4368_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 110:24:@1950.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_3085_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_3085_1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_3085_2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3085_3 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_3085_4 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_3085_5 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_3085_6 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_3085_7 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_3085_8 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_3085_9 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_3085_10 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_3085_11 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_3085_12 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_3085_13 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_3085_14 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_3085_15 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_3085_16 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_3085_17 = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_3085_18 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_3085_19 = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_3085_20 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_3085_21 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_3085_22 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_3085_23 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_3085_24 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_3085_25 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_3085_26 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_3085_27 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_3085_28 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_3085_29 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_3085_30 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_3085_31 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_3085_32 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_3085_33 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_3085_34 = _RAND_34[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_3085_35 = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_3085_36 = _RAND_36[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_3085_37 = _RAND_37[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_3085_38 = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_3085_39 = _RAND_39[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_3085_40 = _RAND_40[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_3085_41 = _RAND_41[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_3085_42 = _RAND_42[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_3085_43 = _RAND_43[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_3085_44 = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_3085_45 = _RAND_45[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_3085_46 = _RAND_46[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_3085_47 = _RAND_47[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_3085_48 = _RAND_48[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_3085_49 = _RAND_49[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_3085_50 = _RAND_50[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_3085_51 = _RAND_51[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_3085_52 = _RAND_52[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_3085_53 = _RAND_53[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_3085_54 = _RAND_54[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_3085_55 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_3085_56 = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_3085_57 = _RAND_57[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_3085_58 = _RAND_58[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_3085_59 = _RAND_59[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_3085_60 = _RAND_60[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_3085_61 = _RAND_61[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_3085_62 = _RAND_62[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_3085_63 = _RAND_63[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_3152_0 = _RAND_64[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_3152_1 = _RAND_65[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_3152_2 = _RAND_66[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_3152_3 = _RAND_67[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_3152_4 = _RAND_68[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_3152_5 = _RAND_69[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_3152_6 = _RAND_70[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_3152_7 = _RAND_71[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_3152_8 = _RAND_72[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_3152_9 = _RAND_73[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_3152_10 = _RAND_74[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_3152_11 = _RAND_75[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_3152_12 = _RAND_76[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_3152_13 = _RAND_77[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_3152_14 = _RAND_78[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_3152_15 = _RAND_79[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_3152_16 = _RAND_80[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_3152_17 = _RAND_81[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_3152_18 = _RAND_82[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_3152_19 = _RAND_83[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_3152_20 = _RAND_84[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_3152_21 = _RAND_85[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_3152_22 = _RAND_86[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_3152_23 = _RAND_87[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_3152_24 = _RAND_88[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_3152_25 = _RAND_89[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_3152_26 = _RAND_90[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_3152_27 = _RAND_91[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_3152_28 = _RAND_92[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_3152_29 = _RAND_93[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_3152_30 = _RAND_94[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_3152_31 = _RAND_95[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_3152_32 = _RAND_96[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_3152_33 = _RAND_97[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_3152_34 = _RAND_98[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_3152_35 = _RAND_99[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_3152_36 = _RAND_100[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_3152_37 = _RAND_101[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_3152_38 = _RAND_102[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_3152_39 = _RAND_103[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_3152_40 = _RAND_104[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_3152_41 = _RAND_105[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_3152_42 = _RAND_106[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_3152_43 = _RAND_107[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_3152_44 = _RAND_108[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_3152_45 = _RAND_109[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_3152_46 = _RAND_110[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_3152_47 = _RAND_111[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_3152_48 = _RAND_112[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_3152_49 = _RAND_113[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_3152_50 = _RAND_114[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_3152_51 = _RAND_115[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_3152_52 = _RAND_116[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_3152_53 = _RAND_117[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_3152_54 = _RAND_118[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_3152_55 = _RAND_119[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_3152_56 = _RAND_120[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_3152_57 = _RAND_121[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_3152_58 = _RAND_122[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_3152_59 = _RAND_123[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_3152_60 = _RAND_124[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_3152_61 = _RAND_125[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_3152_62 = _RAND_126[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_3152_63 = _RAND_127[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_3555_0 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_3555_1 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_3555_2 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_3555_3 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_3555_4 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_3555_5 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_3555_6 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_3555_7 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_3555_8 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_3555_9 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_3555_10 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_3555_11 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_3555_12 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_3555_13 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_3555_14 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_3555_15 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_3555_16 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_3555_17 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_3555_18 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_3555_19 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_3555_20 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_3555_21 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_3555_22 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_3555_23 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_3555_24 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_3555_25 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_3555_26 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_3555_27 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_3555_28 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_3555_29 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_3555_30 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_3555_31 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_3555_32 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_3555_33 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_3555_34 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_3555_35 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_3555_36 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_3555_37 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_3555_38 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_3555_39 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_3555_40 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_3555_41 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_3555_42 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_3555_43 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_3555_44 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_3555_45 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_3555_46 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_3555_47 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_3555_48 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_3555_49 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_3555_50 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_3555_51 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_3555_52 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_3555_53 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_3555_54 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_3555_55 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_3555_56 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_3555_57 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_3555_58 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_3555_59 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_3555_60 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_3555_61 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_3555_62 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_3555_63 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_4018_0 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_4018_1 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_4018_2 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_4018_3 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_4018_4 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_4018_5 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_4018_6 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_4018_7 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_4018_8 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_4018_9 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_4018_10 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_4018_11 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_4018_12 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_4018_13 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_4018_14 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_4018_15 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_4018_16 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_4018_17 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_4018_18 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_4018_19 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_4018_20 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_4018_21 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_4018_22 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_4018_23 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_4018_24 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_4018_25 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_4018_26 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_4018_27 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_4018_28 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_4018_29 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_4018_30 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_4018_31 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_4018_32 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_4018_33 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_4018_34 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_4018_35 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_4018_36 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_4018_37 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_4018_38 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_4018_39 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_4018_40 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_4018_41 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_4018_42 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_4018_43 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_4018_44 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_4018_45 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_4018_46 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_4018_47 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_4018_48 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_4018_49 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_4018_50 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_4018_51 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_4018_52 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_4018_53 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_4018_54 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_4018_55 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_4018_56 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_4018_57 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_4018_58 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_4018_59 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_4018_60 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_4018_61 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_4018_62 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_4018_63 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_4219 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_4222 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_4227 = _RAND_258[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_4230 = _RAND_259[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_4301_0 = _RAND_260[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_4301_1 = _RAND_261[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_4301_2 = _RAND_262[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_4301_3 = _RAND_263[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_4301_4 = _RAND_264[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_4301_5 = _RAND_265[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_4301_6 = _RAND_266[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_4301_7 = _RAND_267[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_4301_8 = _RAND_268[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_4301_9 = _RAND_269[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_4301_10 = _RAND_270[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_4301_11 = _RAND_271[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_4301_12 = _RAND_272[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_4301_13 = _RAND_273[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_4301_14 = _RAND_274[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_4301_15 = _RAND_275[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_4301_16 = _RAND_276[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_4301_17 = _RAND_277[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_4301_18 = _RAND_278[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_4301_19 = _RAND_279[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_4301_20 = _RAND_280[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_4301_21 = _RAND_281[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_4301_22 = _RAND_282[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_4301_23 = _RAND_283[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_4301_24 = _RAND_284[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_4301_25 = _RAND_285[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_4301_26 = _RAND_286[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_4301_27 = _RAND_287[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_4301_28 = _RAND_288[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_4301_29 = _RAND_289[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_4301_30 = _RAND_290[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_4301_31 = _RAND_291[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_4301_32 = _RAND_292[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_4301_33 = _RAND_293[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_4301_34 = _RAND_294[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_4301_35 = _RAND_295[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_4301_36 = _RAND_296[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_4301_37 = _RAND_297[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_4301_38 = _RAND_298[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_4301_39 = _RAND_299[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_4301_40 = _RAND_300[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_4301_41 = _RAND_301[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_4301_42 = _RAND_302[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_4301_43 = _RAND_303[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_4301_44 = _RAND_304[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_4301_45 = _RAND_305[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_4301_46 = _RAND_306[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_4301_47 = _RAND_307[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_4301_48 = _RAND_308[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_4301_49 = _RAND_309[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_4301_50 = _RAND_310[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_4301_51 = _RAND_311[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_4301_52 = _RAND_312[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_4301_53 = _RAND_313[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_4301_54 = _RAND_314[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_4301_55 = _RAND_315[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_4301_56 = _RAND_316[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_4301_57 = _RAND_317[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_4301_58 = _RAND_318[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_4301_59 = _RAND_319[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_4301_60 = _RAND_320[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_4301_61 = _RAND_321[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_4301_62 = _RAND_322[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_4301_63 = _RAND_323[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_4368_0 = _RAND_324[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_4368_1 = _RAND_325[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_4368_2 = _RAND_326[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_4368_3 = _RAND_327[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_4368_4 = _RAND_328[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_4368_5 = _RAND_329[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_4368_6 = _RAND_330[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_4368_7 = _RAND_331[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_4368_8 = _RAND_332[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_4368_9 = _RAND_333[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_4368_10 = _RAND_334[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_4368_11 = _RAND_335[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_4368_12 = _RAND_336[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_4368_13 = _RAND_337[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_4368_14 = _RAND_338[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_4368_15 = _RAND_339[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_4368_16 = _RAND_340[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_4368_17 = _RAND_341[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_4368_18 = _RAND_342[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_4368_19 = _RAND_343[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_4368_20 = _RAND_344[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_4368_21 = _RAND_345[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_4368_22 = _RAND_346[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_4368_23 = _RAND_347[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_4368_24 = _RAND_348[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_4368_25 = _RAND_349[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_4368_26 = _RAND_350[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_4368_27 = _RAND_351[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_4368_28 = _RAND_352[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_4368_29 = _RAND_353[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_4368_30 = _RAND_354[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_4368_31 = _RAND_355[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_4368_32 = _RAND_356[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_4368_33 = _RAND_357[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_4368_34 = _RAND_358[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_4368_35 = _RAND_359[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_4368_36 = _RAND_360[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_4368_37 = _RAND_361[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_4368_38 = _RAND_362[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_4368_39 = _RAND_363[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_4368_40 = _RAND_364[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_4368_41 = _RAND_365[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_4368_42 = _RAND_366[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_4368_43 = _RAND_367[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_4368_44 = _RAND_368[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_4368_45 = _RAND_369[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_4368_46 = _RAND_370[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_4368_47 = _RAND_371[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_4368_48 = _RAND_372[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_4368_49 = _RAND_373[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_4368_50 = _RAND_374[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_4368_51 = _RAND_375[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_4368_52 = _RAND_376[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_4368_53 = _RAND_377[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_4368_54 = _RAND_378[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_4368_55 = _RAND_379[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_4368_56 = _RAND_380[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_4368_57 = _RAND_381[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_4368_58 = _RAND_382[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_4368_59 = _RAND_383[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_4368_60 = _RAND_384[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_4368_61 = _RAND_385[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_4368_62 = _RAND_386[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_4368_63 = _RAND_387[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_4771_0 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_4771_1 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_4771_2 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_4771_3 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_4771_4 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_4771_5 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_4771_6 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_4771_7 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_4771_8 = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_4771_9 = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_4771_10 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_4771_11 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_4771_12 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_4771_13 = _RAND_401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_4771_14 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_4771_15 = _RAND_403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_4771_16 = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_4771_17 = _RAND_405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_4771_18 = _RAND_406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_4771_19 = _RAND_407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_4771_20 = _RAND_408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_4771_21 = _RAND_409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_4771_22 = _RAND_410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_4771_23 = _RAND_411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_4771_24 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_4771_25 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_4771_26 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_4771_27 = _RAND_415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_4771_28 = _RAND_416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_4771_29 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_4771_30 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_4771_31 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_4771_32 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_4771_33 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_4771_34 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_4771_35 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_4771_36 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_4771_37 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_4771_38 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_4771_39 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_4771_40 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_4771_41 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_4771_42 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_4771_43 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_4771_44 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_4771_45 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_4771_46 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_4771_47 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_4771_48 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_4771_49 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_4771_50 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_4771_51 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_4771_52 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_4771_53 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_4771_54 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_4771_55 = _RAND_443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_4771_56 = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_4771_57 = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_4771_58 = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_4771_59 = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_4771_60 = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_4771_61 = _RAND_449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_4771_62 = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_4771_63 = _RAND_451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_5234_0 = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_5234_1 = _RAND_453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_5234_2 = _RAND_454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_5234_3 = _RAND_455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_5234_4 = _RAND_456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_5234_5 = _RAND_457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_5234_6 = _RAND_458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_5234_7 = _RAND_459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_5234_8 = _RAND_460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_5234_9 = _RAND_461[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_5234_10 = _RAND_462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_5234_11 = _RAND_463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_5234_12 = _RAND_464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_5234_13 = _RAND_465[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_5234_14 = _RAND_466[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_5234_15 = _RAND_467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_5234_16 = _RAND_468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_5234_17 = _RAND_469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_5234_18 = _RAND_470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_5234_19 = _RAND_471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_5234_20 = _RAND_472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_5234_21 = _RAND_473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_5234_22 = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_5234_23 = _RAND_475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_5234_24 = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_5234_25 = _RAND_477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_5234_26 = _RAND_478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_5234_27 = _RAND_479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_5234_28 = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_5234_29 = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_5234_30 = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_5234_31 = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_5234_32 = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_5234_33 = _RAND_485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_5234_34 = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_5234_35 = _RAND_487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_5234_36 = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_5234_37 = _RAND_489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_5234_38 = _RAND_490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_5234_39 = _RAND_491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_5234_40 = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_5234_41 = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_5234_42 = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_5234_43 = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_5234_44 = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_5234_45 = _RAND_497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_5234_46 = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_5234_47 = _RAND_499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_5234_48 = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_5234_49 = _RAND_501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_5234_50 = _RAND_502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_5234_51 = _RAND_503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_5234_52 = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_5234_53 = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_5234_54 = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_5234_55 = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_5234_56 = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_5234_57 = _RAND_509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_5234_58 = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_5234_59 = _RAND_511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_5234_60 = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_5234_61 = _RAND_513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_5234_62 = _RAND_514[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_5234_63 = _RAND_515[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_5435 = _RAND_516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_5438 = _RAND_517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_5535_0 = _RAND_518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  _T_5535_1 = _RAND_519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  _T_5535_2 = _RAND_520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  _T_5535_3 = _RAND_521[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  _T_5535_4 = _RAND_522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  _T_5535_5 = _RAND_523[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  _T_5535_6 = _RAND_524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  _T_5535_7 = _RAND_525[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  _T_5535_8 = _RAND_526[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  _T_5535_9 = _RAND_527[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  _T_5535_10 = _RAND_528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  _T_5535_11 = _RAND_529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  _T_5535_12 = _RAND_530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  _T_5535_13 = _RAND_531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  _T_5535_14 = _RAND_532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  _T_5535_15 = _RAND_533[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  _T_5662_0 = _RAND_534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  _T_5662_1 = _RAND_535[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  _T_5662_2 = _RAND_536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  _T_5662_3 = _RAND_537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  _T_5662_4 = _RAND_538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  _T_5662_5 = _RAND_539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  _T_5662_6 = _RAND_540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  _T_5662_7 = _RAND_541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  _T_5662_8 = _RAND_542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  _T_5662_9 = _RAND_543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  _T_5662_10 = _RAND_544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  _T_5662_11 = _RAND_545[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  _T_5662_12 = _RAND_546[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  _T_5662_13 = _RAND_547[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  _T_5662_14 = _RAND_548[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  _T_5662_15 = _RAND_549[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (io_sc2mac_dat_bits_mask_0) begin
      _T_3085_0 <= io_sc2mac_dat_bits_data_0;
    end
    if (io_sc2mac_dat_bits_mask_1) begin
      _T_3085_1 <= io_sc2mac_dat_bits_data_1;
    end
    if (io_sc2mac_dat_bits_mask_2) begin
      _T_3085_2 <= io_sc2mac_dat_bits_data_2;
    end
    if (io_sc2mac_dat_bits_mask_3) begin
      _T_3085_3 <= io_sc2mac_dat_bits_data_3;
    end
    if (io_sc2mac_dat_bits_mask_4) begin
      _T_3085_4 <= io_sc2mac_dat_bits_data_4;
    end
    if (io_sc2mac_dat_bits_mask_5) begin
      _T_3085_5 <= io_sc2mac_dat_bits_data_5;
    end
    if (io_sc2mac_dat_bits_mask_6) begin
      _T_3085_6 <= io_sc2mac_dat_bits_data_6;
    end
    if (io_sc2mac_dat_bits_mask_7) begin
      _T_3085_7 <= io_sc2mac_dat_bits_data_7;
    end
    if (io_sc2mac_dat_bits_mask_8) begin
      _T_3085_8 <= io_sc2mac_dat_bits_data_8;
    end
    if (io_sc2mac_dat_bits_mask_9) begin
      _T_3085_9 <= io_sc2mac_dat_bits_data_9;
    end
    if (io_sc2mac_dat_bits_mask_10) begin
      _T_3085_10 <= io_sc2mac_dat_bits_data_10;
    end
    if (io_sc2mac_dat_bits_mask_11) begin
      _T_3085_11 <= io_sc2mac_dat_bits_data_11;
    end
    if (io_sc2mac_dat_bits_mask_12) begin
      _T_3085_12 <= io_sc2mac_dat_bits_data_12;
    end
    if (io_sc2mac_dat_bits_mask_13) begin
      _T_3085_13 <= io_sc2mac_dat_bits_data_13;
    end
    if (io_sc2mac_dat_bits_mask_14) begin
      _T_3085_14 <= io_sc2mac_dat_bits_data_14;
    end
    if (io_sc2mac_dat_bits_mask_15) begin
      _T_3085_15 <= io_sc2mac_dat_bits_data_15;
    end
    if (io_sc2mac_dat_bits_mask_16) begin
      _T_3085_16 <= io_sc2mac_dat_bits_data_16;
    end
    if (io_sc2mac_dat_bits_mask_17) begin
      _T_3085_17 <= io_sc2mac_dat_bits_data_17;
    end
    if (io_sc2mac_dat_bits_mask_18) begin
      _T_3085_18 <= io_sc2mac_dat_bits_data_18;
    end
    if (io_sc2mac_dat_bits_mask_19) begin
      _T_3085_19 <= io_sc2mac_dat_bits_data_19;
    end
    if (io_sc2mac_dat_bits_mask_20) begin
      _T_3085_20 <= io_sc2mac_dat_bits_data_20;
    end
    if (io_sc2mac_dat_bits_mask_21) begin
      _T_3085_21 <= io_sc2mac_dat_bits_data_21;
    end
    if (io_sc2mac_dat_bits_mask_22) begin
      _T_3085_22 <= io_sc2mac_dat_bits_data_22;
    end
    if (io_sc2mac_dat_bits_mask_23) begin
      _T_3085_23 <= io_sc2mac_dat_bits_data_23;
    end
    if (io_sc2mac_dat_bits_mask_24) begin
      _T_3085_24 <= io_sc2mac_dat_bits_data_24;
    end
    if (io_sc2mac_dat_bits_mask_25) begin
      _T_3085_25 <= io_sc2mac_dat_bits_data_25;
    end
    if (io_sc2mac_dat_bits_mask_26) begin
      _T_3085_26 <= io_sc2mac_dat_bits_data_26;
    end
    if (io_sc2mac_dat_bits_mask_27) begin
      _T_3085_27 <= io_sc2mac_dat_bits_data_27;
    end
    if (io_sc2mac_dat_bits_mask_28) begin
      _T_3085_28 <= io_sc2mac_dat_bits_data_28;
    end
    if (io_sc2mac_dat_bits_mask_29) begin
      _T_3085_29 <= io_sc2mac_dat_bits_data_29;
    end
    if (io_sc2mac_dat_bits_mask_30) begin
      _T_3085_30 <= io_sc2mac_dat_bits_data_30;
    end
    if (io_sc2mac_dat_bits_mask_31) begin
      _T_3085_31 <= io_sc2mac_dat_bits_data_31;
    end
    if (io_sc2mac_dat_bits_mask_32) begin
      _T_3085_32 <= io_sc2mac_dat_bits_data_32;
    end
    if (io_sc2mac_dat_bits_mask_33) begin
      _T_3085_33 <= io_sc2mac_dat_bits_data_33;
    end
    if (io_sc2mac_dat_bits_mask_34) begin
      _T_3085_34 <= io_sc2mac_dat_bits_data_34;
    end
    if (io_sc2mac_dat_bits_mask_35) begin
      _T_3085_35 <= io_sc2mac_dat_bits_data_35;
    end
    if (io_sc2mac_dat_bits_mask_36) begin
      _T_3085_36 <= io_sc2mac_dat_bits_data_36;
    end
    if (io_sc2mac_dat_bits_mask_37) begin
      _T_3085_37 <= io_sc2mac_dat_bits_data_37;
    end
    if (io_sc2mac_dat_bits_mask_38) begin
      _T_3085_38 <= io_sc2mac_dat_bits_data_38;
    end
    if (io_sc2mac_dat_bits_mask_39) begin
      _T_3085_39 <= io_sc2mac_dat_bits_data_39;
    end
    if (io_sc2mac_dat_bits_mask_40) begin
      _T_3085_40 <= io_sc2mac_dat_bits_data_40;
    end
    if (io_sc2mac_dat_bits_mask_41) begin
      _T_3085_41 <= io_sc2mac_dat_bits_data_41;
    end
    if (io_sc2mac_dat_bits_mask_42) begin
      _T_3085_42 <= io_sc2mac_dat_bits_data_42;
    end
    if (io_sc2mac_dat_bits_mask_43) begin
      _T_3085_43 <= io_sc2mac_dat_bits_data_43;
    end
    if (io_sc2mac_dat_bits_mask_44) begin
      _T_3085_44 <= io_sc2mac_dat_bits_data_44;
    end
    if (io_sc2mac_dat_bits_mask_45) begin
      _T_3085_45 <= io_sc2mac_dat_bits_data_45;
    end
    if (io_sc2mac_dat_bits_mask_46) begin
      _T_3085_46 <= io_sc2mac_dat_bits_data_46;
    end
    if (io_sc2mac_dat_bits_mask_47) begin
      _T_3085_47 <= io_sc2mac_dat_bits_data_47;
    end
    if (io_sc2mac_dat_bits_mask_48) begin
      _T_3085_48 <= io_sc2mac_dat_bits_data_48;
    end
    if (io_sc2mac_dat_bits_mask_49) begin
      _T_3085_49 <= io_sc2mac_dat_bits_data_49;
    end
    if (io_sc2mac_dat_bits_mask_50) begin
      _T_3085_50 <= io_sc2mac_dat_bits_data_50;
    end
    if (io_sc2mac_dat_bits_mask_51) begin
      _T_3085_51 <= io_sc2mac_dat_bits_data_51;
    end
    if (io_sc2mac_dat_bits_mask_52) begin
      _T_3085_52 <= io_sc2mac_dat_bits_data_52;
    end
    if (io_sc2mac_dat_bits_mask_53) begin
      _T_3085_53 <= io_sc2mac_dat_bits_data_53;
    end
    if (io_sc2mac_dat_bits_mask_54) begin
      _T_3085_54 <= io_sc2mac_dat_bits_data_54;
    end
    if (io_sc2mac_dat_bits_mask_55) begin
      _T_3085_55 <= io_sc2mac_dat_bits_data_55;
    end
    if (io_sc2mac_dat_bits_mask_56) begin
      _T_3085_56 <= io_sc2mac_dat_bits_data_56;
    end
    if (io_sc2mac_dat_bits_mask_57) begin
      _T_3085_57 <= io_sc2mac_dat_bits_data_57;
    end
    if (io_sc2mac_dat_bits_mask_58) begin
      _T_3085_58 <= io_sc2mac_dat_bits_data_58;
    end
    if (io_sc2mac_dat_bits_mask_59) begin
      _T_3085_59 <= io_sc2mac_dat_bits_data_59;
    end
    if (io_sc2mac_dat_bits_mask_60) begin
      _T_3085_60 <= io_sc2mac_dat_bits_data_60;
    end
    if (io_sc2mac_dat_bits_mask_61) begin
      _T_3085_61 <= io_sc2mac_dat_bits_data_61;
    end
    if (io_sc2mac_dat_bits_mask_62) begin
      _T_3085_62 <= io_sc2mac_dat_bits_data_62;
    end
    if (io_sc2mac_dat_bits_mask_63) begin
      _T_3085_63 <= io_sc2mac_dat_bits_data_63;
    end
    if (_T_3555_0) begin
      _T_3152_0 <= _T_3085_0;
    end
    if (_T_3555_1) begin
      _T_3152_1 <= _T_3085_1;
    end
    if (_T_3555_2) begin
      _T_3152_2 <= _T_3085_2;
    end
    if (_T_3555_3) begin
      _T_3152_3 <= _T_3085_3;
    end
    if (_T_3555_4) begin
      _T_3152_4 <= _T_3085_4;
    end
    if (_T_3555_5) begin
      _T_3152_5 <= _T_3085_5;
    end
    if (_T_3555_6) begin
      _T_3152_6 <= _T_3085_6;
    end
    if (_T_3555_7) begin
      _T_3152_7 <= _T_3085_7;
    end
    if (_T_3555_8) begin
      _T_3152_8 <= _T_3085_8;
    end
    if (_T_3555_9) begin
      _T_3152_9 <= _T_3085_9;
    end
    if (_T_3555_10) begin
      _T_3152_10 <= _T_3085_10;
    end
    if (_T_3555_11) begin
      _T_3152_11 <= _T_3085_11;
    end
    if (_T_3555_12) begin
      _T_3152_12 <= _T_3085_12;
    end
    if (_T_3555_13) begin
      _T_3152_13 <= _T_3085_13;
    end
    if (_T_3555_14) begin
      _T_3152_14 <= _T_3085_14;
    end
    if (_T_3555_15) begin
      _T_3152_15 <= _T_3085_15;
    end
    if (_T_3555_16) begin
      _T_3152_16 <= _T_3085_16;
    end
    if (_T_3555_17) begin
      _T_3152_17 <= _T_3085_17;
    end
    if (_T_3555_18) begin
      _T_3152_18 <= _T_3085_18;
    end
    if (_T_3555_19) begin
      _T_3152_19 <= _T_3085_19;
    end
    if (_T_3555_20) begin
      _T_3152_20 <= _T_3085_20;
    end
    if (_T_3555_21) begin
      _T_3152_21 <= _T_3085_21;
    end
    if (_T_3555_22) begin
      _T_3152_22 <= _T_3085_22;
    end
    if (_T_3555_23) begin
      _T_3152_23 <= _T_3085_23;
    end
    if (_T_3555_24) begin
      _T_3152_24 <= _T_3085_24;
    end
    if (_T_3555_25) begin
      _T_3152_25 <= _T_3085_25;
    end
    if (_T_3555_26) begin
      _T_3152_26 <= _T_3085_26;
    end
    if (_T_3555_27) begin
      _T_3152_27 <= _T_3085_27;
    end
    if (_T_3555_28) begin
      _T_3152_28 <= _T_3085_28;
    end
    if (_T_3555_29) begin
      _T_3152_29 <= _T_3085_29;
    end
    if (_T_3555_30) begin
      _T_3152_30 <= _T_3085_30;
    end
    if (_T_3555_31) begin
      _T_3152_31 <= _T_3085_31;
    end
    if (_T_3555_32) begin
      _T_3152_32 <= _T_3085_32;
    end
    if (_T_3555_33) begin
      _T_3152_33 <= _T_3085_33;
    end
    if (_T_3555_34) begin
      _T_3152_34 <= _T_3085_34;
    end
    if (_T_3555_35) begin
      _T_3152_35 <= _T_3085_35;
    end
    if (_T_3555_36) begin
      _T_3152_36 <= _T_3085_36;
    end
    if (_T_3555_37) begin
      _T_3152_37 <= _T_3085_37;
    end
    if (_T_3555_38) begin
      _T_3152_38 <= _T_3085_38;
    end
    if (_T_3555_39) begin
      _T_3152_39 <= _T_3085_39;
    end
    if (_T_3555_40) begin
      _T_3152_40 <= _T_3085_40;
    end
    if (_T_3555_41) begin
      _T_3152_41 <= _T_3085_41;
    end
    if (_T_3555_42) begin
      _T_3152_42 <= _T_3085_42;
    end
    if (_T_3555_43) begin
      _T_3152_43 <= _T_3085_43;
    end
    if (_T_3555_44) begin
      _T_3152_44 <= _T_3085_44;
    end
    if (_T_3555_45) begin
      _T_3152_45 <= _T_3085_45;
    end
    if (_T_3555_46) begin
      _T_3152_46 <= _T_3085_46;
    end
    if (_T_3555_47) begin
      _T_3152_47 <= _T_3085_47;
    end
    if (_T_3555_48) begin
      _T_3152_48 <= _T_3085_48;
    end
    if (_T_3555_49) begin
      _T_3152_49 <= _T_3085_49;
    end
    if (_T_3555_50) begin
      _T_3152_50 <= _T_3085_50;
    end
    if (_T_3555_51) begin
      _T_3152_51 <= _T_3085_51;
    end
    if (_T_3555_52) begin
      _T_3152_52 <= _T_3085_52;
    end
    if (_T_3555_53) begin
      _T_3152_53 <= _T_3085_53;
    end
    if (_T_3555_54) begin
      _T_3152_54 <= _T_3085_54;
    end
    if (_T_3555_55) begin
      _T_3152_55 <= _T_3085_55;
    end
    if (_T_3555_56) begin
      _T_3152_56 <= _T_3085_56;
    end
    if (_T_3555_57) begin
      _T_3152_57 <= _T_3085_57;
    end
    if (_T_3555_58) begin
      _T_3152_58 <= _T_3085_58;
    end
    if (_T_3555_59) begin
      _T_3152_59 <= _T_3085_59;
    end
    if (_T_3555_60) begin
      _T_3152_60 <= _T_3085_60;
    end
    if (_T_3555_61) begin
      _T_3152_61 <= _T_3085_61;
    end
    if (_T_3555_62) begin
      _T_3152_62 <= _T_3085_62;
    end
    if (_T_3555_63) begin
      _T_3152_63 <= _T_3085_63;
    end
    if (_T_3014) begin
      _T_3555_0 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_0 <= io_sc2mac_dat_bits_mask_0;
      end
    end
    if (_T_3014) begin
      _T_3555_1 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_1 <= io_sc2mac_dat_bits_mask_1;
      end
    end
    if (_T_3014) begin
      _T_3555_2 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_2 <= io_sc2mac_dat_bits_mask_2;
      end
    end
    if (_T_3014) begin
      _T_3555_3 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_3 <= io_sc2mac_dat_bits_mask_3;
      end
    end
    if (_T_3014) begin
      _T_3555_4 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_4 <= io_sc2mac_dat_bits_mask_4;
      end
    end
    if (_T_3014) begin
      _T_3555_5 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_5 <= io_sc2mac_dat_bits_mask_5;
      end
    end
    if (_T_3014) begin
      _T_3555_6 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_6 <= io_sc2mac_dat_bits_mask_6;
      end
    end
    if (_T_3014) begin
      _T_3555_7 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_7 <= io_sc2mac_dat_bits_mask_7;
      end
    end
    if (_T_3014) begin
      _T_3555_8 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_8 <= io_sc2mac_dat_bits_mask_8;
      end
    end
    if (_T_3014) begin
      _T_3555_9 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_9 <= io_sc2mac_dat_bits_mask_9;
      end
    end
    if (_T_3014) begin
      _T_3555_10 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_10 <= io_sc2mac_dat_bits_mask_10;
      end
    end
    if (_T_3014) begin
      _T_3555_11 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_11 <= io_sc2mac_dat_bits_mask_11;
      end
    end
    if (_T_3014) begin
      _T_3555_12 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_12 <= io_sc2mac_dat_bits_mask_12;
      end
    end
    if (_T_3014) begin
      _T_3555_13 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_13 <= io_sc2mac_dat_bits_mask_13;
      end
    end
    if (_T_3014) begin
      _T_3555_14 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_14 <= io_sc2mac_dat_bits_mask_14;
      end
    end
    if (_T_3014) begin
      _T_3555_15 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_15 <= io_sc2mac_dat_bits_mask_15;
      end
    end
    if (_T_3014) begin
      _T_3555_16 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_16 <= io_sc2mac_dat_bits_mask_16;
      end
    end
    if (_T_3014) begin
      _T_3555_17 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_17 <= io_sc2mac_dat_bits_mask_17;
      end
    end
    if (_T_3014) begin
      _T_3555_18 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_18 <= io_sc2mac_dat_bits_mask_18;
      end
    end
    if (_T_3014) begin
      _T_3555_19 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_19 <= io_sc2mac_dat_bits_mask_19;
      end
    end
    if (_T_3014) begin
      _T_3555_20 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_20 <= io_sc2mac_dat_bits_mask_20;
      end
    end
    if (_T_3014) begin
      _T_3555_21 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_21 <= io_sc2mac_dat_bits_mask_21;
      end
    end
    if (_T_3014) begin
      _T_3555_22 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_22 <= io_sc2mac_dat_bits_mask_22;
      end
    end
    if (_T_3014) begin
      _T_3555_23 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_23 <= io_sc2mac_dat_bits_mask_23;
      end
    end
    if (_T_3014) begin
      _T_3555_24 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_24 <= io_sc2mac_dat_bits_mask_24;
      end
    end
    if (_T_3014) begin
      _T_3555_25 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_25 <= io_sc2mac_dat_bits_mask_25;
      end
    end
    if (_T_3014) begin
      _T_3555_26 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_26 <= io_sc2mac_dat_bits_mask_26;
      end
    end
    if (_T_3014) begin
      _T_3555_27 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_27 <= io_sc2mac_dat_bits_mask_27;
      end
    end
    if (_T_3014) begin
      _T_3555_28 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_28 <= io_sc2mac_dat_bits_mask_28;
      end
    end
    if (_T_3014) begin
      _T_3555_29 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_29 <= io_sc2mac_dat_bits_mask_29;
      end
    end
    if (_T_3014) begin
      _T_3555_30 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_30 <= io_sc2mac_dat_bits_mask_30;
      end
    end
    if (_T_3014) begin
      _T_3555_31 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_31 <= io_sc2mac_dat_bits_mask_31;
      end
    end
    if (_T_3014) begin
      _T_3555_32 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_32 <= io_sc2mac_dat_bits_mask_32;
      end
    end
    if (_T_3014) begin
      _T_3555_33 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_33 <= io_sc2mac_dat_bits_mask_33;
      end
    end
    if (_T_3014) begin
      _T_3555_34 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_34 <= io_sc2mac_dat_bits_mask_34;
      end
    end
    if (_T_3014) begin
      _T_3555_35 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_35 <= io_sc2mac_dat_bits_mask_35;
      end
    end
    if (_T_3014) begin
      _T_3555_36 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_36 <= io_sc2mac_dat_bits_mask_36;
      end
    end
    if (_T_3014) begin
      _T_3555_37 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_37 <= io_sc2mac_dat_bits_mask_37;
      end
    end
    if (_T_3014) begin
      _T_3555_38 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_38 <= io_sc2mac_dat_bits_mask_38;
      end
    end
    if (_T_3014) begin
      _T_3555_39 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_39 <= io_sc2mac_dat_bits_mask_39;
      end
    end
    if (_T_3014) begin
      _T_3555_40 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_40 <= io_sc2mac_dat_bits_mask_40;
      end
    end
    if (_T_3014) begin
      _T_3555_41 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_41 <= io_sc2mac_dat_bits_mask_41;
      end
    end
    if (_T_3014) begin
      _T_3555_42 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_42 <= io_sc2mac_dat_bits_mask_42;
      end
    end
    if (_T_3014) begin
      _T_3555_43 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_43 <= io_sc2mac_dat_bits_mask_43;
      end
    end
    if (_T_3014) begin
      _T_3555_44 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_44 <= io_sc2mac_dat_bits_mask_44;
      end
    end
    if (_T_3014) begin
      _T_3555_45 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_45 <= io_sc2mac_dat_bits_mask_45;
      end
    end
    if (_T_3014) begin
      _T_3555_46 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_46 <= io_sc2mac_dat_bits_mask_46;
      end
    end
    if (_T_3014) begin
      _T_3555_47 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_47 <= io_sc2mac_dat_bits_mask_47;
      end
    end
    if (_T_3014) begin
      _T_3555_48 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_48 <= io_sc2mac_dat_bits_mask_48;
      end
    end
    if (_T_3014) begin
      _T_3555_49 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_49 <= io_sc2mac_dat_bits_mask_49;
      end
    end
    if (_T_3014) begin
      _T_3555_50 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_50 <= io_sc2mac_dat_bits_mask_50;
      end
    end
    if (_T_3014) begin
      _T_3555_51 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_51 <= io_sc2mac_dat_bits_mask_51;
      end
    end
    if (_T_3014) begin
      _T_3555_52 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_52 <= io_sc2mac_dat_bits_mask_52;
      end
    end
    if (_T_3014) begin
      _T_3555_53 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_53 <= io_sc2mac_dat_bits_mask_53;
      end
    end
    if (_T_3014) begin
      _T_3555_54 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_54 <= io_sc2mac_dat_bits_mask_54;
      end
    end
    if (_T_3014) begin
      _T_3555_55 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_55 <= io_sc2mac_dat_bits_mask_55;
      end
    end
    if (_T_3014) begin
      _T_3555_56 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_56 <= io_sc2mac_dat_bits_mask_56;
      end
    end
    if (_T_3014) begin
      _T_3555_57 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_57 <= io_sc2mac_dat_bits_mask_57;
      end
    end
    if (_T_3014) begin
      _T_3555_58 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_58 <= io_sc2mac_dat_bits_mask_58;
      end
    end
    if (_T_3014) begin
      _T_3555_59 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_59 <= io_sc2mac_dat_bits_mask_59;
      end
    end
    if (_T_3014) begin
      _T_3555_60 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_60 <= io_sc2mac_dat_bits_mask_60;
      end
    end
    if (_T_3014) begin
      _T_3555_61 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_61 <= io_sc2mac_dat_bits_mask_61;
      end
    end
    if (_T_3014) begin
      _T_3555_62 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_62 <= io_sc2mac_dat_bits_mask_62;
      end
    end
    if (_T_3014) begin
      _T_3555_63 <= 1'h0;
    end else begin
      if (_T_5715) begin
        _T_3555_63 <= io_sc2mac_dat_bits_mask_63;
      end
    end
    if (_T_3014) begin
      _T_4018_0 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_0 <= _T_3555_0;
      end
    end
    if (_T_3014) begin
      _T_4018_1 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_1 <= _T_3555_1;
      end
    end
    if (_T_3014) begin
      _T_4018_2 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_2 <= _T_3555_2;
      end
    end
    if (_T_3014) begin
      _T_4018_3 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_3 <= _T_3555_3;
      end
    end
    if (_T_3014) begin
      _T_4018_4 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_4 <= _T_3555_4;
      end
    end
    if (_T_3014) begin
      _T_4018_5 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_5 <= _T_3555_5;
      end
    end
    if (_T_3014) begin
      _T_4018_6 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_6 <= _T_3555_6;
      end
    end
    if (_T_3014) begin
      _T_4018_7 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_7 <= _T_3555_7;
      end
    end
    if (_T_3014) begin
      _T_4018_8 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_8 <= _T_3555_8;
      end
    end
    if (_T_3014) begin
      _T_4018_9 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_9 <= _T_3555_9;
      end
    end
    if (_T_3014) begin
      _T_4018_10 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_10 <= _T_3555_10;
      end
    end
    if (_T_3014) begin
      _T_4018_11 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_11 <= _T_3555_11;
      end
    end
    if (_T_3014) begin
      _T_4018_12 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_12 <= _T_3555_12;
      end
    end
    if (_T_3014) begin
      _T_4018_13 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_13 <= _T_3555_13;
      end
    end
    if (_T_3014) begin
      _T_4018_14 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_14 <= _T_3555_14;
      end
    end
    if (_T_3014) begin
      _T_4018_15 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_15 <= _T_3555_15;
      end
    end
    if (_T_3014) begin
      _T_4018_16 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_16 <= _T_3555_16;
      end
    end
    if (_T_3014) begin
      _T_4018_17 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_17 <= _T_3555_17;
      end
    end
    if (_T_3014) begin
      _T_4018_18 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_18 <= _T_3555_18;
      end
    end
    if (_T_3014) begin
      _T_4018_19 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_19 <= _T_3555_19;
      end
    end
    if (_T_3014) begin
      _T_4018_20 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_20 <= _T_3555_20;
      end
    end
    if (_T_3014) begin
      _T_4018_21 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_21 <= _T_3555_21;
      end
    end
    if (_T_3014) begin
      _T_4018_22 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_22 <= _T_3555_22;
      end
    end
    if (_T_3014) begin
      _T_4018_23 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_23 <= _T_3555_23;
      end
    end
    if (_T_3014) begin
      _T_4018_24 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_24 <= _T_3555_24;
      end
    end
    if (_T_3014) begin
      _T_4018_25 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_25 <= _T_3555_25;
      end
    end
    if (_T_3014) begin
      _T_4018_26 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_26 <= _T_3555_26;
      end
    end
    if (_T_3014) begin
      _T_4018_27 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_27 <= _T_3555_27;
      end
    end
    if (_T_3014) begin
      _T_4018_28 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_28 <= _T_3555_28;
      end
    end
    if (_T_3014) begin
      _T_4018_29 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_29 <= _T_3555_29;
      end
    end
    if (_T_3014) begin
      _T_4018_30 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_30 <= _T_3555_30;
      end
    end
    if (_T_3014) begin
      _T_4018_31 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_31 <= _T_3555_31;
      end
    end
    if (_T_3014) begin
      _T_4018_32 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_32 <= _T_3555_32;
      end
    end
    if (_T_3014) begin
      _T_4018_33 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_33 <= _T_3555_33;
      end
    end
    if (_T_3014) begin
      _T_4018_34 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_34 <= _T_3555_34;
      end
    end
    if (_T_3014) begin
      _T_4018_35 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_35 <= _T_3555_35;
      end
    end
    if (_T_3014) begin
      _T_4018_36 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_36 <= _T_3555_36;
      end
    end
    if (_T_3014) begin
      _T_4018_37 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_37 <= _T_3555_37;
      end
    end
    if (_T_3014) begin
      _T_4018_38 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_38 <= _T_3555_38;
      end
    end
    if (_T_3014) begin
      _T_4018_39 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_39 <= _T_3555_39;
      end
    end
    if (_T_3014) begin
      _T_4018_40 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_40 <= _T_3555_40;
      end
    end
    if (_T_3014) begin
      _T_4018_41 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_41 <= _T_3555_41;
      end
    end
    if (_T_3014) begin
      _T_4018_42 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_42 <= _T_3555_42;
      end
    end
    if (_T_3014) begin
      _T_4018_43 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_43 <= _T_3555_43;
      end
    end
    if (_T_3014) begin
      _T_4018_44 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_44 <= _T_3555_44;
      end
    end
    if (_T_3014) begin
      _T_4018_45 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_45 <= _T_3555_45;
      end
    end
    if (_T_3014) begin
      _T_4018_46 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_46 <= _T_3555_46;
      end
    end
    if (_T_3014) begin
      _T_4018_47 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_47 <= _T_3555_47;
      end
    end
    if (_T_3014) begin
      _T_4018_48 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_48 <= _T_3555_48;
      end
    end
    if (_T_3014) begin
      _T_4018_49 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_49 <= _T_3555_49;
      end
    end
    if (_T_3014) begin
      _T_4018_50 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_50 <= _T_3555_50;
      end
    end
    if (_T_3014) begin
      _T_4018_51 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_51 <= _T_3555_51;
      end
    end
    if (_T_3014) begin
      _T_4018_52 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_52 <= _T_3555_52;
      end
    end
    if (_T_3014) begin
      _T_4018_53 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_53 <= _T_3555_53;
      end
    end
    if (_T_3014) begin
      _T_4018_54 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_54 <= _T_3555_54;
      end
    end
    if (_T_3014) begin
      _T_4018_55 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_55 <= _T_3555_55;
      end
    end
    if (_T_3014) begin
      _T_4018_56 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_56 <= _T_3555_56;
      end
    end
    if (_T_3014) begin
      _T_4018_57 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_57 <= _T_3555_57;
      end
    end
    if (_T_3014) begin
      _T_4018_58 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_58 <= _T_3555_58;
      end
    end
    if (_T_3014) begin
      _T_4018_59 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_59 <= _T_3555_59;
      end
    end
    if (_T_3014) begin
      _T_4018_60 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_60 <= _T_3555_60;
      end
    end
    if (_T_3014) begin
      _T_4018_61 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_61 <= _T_3555_61;
      end
    end
    if (_T_3014) begin
      _T_4018_62 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_62 <= _T_3555_62;
      end
    end
    if (_T_3014) begin
      _T_4018_63 <= 1'h0;
    end else begin
      if (_T_5717) begin
        _T_4018_63 <= _T_3555_63;
      end
    end
    if (_T_3014) begin
      _T_4219 <= 1'h0;
    end else begin
      _T_4219 <= io_sc2mac_dat_valid;
    end
    if (_T_3014) begin
      _T_4222 <= 1'h0;
    end else begin
      _T_4222 <= _T_4219;
    end
    if (_T_3014) begin
      _T_4227 <= 9'h0;
    end else begin
      if (_T_5715) begin
        _T_4227 <= io_sc2mac_dat_bits_pd;
      end
    end
    if (_T_3014) begin
      _T_4230 <= 9'h0;
    end else begin
      if (_T_5717) begin
        _T_4230 <= _T_4227;
      end
    end
    if (io_sc2mac_wt_bits_mask_0) begin
      _T_4301_0 <= io_sc2mac_wt_bits_data_0;
    end
    if (io_sc2mac_wt_bits_mask_1) begin
      _T_4301_1 <= io_sc2mac_wt_bits_data_1;
    end
    if (io_sc2mac_wt_bits_mask_2) begin
      _T_4301_2 <= io_sc2mac_wt_bits_data_2;
    end
    if (io_sc2mac_wt_bits_mask_3) begin
      _T_4301_3 <= io_sc2mac_wt_bits_data_3;
    end
    if (io_sc2mac_wt_bits_mask_4) begin
      _T_4301_4 <= io_sc2mac_wt_bits_data_4;
    end
    if (io_sc2mac_wt_bits_mask_5) begin
      _T_4301_5 <= io_sc2mac_wt_bits_data_5;
    end
    if (io_sc2mac_wt_bits_mask_6) begin
      _T_4301_6 <= io_sc2mac_wt_bits_data_6;
    end
    if (io_sc2mac_wt_bits_mask_7) begin
      _T_4301_7 <= io_sc2mac_wt_bits_data_7;
    end
    if (io_sc2mac_wt_bits_mask_8) begin
      _T_4301_8 <= io_sc2mac_wt_bits_data_8;
    end
    if (io_sc2mac_wt_bits_mask_9) begin
      _T_4301_9 <= io_sc2mac_wt_bits_data_9;
    end
    if (io_sc2mac_wt_bits_mask_10) begin
      _T_4301_10 <= io_sc2mac_wt_bits_data_10;
    end
    if (io_sc2mac_wt_bits_mask_11) begin
      _T_4301_11 <= io_sc2mac_wt_bits_data_11;
    end
    if (io_sc2mac_wt_bits_mask_12) begin
      _T_4301_12 <= io_sc2mac_wt_bits_data_12;
    end
    if (io_sc2mac_wt_bits_mask_13) begin
      _T_4301_13 <= io_sc2mac_wt_bits_data_13;
    end
    if (io_sc2mac_wt_bits_mask_14) begin
      _T_4301_14 <= io_sc2mac_wt_bits_data_14;
    end
    if (io_sc2mac_wt_bits_mask_15) begin
      _T_4301_15 <= io_sc2mac_wt_bits_data_15;
    end
    if (io_sc2mac_wt_bits_mask_16) begin
      _T_4301_16 <= io_sc2mac_wt_bits_data_16;
    end
    if (io_sc2mac_wt_bits_mask_17) begin
      _T_4301_17 <= io_sc2mac_wt_bits_data_17;
    end
    if (io_sc2mac_wt_bits_mask_18) begin
      _T_4301_18 <= io_sc2mac_wt_bits_data_18;
    end
    if (io_sc2mac_wt_bits_mask_19) begin
      _T_4301_19 <= io_sc2mac_wt_bits_data_19;
    end
    if (io_sc2mac_wt_bits_mask_20) begin
      _T_4301_20 <= io_sc2mac_wt_bits_data_20;
    end
    if (io_sc2mac_wt_bits_mask_21) begin
      _T_4301_21 <= io_sc2mac_wt_bits_data_21;
    end
    if (io_sc2mac_wt_bits_mask_22) begin
      _T_4301_22 <= io_sc2mac_wt_bits_data_22;
    end
    if (io_sc2mac_wt_bits_mask_23) begin
      _T_4301_23 <= io_sc2mac_wt_bits_data_23;
    end
    if (io_sc2mac_wt_bits_mask_24) begin
      _T_4301_24 <= io_sc2mac_wt_bits_data_24;
    end
    if (io_sc2mac_wt_bits_mask_25) begin
      _T_4301_25 <= io_sc2mac_wt_bits_data_25;
    end
    if (io_sc2mac_wt_bits_mask_26) begin
      _T_4301_26 <= io_sc2mac_wt_bits_data_26;
    end
    if (io_sc2mac_wt_bits_mask_27) begin
      _T_4301_27 <= io_sc2mac_wt_bits_data_27;
    end
    if (io_sc2mac_wt_bits_mask_28) begin
      _T_4301_28 <= io_sc2mac_wt_bits_data_28;
    end
    if (io_sc2mac_wt_bits_mask_29) begin
      _T_4301_29 <= io_sc2mac_wt_bits_data_29;
    end
    if (io_sc2mac_wt_bits_mask_30) begin
      _T_4301_30 <= io_sc2mac_wt_bits_data_30;
    end
    if (io_sc2mac_wt_bits_mask_31) begin
      _T_4301_31 <= io_sc2mac_wt_bits_data_31;
    end
    if (io_sc2mac_wt_bits_mask_32) begin
      _T_4301_32 <= io_sc2mac_wt_bits_data_32;
    end
    if (io_sc2mac_wt_bits_mask_33) begin
      _T_4301_33 <= io_sc2mac_wt_bits_data_33;
    end
    if (io_sc2mac_wt_bits_mask_34) begin
      _T_4301_34 <= io_sc2mac_wt_bits_data_34;
    end
    if (io_sc2mac_wt_bits_mask_35) begin
      _T_4301_35 <= io_sc2mac_wt_bits_data_35;
    end
    if (io_sc2mac_wt_bits_mask_36) begin
      _T_4301_36 <= io_sc2mac_wt_bits_data_36;
    end
    if (io_sc2mac_wt_bits_mask_37) begin
      _T_4301_37 <= io_sc2mac_wt_bits_data_37;
    end
    if (io_sc2mac_wt_bits_mask_38) begin
      _T_4301_38 <= io_sc2mac_wt_bits_data_38;
    end
    if (io_sc2mac_wt_bits_mask_39) begin
      _T_4301_39 <= io_sc2mac_wt_bits_data_39;
    end
    if (io_sc2mac_wt_bits_mask_40) begin
      _T_4301_40 <= io_sc2mac_wt_bits_data_40;
    end
    if (io_sc2mac_wt_bits_mask_41) begin
      _T_4301_41 <= io_sc2mac_wt_bits_data_41;
    end
    if (io_sc2mac_wt_bits_mask_42) begin
      _T_4301_42 <= io_sc2mac_wt_bits_data_42;
    end
    if (io_sc2mac_wt_bits_mask_43) begin
      _T_4301_43 <= io_sc2mac_wt_bits_data_43;
    end
    if (io_sc2mac_wt_bits_mask_44) begin
      _T_4301_44 <= io_sc2mac_wt_bits_data_44;
    end
    if (io_sc2mac_wt_bits_mask_45) begin
      _T_4301_45 <= io_sc2mac_wt_bits_data_45;
    end
    if (io_sc2mac_wt_bits_mask_46) begin
      _T_4301_46 <= io_sc2mac_wt_bits_data_46;
    end
    if (io_sc2mac_wt_bits_mask_47) begin
      _T_4301_47 <= io_sc2mac_wt_bits_data_47;
    end
    if (io_sc2mac_wt_bits_mask_48) begin
      _T_4301_48 <= io_sc2mac_wt_bits_data_48;
    end
    if (io_sc2mac_wt_bits_mask_49) begin
      _T_4301_49 <= io_sc2mac_wt_bits_data_49;
    end
    if (io_sc2mac_wt_bits_mask_50) begin
      _T_4301_50 <= io_sc2mac_wt_bits_data_50;
    end
    if (io_sc2mac_wt_bits_mask_51) begin
      _T_4301_51 <= io_sc2mac_wt_bits_data_51;
    end
    if (io_sc2mac_wt_bits_mask_52) begin
      _T_4301_52 <= io_sc2mac_wt_bits_data_52;
    end
    if (io_sc2mac_wt_bits_mask_53) begin
      _T_4301_53 <= io_sc2mac_wt_bits_data_53;
    end
    if (io_sc2mac_wt_bits_mask_54) begin
      _T_4301_54 <= io_sc2mac_wt_bits_data_54;
    end
    if (io_sc2mac_wt_bits_mask_55) begin
      _T_4301_55 <= io_sc2mac_wt_bits_data_55;
    end
    if (io_sc2mac_wt_bits_mask_56) begin
      _T_4301_56 <= io_sc2mac_wt_bits_data_56;
    end
    if (io_sc2mac_wt_bits_mask_57) begin
      _T_4301_57 <= io_sc2mac_wt_bits_data_57;
    end
    if (io_sc2mac_wt_bits_mask_58) begin
      _T_4301_58 <= io_sc2mac_wt_bits_data_58;
    end
    if (io_sc2mac_wt_bits_mask_59) begin
      _T_4301_59 <= io_sc2mac_wt_bits_data_59;
    end
    if (io_sc2mac_wt_bits_mask_60) begin
      _T_4301_60 <= io_sc2mac_wt_bits_data_60;
    end
    if (io_sc2mac_wt_bits_mask_61) begin
      _T_4301_61 <= io_sc2mac_wt_bits_data_61;
    end
    if (io_sc2mac_wt_bits_mask_62) begin
      _T_4301_62 <= io_sc2mac_wt_bits_data_62;
    end
    if (io_sc2mac_wt_bits_mask_63) begin
      _T_4301_63 <= io_sc2mac_wt_bits_data_63;
    end
    if (_T_4771_0) begin
      _T_4368_0 <= _T_4301_0;
    end
    if (_T_4771_1) begin
      _T_4368_1 <= _T_4301_1;
    end
    if (_T_4771_2) begin
      _T_4368_2 <= _T_4301_2;
    end
    if (_T_4771_3) begin
      _T_4368_3 <= _T_4301_3;
    end
    if (_T_4771_4) begin
      _T_4368_4 <= _T_4301_4;
    end
    if (_T_4771_5) begin
      _T_4368_5 <= _T_4301_5;
    end
    if (_T_4771_6) begin
      _T_4368_6 <= _T_4301_6;
    end
    if (_T_4771_7) begin
      _T_4368_7 <= _T_4301_7;
    end
    if (_T_4771_8) begin
      _T_4368_8 <= _T_4301_8;
    end
    if (_T_4771_9) begin
      _T_4368_9 <= _T_4301_9;
    end
    if (_T_4771_10) begin
      _T_4368_10 <= _T_4301_10;
    end
    if (_T_4771_11) begin
      _T_4368_11 <= _T_4301_11;
    end
    if (_T_4771_12) begin
      _T_4368_12 <= _T_4301_12;
    end
    if (_T_4771_13) begin
      _T_4368_13 <= _T_4301_13;
    end
    if (_T_4771_14) begin
      _T_4368_14 <= _T_4301_14;
    end
    if (_T_4771_15) begin
      _T_4368_15 <= _T_4301_15;
    end
    if (_T_4771_16) begin
      _T_4368_16 <= _T_4301_16;
    end
    if (_T_4771_17) begin
      _T_4368_17 <= _T_4301_17;
    end
    if (_T_4771_18) begin
      _T_4368_18 <= _T_4301_18;
    end
    if (_T_4771_19) begin
      _T_4368_19 <= _T_4301_19;
    end
    if (_T_4771_20) begin
      _T_4368_20 <= _T_4301_20;
    end
    if (_T_4771_21) begin
      _T_4368_21 <= _T_4301_21;
    end
    if (_T_4771_22) begin
      _T_4368_22 <= _T_4301_22;
    end
    if (_T_4771_23) begin
      _T_4368_23 <= _T_4301_23;
    end
    if (_T_4771_24) begin
      _T_4368_24 <= _T_4301_24;
    end
    if (_T_4771_25) begin
      _T_4368_25 <= _T_4301_25;
    end
    if (_T_4771_26) begin
      _T_4368_26 <= _T_4301_26;
    end
    if (_T_4771_27) begin
      _T_4368_27 <= _T_4301_27;
    end
    if (_T_4771_28) begin
      _T_4368_28 <= _T_4301_28;
    end
    if (_T_4771_29) begin
      _T_4368_29 <= _T_4301_29;
    end
    if (_T_4771_30) begin
      _T_4368_30 <= _T_4301_30;
    end
    if (_T_4771_31) begin
      _T_4368_31 <= _T_4301_31;
    end
    if (_T_4771_32) begin
      _T_4368_32 <= _T_4301_32;
    end
    if (_T_4771_33) begin
      _T_4368_33 <= _T_4301_33;
    end
    if (_T_4771_34) begin
      _T_4368_34 <= _T_4301_34;
    end
    if (_T_4771_35) begin
      _T_4368_35 <= _T_4301_35;
    end
    if (_T_4771_36) begin
      _T_4368_36 <= _T_4301_36;
    end
    if (_T_4771_37) begin
      _T_4368_37 <= _T_4301_37;
    end
    if (_T_4771_38) begin
      _T_4368_38 <= _T_4301_38;
    end
    if (_T_4771_39) begin
      _T_4368_39 <= _T_4301_39;
    end
    if (_T_4771_40) begin
      _T_4368_40 <= _T_4301_40;
    end
    if (_T_4771_41) begin
      _T_4368_41 <= _T_4301_41;
    end
    if (_T_4771_42) begin
      _T_4368_42 <= _T_4301_42;
    end
    if (_T_4771_43) begin
      _T_4368_43 <= _T_4301_43;
    end
    if (_T_4771_44) begin
      _T_4368_44 <= _T_4301_44;
    end
    if (_T_4771_45) begin
      _T_4368_45 <= _T_4301_45;
    end
    if (_T_4771_46) begin
      _T_4368_46 <= _T_4301_46;
    end
    if (_T_4771_47) begin
      _T_4368_47 <= _T_4301_47;
    end
    if (_T_4771_48) begin
      _T_4368_48 <= _T_4301_48;
    end
    if (_T_4771_49) begin
      _T_4368_49 <= _T_4301_49;
    end
    if (_T_4771_50) begin
      _T_4368_50 <= _T_4301_50;
    end
    if (_T_4771_51) begin
      _T_4368_51 <= _T_4301_51;
    end
    if (_T_4771_52) begin
      _T_4368_52 <= _T_4301_52;
    end
    if (_T_4771_53) begin
      _T_4368_53 <= _T_4301_53;
    end
    if (_T_4771_54) begin
      _T_4368_54 <= _T_4301_54;
    end
    if (_T_4771_55) begin
      _T_4368_55 <= _T_4301_55;
    end
    if (_T_4771_56) begin
      _T_4368_56 <= _T_4301_56;
    end
    if (_T_4771_57) begin
      _T_4368_57 <= _T_4301_57;
    end
    if (_T_4771_58) begin
      _T_4368_58 <= _T_4301_58;
    end
    if (_T_4771_59) begin
      _T_4368_59 <= _T_4301_59;
    end
    if (_T_4771_60) begin
      _T_4368_60 <= _T_4301_60;
    end
    if (_T_4771_61) begin
      _T_4368_61 <= _T_4301_61;
    end
    if (_T_4771_62) begin
      _T_4368_62 <= _T_4301_62;
    end
    if (_T_4771_63) begin
      _T_4368_63 <= _T_4301_63;
    end
    if (_T_3014) begin
      _T_4771_0 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_0 <= io_sc2mac_wt_bits_mask_0;
      end
    end
    if (_T_3014) begin
      _T_4771_1 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_1 <= io_sc2mac_wt_bits_mask_1;
      end
    end
    if (_T_3014) begin
      _T_4771_2 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_2 <= io_sc2mac_wt_bits_mask_2;
      end
    end
    if (_T_3014) begin
      _T_4771_3 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_3 <= io_sc2mac_wt_bits_mask_3;
      end
    end
    if (_T_3014) begin
      _T_4771_4 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_4 <= io_sc2mac_wt_bits_mask_4;
      end
    end
    if (_T_3014) begin
      _T_4771_5 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_5 <= io_sc2mac_wt_bits_mask_5;
      end
    end
    if (_T_3014) begin
      _T_4771_6 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_6 <= io_sc2mac_wt_bits_mask_6;
      end
    end
    if (_T_3014) begin
      _T_4771_7 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_7 <= io_sc2mac_wt_bits_mask_7;
      end
    end
    if (_T_3014) begin
      _T_4771_8 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_8 <= io_sc2mac_wt_bits_mask_8;
      end
    end
    if (_T_3014) begin
      _T_4771_9 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_9 <= io_sc2mac_wt_bits_mask_9;
      end
    end
    if (_T_3014) begin
      _T_4771_10 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_10 <= io_sc2mac_wt_bits_mask_10;
      end
    end
    if (_T_3014) begin
      _T_4771_11 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_11 <= io_sc2mac_wt_bits_mask_11;
      end
    end
    if (_T_3014) begin
      _T_4771_12 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_12 <= io_sc2mac_wt_bits_mask_12;
      end
    end
    if (_T_3014) begin
      _T_4771_13 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_13 <= io_sc2mac_wt_bits_mask_13;
      end
    end
    if (_T_3014) begin
      _T_4771_14 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_14 <= io_sc2mac_wt_bits_mask_14;
      end
    end
    if (_T_3014) begin
      _T_4771_15 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_15 <= io_sc2mac_wt_bits_mask_15;
      end
    end
    if (_T_3014) begin
      _T_4771_16 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_16 <= io_sc2mac_wt_bits_mask_16;
      end
    end
    if (_T_3014) begin
      _T_4771_17 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_17 <= io_sc2mac_wt_bits_mask_17;
      end
    end
    if (_T_3014) begin
      _T_4771_18 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_18 <= io_sc2mac_wt_bits_mask_18;
      end
    end
    if (_T_3014) begin
      _T_4771_19 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_19 <= io_sc2mac_wt_bits_mask_19;
      end
    end
    if (_T_3014) begin
      _T_4771_20 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_20 <= io_sc2mac_wt_bits_mask_20;
      end
    end
    if (_T_3014) begin
      _T_4771_21 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_21 <= io_sc2mac_wt_bits_mask_21;
      end
    end
    if (_T_3014) begin
      _T_4771_22 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_22 <= io_sc2mac_wt_bits_mask_22;
      end
    end
    if (_T_3014) begin
      _T_4771_23 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_23 <= io_sc2mac_wt_bits_mask_23;
      end
    end
    if (_T_3014) begin
      _T_4771_24 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_24 <= io_sc2mac_wt_bits_mask_24;
      end
    end
    if (_T_3014) begin
      _T_4771_25 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_25 <= io_sc2mac_wt_bits_mask_25;
      end
    end
    if (_T_3014) begin
      _T_4771_26 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_26 <= io_sc2mac_wt_bits_mask_26;
      end
    end
    if (_T_3014) begin
      _T_4771_27 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_27 <= io_sc2mac_wt_bits_mask_27;
      end
    end
    if (_T_3014) begin
      _T_4771_28 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_28 <= io_sc2mac_wt_bits_mask_28;
      end
    end
    if (_T_3014) begin
      _T_4771_29 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_29 <= io_sc2mac_wt_bits_mask_29;
      end
    end
    if (_T_3014) begin
      _T_4771_30 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_30 <= io_sc2mac_wt_bits_mask_30;
      end
    end
    if (_T_3014) begin
      _T_4771_31 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_31 <= io_sc2mac_wt_bits_mask_31;
      end
    end
    if (_T_3014) begin
      _T_4771_32 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_32 <= io_sc2mac_wt_bits_mask_32;
      end
    end
    if (_T_3014) begin
      _T_4771_33 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_33 <= io_sc2mac_wt_bits_mask_33;
      end
    end
    if (_T_3014) begin
      _T_4771_34 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_34 <= io_sc2mac_wt_bits_mask_34;
      end
    end
    if (_T_3014) begin
      _T_4771_35 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_35 <= io_sc2mac_wt_bits_mask_35;
      end
    end
    if (_T_3014) begin
      _T_4771_36 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_36 <= io_sc2mac_wt_bits_mask_36;
      end
    end
    if (_T_3014) begin
      _T_4771_37 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_37 <= io_sc2mac_wt_bits_mask_37;
      end
    end
    if (_T_3014) begin
      _T_4771_38 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_38 <= io_sc2mac_wt_bits_mask_38;
      end
    end
    if (_T_3014) begin
      _T_4771_39 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_39 <= io_sc2mac_wt_bits_mask_39;
      end
    end
    if (_T_3014) begin
      _T_4771_40 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_40 <= io_sc2mac_wt_bits_mask_40;
      end
    end
    if (_T_3014) begin
      _T_4771_41 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_41 <= io_sc2mac_wt_bits_mask_41;
      end
    end
    if (_T_3014) begin
      _T_4771_42 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_42 <= io_sc2mac_wt_bits_mask_42;
      end
    end
    if (_T_3014) begin
      _T_4771_43 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_43 <= io_sc2mac_wt_bits_mask_43;
      end
    end
    if (_T_3014) begin
      _T_4771_44 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_44 <= io_sc2mac_wt_bits_mask_44;
      end
    end
    if (_T_3014) begin
      _T_4771_45 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_45 <= io_sc2mac_wt_bits_mask_45;
      end
    end
    if (_T_3014) begin
      _T_4771_46 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_46 <= io_sc2mac_wt_bits_mask_46;
      end
    end
    if (_T_3014) begin
      _T_4771_47 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_47 <= io_sc2mac_wt_bits_mask_47;
      end
    end
    if (_T_3014) begin
      _T_4771_48 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_48 <= io_sc2mac_wt_bits_mask_48;
      end
    end
    if (_T_3014) begin
      _T_4771_49 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_49 <= io_sc2mac_wt_bits_mask_49;
      end
    end
    if (_T_3014) begin
      _T_4771_50 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_50 <= io_sc2mac_wt_bits_mask_50;
      end
    end
    if (_T_3014) begin
      _T_4771_51 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_51 <= io_sc2mac_wt_bits_mask_51;
      end
    end
    if (_T_3014) begin
      _T_4771_52 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_52 <= io_sc2mac_wt_bits_mask_52;
      end
    end
    if (_T_3014) begin
      _T_4771_53 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_53 <= io_sc2mac_wt_bits_mask_53;
      end
    end
    if (_T_3014) begin
      _T_4771_54 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_54 <= io_sc2mac_wt_bits_mask_54;
      end
    end
    if (_T_3014) begin
      _T_4771_55 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_55 <= io_sc2mac_wt_bits_mask_55;
      end
    end
    if (_T_3014) begin
      _T_4771_56 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_56 <= io_sc2mac_wt_bits_mask_56;
      end
    end
    if (_T_3014) begin
      _T_4771_57 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_57 <= io_sc2mac_wt_bits_mask_57;
      end
    end
    if (_T_3014) begin
      _T_4771_58 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_58 <= io_sc2mac_wt_bits_mask_58;
      end
    end
    if (_T_3014) begin
      _T_4771_59 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_59 <= io_sc2mac_wt_bits_mask_59;
      end
    end
    if (_T_3014) begin
      _T_4771_60 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_60 <= io_sc2mac_wt_bits_mask_60;
      end
    end
    if (_T_3014) begin
      _T_4771_61 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_61 <= io_sc2mac_wt_bits_mask_61;
      end
    end
    if (_T_3014) begin
      _T_4771_62 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_62 <= io_sc2mac_wt_bits_mask_62;
      end
    end
    if (_T_3014) begin
      _T_4771_63 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_4771_63 <= io_sc2mac_wt_bits_mask_63;
      end
    end
    if (_T_3014) begin
      _T_5234_0 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_0 <= _T_4771_0;
      end
    end
    if (_T_3014) begin
      _T_5234_1 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_1 <= _T_4771_1;
      end
    end
    if (_T_3014) begin
      _T_5234_2 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_2 <= _T_4771_2;
      end
    end
    if (_T_3014) begin
      _T_5234_3 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_3 <= _T_4771_3;
      end
    end
    if (_T_3014) begin
      _T_5234_4 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_4 <= _T_4771_4;
      end
    end
    if (_T_3014) begin
      _T_5234_5 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_5 <= _T_4771_5;
      end
    end
    if (_T_3014) begin
      _T_5234_6 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_6 <= _T_4771_6;
      end
    end
    if (_T_3014) begin
      _T_5234_7 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_7 <= _T_4771_7;
      end
    end
    if (_T_3014) begin
      _T_5234_8 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_8 <= _T_4771_8;
      end
    end
    if (_T_3014) begin
      _T_5234_9 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_9 <= _T_4771_9;
      end
    end
    if (_T_3014) begin
      _T_5234_10 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_10 <= _T_4771_10;
      end
    end
    if (_T_3014) begin
      _T_5234_11 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_11 <= _T_4771_11;
      end
    end
    if (_T_3014) begin
      _T_5234_12 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_12 <= _T_4771_12;
      end
    end
    if (_T_3014) begin
      _T_5234_13 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_13 <= _T_4771_13;
      end
    end
    if (_T_3014) begin
      _T_5234_14 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_14 <= _T_4771_14;
      end
    end
    if (_T_3014) begin
      _T_5234_15 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_15 <= _T_4771_15;
      end
    end
    if (_T_3014) begin
      _T_5234_16 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_16 <= _T_4771_16;
      end
    end
    if (_T_3014) begin
      _T_5234_17 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_17 <= _T_4771_17;
      end
    end
    if (_T_3014) begin
      _T_5234_18 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_18 <= _T_4771_18;
      end
    end
    if (_T_3014) begin
      _T_5234_19 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_19 <= _T_4771_19;
      end
    end
    if (_T_3014) begin
      _T_5234_20 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_20 <= _T_4771_20;
      end
    end
    if (_T_3014) begin
      _T_5234_21 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_21 <= _T_4771_21;
      end
    end
    if (_T_3014) begin
      _T_5234_22 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_22 <= _T_4771_22;
      end
    end
    if (_T_3014) begin
      _T_5234_23 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_23 <= _T_4771_23;
      end
    end
    if (_T_3014) begin
      _T_5234_24 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_24 <= _T_4771_24;
      end
    end
    if (_T_3014) begin
      _T_5234_25 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_25 <= _T_4771_25;
      end
    end
    if (_T_3014) begin
      _T_5234_26 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_26 <= _T_4771_26;
      end
    end
    if (_T_3014) begin
      _T_5234_27 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_27 <= _T_4771_27;
      end
    end
    if (_T_3014) begin
      _T_5234_28 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_28 <= _T_4771_28;
      end
    end
    if (_T_3014) begin
      _T_5234_29 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_29 <= _T_4771_29;
      end
    end
    if (_T_3014) begin
      _T_5234_30 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_30 <= _T_4771_30;
      end
    end
    if (_T_3014) begin
      _T_5234_31 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_31 <= _T_4771_31;
      end
    end
    if (_T_3014) begin
      _T_5234_32 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_32 <= _T_4771_32;
      end
    end
    if (_T_3014) begin
      _T_5234_33 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_33 <= _T_4771_33;
      end
    end
    if (_T_3014) begin
      _T_5234_34 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_34 <= _T_4771_34;
      end
    end
    if (_T_3014) begin
      _T_5234_35 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_35 <= _T_4771_35;
      end
    end
    if (_T_3014) begin
      _T_5234_36 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_36 <= _T_4771_36;
      end
    end
    if (_T_3014) begin
      _T_5234_37 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_37 <= _T_4771_37;
      end
    end
    if (_T_3014) begin
      _T_5234_38 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_38 <= _T_4771_38;
      end
    end
    if (_T_3014) begin
      _T_5234_39 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_39 <= _T_4771_39;
      end
    end
    if (_T_3014) begin
      _T_5234_40 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_40 <= _T_4771_40;
      end
    end
    if (_T_3014) begin
      _T_5234_41 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_41 <= _T_4771_41;
      end
    end
    if (_T_3014) begin
      _T_5234_42 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_42 <= _T_4771_42;
      end
    end
    if (_T_3014) begin
      _T_5234_43 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_43 <= _T_4771_43;
      end
    end
    if (_T_3014) begin
      _T_5234_44 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_44 <= _T_4771_44;
      end
    end
    if (_T_3014) begin
      _T_5234_45 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_45 <= _T_4771_45;
      end
    end
    if (_T_3014) begin
      _T_5234_46 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_46 <= _T_4771_46;
      end
    end
    if (_T_3014) begin
      _T_5234_47 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_47 <= _T_4771_47;
      end
    end
    if (_T_3014) begin
      _T_5234_48 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_48 <= _T_4771_48;
      end
    end
    if (_T_3014) begin
      _T_5234_49 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_49 <= _T_4771_49;
      end
    end
    if (_T_3014) begin
      _T_5234_50 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_50 <= _T_4771_50;
      end
    end
    if (_T_3014) begin
      _T_5234_51 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_51 <= _T_4771_51;
      end
    end
    if (_T_3014) begin
      _T_5234_52 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_52 <= _T_4771_52;
      end
    end
    if (_T_3014) begin
      _T_5234_53 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_53 <= _T_4771_53;
      end
    end
    if (_T_3014) begin
      _T_5234_54 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_54 <= _T_4771_54;
      end
    end
    if (_T_3014) begin
      _T_5234_55 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_55 <= _T_4771_55;
      end
    end
    if (_T_3014) begin
      _T_5234_56 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_56 <= _T_4771_56;
      end
    end
    if (_T_3014) begin
      _T_5234_57 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_57 <= _T_4771_57;
      end
    end
    if (_T_3014) begin
      _T_5234_58 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_58 <= _T_4771_58;
      end
    end
    if (_T_3014) begin
      _T_5234_59 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_59 <= _T_4771_59;
      end
    end
    if (_T_3014) begin
      _T_5234_60 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_60 <= _T_4771_60;
      end
    end
    if (_T_3014) begin
      _T_5234_61 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_61 <= _T_4771_61;
      end
    end
    if (_T_3014) begin
      _T_5234_62 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_62 <= _T_4771_62;
      end
    end
    if (_T_3014) begin
      _T_5234_63 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5234_63 <= _T_4771_63;
      end
    end
    if (_T_3014) begin
      _T_5435 <= 1'h0;
    end else begin
      _T_5435 <= io_sc2mac_wt_valid;
    end
    if (_T_3014) begin
      _T_5438 <= 1'h0;
    end else begin
      _T_5438 <= _T_5435;
    end
    if (_T_3014) begin
      _T_5535_0 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_5535_0 <= io_sc2mac_wt_bits_sel_0;
      end
    end
    if (_T_3014) begin
      _T_5535_1 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_5535_1 <= io_sc2mac_wt_bits_sel_1;
      end
    end
    if (_T_3014) begin
      _T_5535_2 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_5535_2 <= io_sc2mac_wt_bits_sel_2;
      end
    end
    if (_T_3014) begin
      _T_5535_3 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_5535_3 <= io_sc2mac_wt_bits_sel_3;
      end
    end
    if (_T_3014) begin
      _T_5535_4 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_5535_4 <= io_sc2mac_wt_bits_sel_4;
      end
    end
    if (_T_3014) begin
      _T_5535_5 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_5535_5 <= io_sc2mac_wt_bits_sel_5;
      end
    end
    if (_T_3014) begin
      _T_5535_6 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_5535_6 <= io_sc2mac_wt_bits_sel_6;
      end
    end
    if (_T_3014) begin
      _T_5535_7 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_5535_7 <= io_sc2mac_wt_bits_sel_7;
      end
    end
    if (_T_3014) begin
      _T_5535_8 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_5535_8 <= io_sc2mac_wt_bits_sel_8;
      end
    end
    if (_T_3014) begin
      _T_5535_9 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_5535_9 <= io_sc2mac_wt_bits_sel_9;
      end
    end
    if (_T_3014) begin
      _T_5535_10 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_5535_10 <= io_sc2mac_wt_bits_sel_10;
      end
    end
    if (_T_3014) begin
      _T_5535_11 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_5535_11 <= io_sc2mac_wt_bits_sel_11;
      end
    end
    if (_T_3014) begin
      _T_5535_12 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_5535_12 <= io_sc2mac_wt_bits_sel_12;
      end
    end
    if (_T_3014) begin
      _T_5535_13 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_5535_13 <= io_sc2mac_wt_bits_sel_13;
      end
    end
    if (_T_3014) begin
      _T_5535_14 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_5535_14 <= io_sc2mac_wt_bits_sel_14;
      end
    end
    if (_T_3014) begin
      _T_5535_15 <= 1'h0;
    end else begin
      if (_T_5716) begin
        _T_5535_15 <= io_sc2mac_wt_bits_sel_15;
      end
    end
    if (_T_3014) begin
      _T_5662_0 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5662_0 <= _T_5535_0;
      end
    end
    if (_T_3014) begin
      _T_5662_1 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5662_1 <= _T_5535_1;
      end
    end
    if (_T_3014) begin
      _T_5662_2 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5662_2 <= _T_5535_2;
      end
    end
    if (_T_3014) begin
      _T_5662_3 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5662_3 <= _T_5535_3;
      end
    end
    if (_T_3014) begin
      _T_5662_4 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5662_4 <= _T_5535_4;
      end
    end
    if (_T_3014) begin
      _T_5662_5 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5662_5 <= _T_5535_5;
      end
    end
    if (_T_3014) begin
      _T_5662_6 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5662_6 <= _T_5535_6;
      end
    end
    if (_T_3014) begin
      _T_5662_7 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5662_7 <= _T_5535_7;
      end
    end
    if (_T_3014) begin
      _T_5662_8 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5662_8 <= _T_5535_8;
      end
    end
    if (_T_3014) begin
      _T_5662_9 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5662_9 <= _T_5535_9;
      end
    end
    if (_T_3014) begin
      _T_5662_10 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5662_10 <= _T_5535_10;
      end
    end
    if (_T_3014) begin
      _T_5662_11 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5662_11 <= _T_5535_11;
      end
    end
    if (_T_3014) begin
      _T_5662_12 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5662_12 <= _T_5535_12;
      end
    end
    if (_T_3014) begin
      _T_5662_13 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5662_13 <= _T_5535_13;
      end
    end
    if (_T_3014) begin
      _T_5662_14 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5662_14 <= _T_5535_14;
      end
    end
    if (_T_3014) begin
      _T_5662_15 <= 1'h0;
    end else begin
      if (_T_5718) begin
        _T_5662_15 <= _T_5535_15;
      end
    end
  end
endmodule
