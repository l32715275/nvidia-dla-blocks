module NV_NVDLA_CMAC_CORE_mac_dft( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input         io_nvdla_core_clk, // @[:@6.4]
  input         io_nvdla_core_rstn, // @[:@6.4]
  input         io_dat_actv_0_valid, // @[:@6.4]
  input         io_dat_actv_0_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_0_bits_data, // @[:@6.4]
  input         io_dat_actv_1_valid, // @[:@6.4]
  input         io_dat_actv_1_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_1_bits_data, // @[:@6.4]
  input         io_dat_actv_2_valid, // @[:@6.4]
  input         io_dat_actv_2_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_2_bits_data, // @[:@6.4]
  input         io_dat_actv_3_valid, // @[:@6.4]
  input         io_dat_actv_3_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_3_bits_data, // @[:@6.4]
  input         io_dat_actv_4_valid, // @[:@6.4]
  input         io_dat_actv_4_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_4_bits_data, // @[:@6.4]
  input         io_dat_actv_5_valid, // @[:@6.4]
  input         io_dat_actv_5_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_5_bits_data, // @[:@6.4]
  input         io_dat_actv_6_valid, // @[:@6.4]
  input         io_dat_actv_6_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_6_bits_data, // @[:@6.4]
  input         io_dat_actv_7_valid, // @[:@6.4]
  input         io_dat_actv_7_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_7_bits_data, // @[:@6.4]
  input         io_dat_actv_8_valid, // @[:@6.4]
  input         io_dat_actv_8_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_8_bits_data, // @[:@6.4]
  input         io_dat_actv_9_valid, // @[:@6.4]
  input         io_dat_actv_9_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_9_bits_data, // @[:@6.4]
  input         io_dat_actv_10_valid, // @[:@6.4]
  input         io_dat_actv_10_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_10_bits_data, // @[:@6.4]
  input         io_dat_actv_11_valid, // @[:@6.4]
  input         io_dat_actv_11_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_11_bits_data, // @[:@6.4]
  input         io_dat_actv_12_valid, // @[:@6.4]
  input         io_dat_actv_12_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_12_bits_data, // @[:@6.4]
  input         io_dat_actv_13_valid, // @[:@6.4]
  input         io_dat_actv_13_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_13_bits_data, // @[:@6.4]
  input         io_dat_actv_14_valid, // @[:@6.4]
  input         io_dat_actv_14_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_14_bits_data, // @[:@6.4]
  input         io_dat_actv_15_valid, // @[:@6.4]
  input         io_dat_actv_15_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_15_bits_data, // @[:@6.4]
  input         io_dat_actv_16_valid, // @[:@6.4]
  input         io_dat_actv_16_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_16_bits_data, // @[:@6.4]
  input         io_dat_actv_17_valid, // @[:@6.4]
  input         io_dat_actv_17_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_17_bits_data, // @[:@6.4]
  input         io_dat_actv_18_valid, // @[:@6.4]
  input         io_dat_actv_18_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_18_bits_data, // @[:@6.4]
  input         io_dat_actv_19_valid, // @[:@6.4]
  input         io_dat_actv_19_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_19_bits_data, // @[:@6.4]
  input         io_dat_actv_20_valid, // @[:@6.4]
  input         io_dat_actv_20_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_20_bits_data, // @[:@6.4]
  input         io_dat_actv_21_valid, // @[:@6.4]
  input         io_dat_actv_21_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_21_bits_data, // @[:@6.4]
  input         io_dat_actv_22_valid, // @[:@6.4]
  input         io_dat_actv_22_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_22_bits_data, // @[:@6.4]
  input         io_dat_actv_23_valid, // @[:@6.4]
  input         io_dat_actv_23_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_23_bits_data, // @[:@6.4]
  input         io_dat_actv_24_valid, // @[:@6.4]
  input         io_dat_actv_24_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_24_bits_data, // @[:@6.4]
  input         io_dat_actv_25_valid, // @[:@6.4]
  input         io_dat_actv_25_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_25_bits_data, // @[:@6.4]
  input         io_dat_actv_26_valid, // @[:@6.4]
  input         io_dat_actv_26_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_26_bits_data, // @[:@6.4]
  input         io_dat_actv_27_valid, // @[:@6.4]
  input         io_dat_actv_27_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_27_bits_data, // @[:@6.4]
  input         io_dat_actv_28_valid, // @[:@6.4]
  input         io_dat_actv_28_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_28_bits_data, // @[:@6.4]
  input         io_dat_actv_29_valid, // @[:@6.4]
  input         io_dat_actv_29_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_29_bits_data, // @[:@6.4]
  input         io_dat_actv_30_valid, // @[:@6.4]
  input         io_dat_actv_30_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_30_bits_data, // @[:@6.4]
  input         io_dat_actv_31_valid, // @[:@6.4]
  input         io_dat_actv_31_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_31_bits_data, // @[:@6.4]
  input         io_dat_actv_32_valid, // @[:@6.4]
  input         io_dat_actv_32_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_32_bits_data, // @[:@6.4]
  input         io_dat_actv_33_valid, // @[:@6.4]
  input         io_dat_actv_33_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_33_bits_data, // @[:@6.4]
  input         io_dat_actv_34_valid, // @[:@6.4]
  input         io_dat_actv_34_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_34_bits_data, // @[:@6.4]
  input         io_dat_actv_35_valid, // @[:@6.4]
  input         io_dat_actv_35_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_35_bits_data, // @[:@6.4]
  input         io_dat_actv_36_valid, // @[:@6.4]
  input         io_dat_actv_36_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_36_bits_data, // @[:@6.4]
  input         io_dat_actv_37_valid, // @[:@6.4]
  input         io_dat_actv_37_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_37_bits_data, // @[:@6.4]
  input         io_dat_actv_38_valid, // @[:@6.4]
  input         io_dat_actv_38_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_38_bits_data, // @[:@6.4]
  input         io_dat_actv_39_valid, // @[:@6.4]
  input         io_dat_actv_39_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_39_bits_data, // @[:@6.4]
  input         io_dat_actv_40_valid, // @[:@6.4]
  input         io_dat_actv_40_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_40_bits_data, // @[:@6.4]
  input         io_dat_actv_41_valid, // @[:@6.4]
  input         io_dat_actv_41_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_41_bits_data, // @[:@6.4]
  input         io_dat_actv_42_valid, // @[:@6.4]
  input         io_dat_actv_42_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_42_bits_data, // @[:@6.4]
  input         io_dat_actv_43_valid, // @[:@6.4]
  input         io_dat_actv_43_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_43_bits_data, // @[:@6.4]
  input         io_dat_actv_44_valid, // @[:@6.4]
  input         io_dat_actv_44_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_44_bits_data, // @[:@6.4]
  input         io_dat_actv_45_valid, // @[:@6.4]
  input         io_dat_actv_45_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_45_bits_data, // @[:@6.4]
  input         io_dat_actv_46_valid, // @[:@6.4]
  input         io_dat_actv_46_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_46_bits_data, // @[:@6.4]
  input         io_dat_actv_47_valid, // @[:@6.4]
  input         io_dat_actv_47_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_47_bits_data, // @[:@6.4]
  input         io_dat_actv_48_valid, // @[:@6.4]
  input         io_dat_actv_48_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_48_bits_data, // @[:@6.4]
  input         io_dat_actv_49_valid, // @[:@6.4]
  input         io_dat_actv_49_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_49_bits_data, // @[:@6.4]
  input         io_dat_actv_50_valid, // @[:@6.4]
  input         io_dat_actv_50_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_50_bits_data, // @[:@6.4]
  input         io_dat_actv_51_valid, // @[:@6.4]
  input         io_dat_actv_51_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_51_bits_data, // @[:@6.4]
  input         io_dat_actv_52_valid, // @[:@6.4]
  input         io_dat_actv_52_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_52_bits_data, // @[:@6.4]
  input         io_dat_actv_53_valid, // @[:@6.4]
  input         io_dat_actv_53_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_53_bits_data, // @[:@6.4]
  input         io_dat_actv_54_valid, // @[:@6.4]
  input         io_dat_actv_54_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_54_bits_data, // @[:@6.4]
  input         io_dat_actv_55_valid, // @[:@6.4]
  input         io_dat_actv_55_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_55_bits_data, // @[:@6.4]
  input         io_dat_actv_56_valid, // @[:@6.4]
  input         io_dat_actv_56_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_56_bits_data, // @[:@6.4]
  input         io_dat_actv_57_valid, // @[:@6.4]
  input         io_dat_actv_57_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_57_bits_data, // @[:@6.4]
  input         io_dat_actv_58_valid, // @[:@6.4]
  input         io_dat_actv_58_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_58_bits_data, // @[:@6.4]
  input         io_dat_actv_59_valid, // @[:@6.4]
  input         io_dat_actv_59_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_59_bits_data, // @[:@6.4]
  input         io_dat_actv_60_valid, // @[:@6.4]
  input         io_dat_actv_60_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_60_bits_data, // @[:@6.4]
  input         io_dat_actv_61_valid, // @[:@6.4]
  input         io_dat_actv_61_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_61_bits_data, // @[:@6.4]
  input         io_dat_actv_62_valid, // @[:@6.4]
  input         io_dat_actv_62_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_62_bits_data, // @[:@6.4]
  input         io_dat_actv_63_valid, // @[:@6.4]
  input         io_dat_actv_63_bits_nz, // @[:@6.4]
  input  [7:0]  io_dat_actv_63_bits_data, // @[:@6.4]
  input         io_wt_actv_0_valid, // @[:@6.4]
  input         io_wt_actv_0_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_0_bits_data, // @[:@6.4]
  input         io_wt_actv_1_valid, // @[:@6.4]
  input         io_wt_actv_1_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_1_bits_data, // @[:@6.4]
  input         io_wt_actv_2_valid, // @[:@6.4]
  input         io_wt_actv_2_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_2_bits_data, // @[:@6.4]
  input         io_wt_actv_3_valid, // @[:@6.4]
  input         io_wt_actv_3_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_3_bits_data, // @[:@6.4]
  input         io_wt_actv_4_valid, // @[:@6.4]
  input         io_wt_actv_4_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_4_bits_data, // @[:@6.4]
  input         io_wt_actv_5_valid, // @[:@6.4]
  input         io_wt_actv_5_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_5_bits_data, // @[:@6.4]
  input         io_wt_actv_6_valid, // @[:@6.4]
  input         io_wt_actv_6_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_6_bits_data, // @[:@6.4]
  input         io_wt_actv_7_valid, // @[:@6.4]
  input         io_wt_actv_7_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_7_bits_data, // @[:@6.4]
  input         io_wt_actv_8_valid, // @[:@6.4]
  input         io_wt_actv_8_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_8_bits_data, // @[:@6.4]
  input         io_wt_actv_9_valid, // @[:@6.4]
  input         io_wt_actv_9_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_9_bits_data, // @[:@6.4]
  input         io_wt_actv_10_valid, // @[:@6.4]
  input         io_wt_actv_10_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_10_bits_data, // @[:@6.4]
  input         io_wt_actv_11_valid, // @[:@6.4]
  input         io_wt_actv_11_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_11_bits_data, // @[:@6.4]
  input         io_wt_actv_12_valid, // @[:@6.4]
  input         io_wt_actv_12_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_12_bits_data, // @[:@6.4]
  input         io_wt_actv_13_valid, // @[:@6.4]
  input         io_wt_actv_13_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_13_bits_data, // @[:@6.4]
  input         io_wt_actv_14_valid, // @[:@6.4]
  input         io_wt_actv_14_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_14_bits_data, // @[:@6.4]
  input         io_wt_actv_15_valid, // @[:@6.4]
  input         io_wt_actv_15_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_15_bits_data, // @[:@6.4]
  input         io_wt_actv_16_valid, // @[:@6.4]
  input         io_wt_actv_16_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_16_bits_data, // @[:@6.4]
  input         io_wt_actv_17_valid, // @[:@6.4]
  input         io_wt_actv_17_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_17_bits_data, // @[:@6.4]
  input         io_wt_actv_18_valid, // @[:@6.4]
  input         io_wt_actv_18_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_18_bits_data, // @[:@6.4]
  input         io_wt_actv_19_valid, // @[:@6.4]
  input         io_wt_actv_19_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_19_bits_data, // @[:@6.4]
  input         io_wt_actv_20_valid, // @[:@6.4]
  input         io_wt_actv_20_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_20_bits_data, // @[:@6.4]
  input         io_wt_actv_21_valid, // @[:@6.4]
  input         io_wt_actv_21_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_21_bits_data, // @[:@6.4]
  input         io_wt_actv_22_valid, // @[:@6.4]
  input         io_wt_actv_22_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_22_bits_data, // @[:@6.4]
  input         io_wt_actv_23_valid, // @[:@6.4]
  input         io_wt_actv_23_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_23_bits_data, // @[:@6.4]
  input         io_wt_actv_24_valid, // @[:@6.4]
  input         io_wt_actv_24_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_24_bits_data, // @[:@6.4]
  input         io_wt_actv_25_valid, // @[:@6.4]
  input         io_wt_actv_25_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_25_bits_data, // @[:@6.4]
  input         io_wt_actv_26_valid, // @[:@6.4]
  input         io_wt_actv_26_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_26_bits_data, // @[:@6.4]
  input         io_wt_actv_27_valid, // @[:@6.4]
  input         io_wt_actv_27_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_27_bits_data, // @[:@6.4]
  input         io_wt_actv_28_valid, // @[:@6.4]
  input         io_wt_actv_28_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_28_bits_data, // @[:@6.4]
  input         io_wt_actv_29_valid, // @[:@6.4]
  input         io_wt_actv_29_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_29_bits_data, // @[:@6.4]
  input         io_wt_actv_30_valid, // @[:@6.4]
  input         io_wt_actv_30_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_30_bits_data, // @[:@6.4]
  input         io_wt_actv_31_valid, // @[:@6.4]
  input         io_wt_actv_31_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_31_bits_data, // @[:@6.4]
  input         io_wt_actv_32_valid, // @[:@6.4]
  input         io_wt_actv_32_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_32_bits_data, // @[:@6.4]
  input         io_wt_actv_33_valid, // @[:@6.4]
  input         io_wt_actv_33_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_33_bits_data, // @[:@6.4]
  input         io_wt_actv_34_valid, // @[:@6.4]
  input         io_wt_actv_34_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_34_bits_data, // @[:@6.4]
  input         io_wt_actv_35_valid, // @[:@6.4]
  input         io_wt_actv_35_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_35_bits_data, // @[:@6.4]
  input         io_wt_actv_36_valid, // @[:@6.4]
  input         io_wt_actv_36_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_36_bits_data, // @[:@6.4]
  input         io_wt_actv_37_valid, // @[:@6.4]
  input         io_wt_actv_37_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_37_bits_data, // @[:@6.4]
  input         io_wt_actv_38_valid, // @[:@6.4]
  input         io_wt_actv_38_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_38_bits_data, // @[:@6.4]
  input         io_wt_actv_39_valid, // @[:@6.4]
  input         io_wt_actv_39_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_39_bits_data, // @[:@6.4]
  input         io_wt_actv_40_valid, // @[:@6.4]
  input         io_wt_actv_40_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_40_bits_data, // @[:@6.4]
  input         io_wt_actv_41_valid, // @[:@6.4]
  input         io_wt_actv_41_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_41_bits_data, // @[:@6.4]
  input         io_wt_actv_42_valid, // @[:@6.4]
  input         io_wt_actv_42_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_42_bits_data, // @[:@6.4]
  input         io_wt_actv_43_valid, // @[:@6.4]
  input         io_wt_actv_43_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_43_bits_data, // @[:@6.4]
  input         io_wt_actv_44_valid, // @[:@6.4]
  input         io_wt_actv_44_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_44_bits_data, // @[:@6.4]
  input         io_wt_actv_45_valid, // @[:@6.4]
  input         io_wt_actv_45_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_45_bits_data, // @[:@6.4]
  input         io_wt_actv_46_valid, // @[:@6.4]
  input         io_wt_actv_46_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_46_bits_data, // @[:@6.4]
  input         io_wt_actv_47_valid, // @[:@6.4]
  input         io_wt_actv_47_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_47_bits_data, // @[:@6.4]
  input         io_wt_actv_48_valid, // @[:@6.4]
  input         io_wt_actv_48_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_48_bits_data, // @[:@6.4]
  input         io_wt_actv_49_valid, // @[:@6.4]
  input         io_wt_actv_49_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_49_bits_data, // @[:@6.4]
  input         io_wt_actv_50_valid, // @[:@6.4]
  input         io_wt_actv_50_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_50_bits_data, // @[:@6.4]
  input         io_wt_actv_51_valid, // @[:@6.4]
  input         io_wt_actv_51_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_51_bits_data, // @[:@6.4]
  input         io_wt_actv_52_valid, // @[:@6.4]
  input         io_wt_actv_52_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_52_bits_data, // @[:@6.4]
  input         io_wt_actv_53_valid, // @[:@6.4]
  input         io_wt_actv_53_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_53_bits_data, // @[:@6.4]
  input         io_wt_actv_54_valid, // @[:@6.4]
  input         io_wt_actv_54_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_54_bits_data, // @[:@6.4]
  input         io_wt_actv_55_valid, // @[:@6.4]
  input         io_wt_actv_55_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_55_bits_data, // @[:@6.4]
  input         io_wt_actv_56_valid, // @[:@6.4]
  input         io_wt_actv_56_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_56_bits_data, // @[:@6.4]
  input         io_wt_actv_57_valid, // @[:@6.4]
  input         io_wt_actv_57_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_57_bits_data, // @[:@6.4]
  input         io_wt_actv_58_valid, // @[:@6.4]
  input         io_wt_actv_58_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_58_bits_data, // @[:@6.4]
  input         io_wt_actv_59_valid, // @[:@6.4]
  input         io_wt_actv_59_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_59_bits_data, // @[:@6.4]
  input         io_wt_actv_60_valid, // @[:@6.4]
  input         io_wt_actv_60_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_60_bits_data, // @[:@6.4]
  input         io_wt_actv_61_valid, // @[:@6.4]
  input         io_wt_actv_61_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_61_bits_data, // @[:@6.4]
  input         io_wt_actv_62_valid, // @[:@6.4]
  input         io_wt_actv_62_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_62_bits_data, // @[:@6.4]
  input         io_wt_actv_63_valid, // @[:@6.4]
  input         io_wt_actv_63_bits_nz, // @[:@6.4]
  input  [7:0]  io_wt_actv_63_bits_data, // @[:@6.4]
  output        io_mac_out_valid, // @[:@6.4]
  output [21:0] io_mac_out_bits // @[:@6.4]
);
  wire  _T_977; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@74.4]
  wire  _T_978; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@75.4]
  wire  _T_979; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@76.4]
  wire [7:0] _T_980; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@78.6]
  wire [7:0] _T_981; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@79.6]
  wire [15:0] _T_982; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@80.6]
  wire [15:0] _GEN_0; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@77.4]
  wire  _T_983; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@83.4]
  wire  _T_984; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@84.4]
  wire  _T_985; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@85.4]
  wire [7:0] _T_986; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@87.6]
  wire [7:0] _T_987; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@88.6]
  wire [15:0] _T_988; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@89.6]
  wire [15:0] _GEN_1; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@86.4]
  wire  _T_989; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@92.4]
  wire  _T_990; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@93.4]
  wire  _T_991; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@94.4]
  wire [7:0] _T_992; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@96.6]
  wire [7:0] _T_993; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@97.6]
  wire [15:0] _T_994; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@98.6]
  wire [15:0] _GEN_2; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@95.4]
  wire  _T_995; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@101.4]
  wire  _T_996; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@102.4]
  wire  _T_997; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@103.4]
  wire [7:0] _T_998; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@105.6]
  wire [7:0] _T_999; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@106.6]
  wire [15:0] _T_1000; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@107.6]
  wire [15:0] _GEN_3; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@104.4]
  wire  _T_1001; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@110.4]
  wire  _T_1002; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@111.4]
  wire  _T_1003; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@112.4]
  wire [7:0] _T_1004; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@114.6]
  wire [7:0] _T_1005; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@115.6]
  wire [15:0] _T_1006; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@116.6]
  wire [15:0] _GEN_4; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@113.4]
  wire  _T_1007; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@119.4]
  wire  _T_1008; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@120.4]
  wire  _T_1009; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@121.4]
  wire [7:0] _T_1010; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@123.6]
  wire [7:0] _T_1011; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@124.6]
  wire [15:0] _T_1012; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@125.6]
  wire [15:0] _GEN_5; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@122.4]
  wire  _T_1013; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@128.4]
  wire  _T_1014; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@129.4]
  wire  _T_1015; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@130.4]
  wire [7:0] _T_1016; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@132.6]
  wire [7:0] _T_1017; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@133.6]
  wire [15:0] _T_1018; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@134.6]
  wire [15:0] _GEN_6; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@131.4]
  wire  _T_1019; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@137.4]
  wire  _T_1020; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@138.4]
  wire  _T_1021; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@139.4]
  wire [7:0] _T_1022; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@141.6]
  wire [7:0] _T_1023; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@142.6]
  wire [15:0] _T_1024; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@143.6]
  wire [15:0] _GEN_7; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@140.4]
  wire  _T_1025; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@146.4]
  wire  _T_1026; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@147.4]
  wire  _T_1027; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@148.4]
  wire [7:0] _T_1028; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@150.6]
  wire [7:0] _T_1029; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@151.6]
  wire [15:0] _T_1030; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@152.6]
  wire [15:0] _GEN_8; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@149.4]
  wire  _T_1031; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@155.4]
  wire  _T_1032; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@156.4]
  wire  _T_1033; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@157.4]
  wire [7:0] _T_1034; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@159.6]
  wire [7:0] _T_1035; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@160.6]
  wire [15:0] _T_1036; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@161.6]
  wire [15:0] _GEN_9; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@158.4]
  wire  _T_1037; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@164.4]
  wire  _T_1038; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@165.4]
  wire  _T_1039; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@166.4]
  wire [7:0] _T_1040; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@168.6]
  wire [7:0] _T_1041; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@169.6]
  wire [15:0] _T_1042; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@170.6]
  wire [15:0] _GEN_10; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@167.4]
  wire  _T_1043; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@173.4]
  wire  _T_1044; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@174.4]
  wire  _T_1045; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@175.4]
  wire [7:0] _T_1046; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@177.6]
  wire [7:0] _T_1047; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@178.6]
  wire [15:0] _T_1048; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@179.6]
  wire [15:0] _GEN_11; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@176.4]
  wire  _T_1049; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@182.4]
  wire  _T_1050; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@183.4]
  wire  _T_1051; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@184.4]
  wire [7:0] _T_1052; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@186.6]
  wire [7:0] _T_1053; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@187.6]
  wire [15:0] _T_1054; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@188.6]
  wire [15:0] _GEN_12; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@185.4]
  wire  _T_1055; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@191.4]
  wire  _T_1056; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@192.4]
  wire  _T_1057; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@193.4]
  wire [7:0] _T_1058; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@195.6]
  wire [7:0] _T_1059; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@196.6]
  wire [15:0] _T_1060; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@197.6]
  wire [15:0] _GEN_13; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@194.4]
  wire  _T_1061; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@200.4]
  wire  _T_1062; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@201.4]
  wire  _T_1063; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@202.4]
  wire [7:0] _T_1064; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@204.6]
  wire [7:0] _T_1065; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@205.6]
  wire [15:0] _T_1066; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@206.6]
  wire [15:0] _GEN_14; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@203.4]
  wire  _T_1067; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@209.4]
  wire  _T_1068; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@210.4]
  wire  _T_1069; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@211.4]
  wire [7:0] _T_1070; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@213.6]
  wire [7:0] _T_1071; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@214.6]
  wire [15:0] _T_1072; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@215.6]
  wire [15:0] _GEN_15; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@212.4]
  wire  _T_1073; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@218.4]
  wire  _T_1074; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@219.4]
  wire  _T_1075; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@220.4]
  wire [7:0] _T_1076; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@222.6]
  wire [7:0] _T_1077; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@223.6]
  wire [15:0] _T_1078; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@224.6]
  wire [15:0] _GEN_16; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@221.4]
  wire  _T_1079; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@227.4]
  wire  _T_1080; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@228.4]
  wire  _T_1081; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@229.4]
  wire [7:0] _T_1082; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@231.6]
  wire [7:0] _T_1083; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@232.6]
  wire [15:0] _T_1084; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@233.6]
  wire [15:0] _GEN_17; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@230.4]
  wire  _T_1085; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@236.4]
  wire  _T_1086; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@237.4]
  wire  _T_1087; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@238.4]
  wire [7:0] _T_1088; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@240.6]
  wire [7:0] _T_1089; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@241.6]
  wire [15:0] _T_1090; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@242.6]
  wire [15:0] _GEN_18; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@239.4]
  wire  _T_1091; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@245.4]
  wire  _T_1092; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@246.4]
  wire  _T_1093; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@247.4]
  wire [7:0] _T_1094; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@249.6]
  wire [7:0] _T_1095; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@250.6]
  wire [15:0] _T_1096; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@251.6]
  wire [15:0] _GEN_19; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@248.4]
  wire  _T_1097; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@254.4]
  wire  _T_1098; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@255.4]
  wire  _T_1099; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@256.4]
  wire [7:0] _T_1100; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@258.6]
  wire [7:0] _T_1101; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@259.6]
  wire [15:0] _T_1102; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@260.6]
  wire [15:0] _GEN_20; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@257.4]
  wire  _T_1103; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@263.4]
  wire  _T_1104; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@264.4]
  wire  _T_1105; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@265.4]
  wire [7:0] _T_1106; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@267.6]
  wire [7:0] _T_1107; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@268.6]
  wire [15:0] _T_1108; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@269.6]
  wire [15:0] _GEN_21; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@266.4]
  wire  _T_1109; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@272.4]
  wire  _T_1110; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@273.4]
  wire  _T_1111; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@274.4]
  wire [7:0] _T_1112; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@276.6]
  wire [7:0] _T_1113; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@277.6]
  wire [15:0] _T_1114; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@278.6]
  wire [15:0] _GEN_22; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@275.4]
  wire  _T_1115; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@281.4]
  wire  _T_1116; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@282.4]
  wire  _T_1117; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@283.4]
  wire [7:0] _T_1118; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@285.6]
  wire [7:0] _T_1119; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@286.6]
  wire [15:0] _T_1120; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@287.6]
  wire [15:0] _GEN_23; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@284.4]
  wire  _T_1121; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@290.4]
  wire  _T_1122; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@291.4]
  wire  _T_1123; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@292.4]
  wire [7:0] _T_1124; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@294.6]
  wire [7:0] _T_1125; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@295.6]
  wire [15:0] _T_1126; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@296.6]
  wire [15:0] _GEN_24; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@293.4]
  wire  _T_1127; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@299.4]
  wire  _T_1128; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@300.4]
  wire  _T_1129; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@301.4]
  wire [7:0] _T_1130; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@303.6]
  wire [7:0] _T_1131; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@304.6]
  wire [15:0] _T_1132; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@305.6]
  wire [15:0] _GEN_25; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@302.4]
  wire  _T_1133; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@308.4]
  wire  _T_1134; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@309.4]
  wire  _T_1135; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@310.4]
  wire [7:0] _T_1136; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@312.6]
  wire [7:0] _T_1137; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@313.6]
  wire [15:0] _T_1138; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@314.6]
  wire [15:0] _GEN_26; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@311.4]
  wire  _T_1139; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@317.4]
  wire  _T_1140; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@318.4]
  wire  _T_1141; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@319.4]
  wire [7:0] _T_1142; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@321.6]
  wire [7:0] _T_1143; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@322.6]
  wire [15:0] _T_1144; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@323.6]
  wire [15:0] _GEN_27; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@320.4]
  wire  _T_1145; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@326.4]
  wire  _T_1146; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@327.4]
  wire  _T_1147; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@328.4]
  wire [7:0] _T_1148; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@330.6]
  wire [7:0] _T_1149; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@331.6]
  wire [15:0] _T_1150; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@332.6]
  wire [15:0] _GEN_28; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@329.4]
  wire  _T_1151; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@335.4]
  wire  _T_1152; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@336.4]
  wire  _T_1153; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@337.4]
  wire [7:0] _T_1154; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@339.6]
  wire [7:0] _T_1155; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@340.6]
  wire [15:0] _T_1156; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@341.6]
  wire [15:0] _GEN_29; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@338.4]
  wire  _T_1157; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@344.4]
  wire  _T_1158; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@345.4]
  wire  _T_1159; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@346.4]
  wire [7:0] _T_1160; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@348.6]
  wire [7:0] _T_1161; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@349.6]
  wire [15:0] _T_1162; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@350.6]
  wire [15:0] _GEN_30; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@347.4]
  wire  _T_1163; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@353.4]
  wire  _T_1164; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@354.4]
  wire  _T_1165; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@355.4]
  wire [7:0] _T_1166; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@357.6]
  wire [7:0] _T_1167; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@358.6]
  wire [15:0] _T_1168; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@359.6]
  wire [15:0] _GEN_31; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@356.4]
  wire  _T_1169; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@362.4]
  wire  _T_1170; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@363.4]
  wire  _T_1171; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@364.4]
  wire [7:0] _T_1172; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@366.6]
  wire [7:0] _T_1173; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@367.6]
  wire [15:0] _T_1174; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@368.6]
  wire [15:0] _GEN_32; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@365.4]
  wire  _T_1175; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@371.4]
  wire  _T_1176; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@372.4]
  wire  _T_1177; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@373.4]
  wire [7:0] _T_1178; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@375.6]
  wire [7:0] _T_1179; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@376.6]
  wire [15:0] _T_1180; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@377.6]
  wire [15:0] _GEN_33; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@374.4]
  wire  _T_1181; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@380.4]
  wire  _T_1182; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@381.4]
  wire  _T_1183; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@382.4]
  wire [7:0] _T_1184; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@384.6]
  wire [7:0] _T_1185; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@385.6]
  wire [15:0] _T_1186; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@386.6]
  wire [15:0] _GEN_34; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@383.4]
  wire  _T_1187; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@389.4]
  wire  _T_1188; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@390.4]
  wire  _T_1189; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@391.4]
  wire [7:0] _T_1190; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@393.6]
  wire [7:0] _T_1191; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@394.6]
  wire [15:0] _T_1192; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@395.6]
  wire [15:0] _GEN_35; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@392.4]
  wire  _T_1193; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@398.4]
  wire  _T_1194; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@399.4]
  wire  _T_1195; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@400.4]
  wire [7:0] _T_1196; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@402.6]
  wire [7:0] _T_1197; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@403.6]
  wire [15:0] _T_1198; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@404.6]
  wire [15:0] _GEN_36; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@401.4]
  wire  _T_1199; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@407.4]
  wire  _T_1200; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@408.4]
  wire  _T_1201; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@409.4]
  wire [7:0] _T_1202; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@411.6]
  wire [7:0] _T_1203; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@412.6]
  wire [15:0] _T_1204; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@413.6]
  wire [15:0] _GEN_37; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@410.4]
  wire  _T_1205; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@416.4]
  wire  _T_1206; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@417.4]
  wire  _T_1207; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@418.4]
  wire [7:0] _T_1208; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@420.6]
  wire [7:0] _T_1209; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@421.6]
  wire [15:0] _T_1210; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@422.6]
  wire [15:0] _GEN_38; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@419.4]
  wire  _T_1211; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@425.4]
  wire  _T_1212; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@426.4]
  wire  _T_1213; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@427.4]
  wire [7:0] _T_1214; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@429.6]
  wire [7:0] _T_1215; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@430.6]
  wire [15:0] _T_1216; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@431.6]
  wire [15:0] _GEN_39; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@428.4]
  wire  _T_1217; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@434.4]
  wire  _T_1218; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@435.4]
  wire  _T_1219; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@436.4]
  wire [7:0] _T_1220; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@438.6]
  wire [7:0] _T_1221; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@439.6]
  wire [15:0] _T_1222; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@440.6]
  wire [15:0] _GEN_40; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@437.4]
  wire  _T_1223; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@443.4]
  wire  _T_1224; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@444.4]
  wire  _T_1225; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@445.4]
  wire [7:0] _T_1226; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@447.6]
  wire [7:0] _T_1227; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@448.6]
  wire [15:0] _T_1228; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@449.6]
  wire [15:0] _GEN_41; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@446.4]
  wire  _T_1229; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@452.4]
  wire  _T_1230; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@453.4]
  wire  _T_1231; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@454.4]
  wire [7:0] _T_1232; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@456.6]
  wire [7:0] _T_1233; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@457.6]
  wire [15:0] _T_1234; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@458.6]
  wire [15:0] _GEN_42; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@455.4]
  wire  _T_1235; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@461.4]
  wire  _T_1236; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@462.4]
  wire  _T_1237; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@463.4]
  wire [7:0] _T_1238; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@465.6]
  wire [7:0] _T_1239; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@466.6]
  wire [15:0] _T_1240; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@467.6]
  wire [15:0] _GEN_43; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@464.4]
  wire  _T_1241; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@470.4]
  wire  _T_1242; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@471.4]
  wire  _T_1243; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@472.4]
  wire [7:0] _T_1244; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@474.6]
  wire [7:0] _T_1245; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@475.6]
  wire [15:0] _T_1246; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@476.6]
  wire [15:0] _GEN_44; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@473.4]
  wire  _T_1247; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@479.4]
  wire  _T_1248; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@480.4]
  wire  _T_1249; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@481.4]
  wire [7:0] _T_1250; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@483.6]
  wire [7:0] _T_1251; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@484.6]
  wire [15:0] _T_1252; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@485.6]
  wire [15:0] _GEN_45; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@482.4]
  wire  _T_1253; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@488.4]
  wire  _T_1254; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@489.4]
  wire  _T_1255; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@490.4]
  wire [7:0] _T_1256; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@492.6]
  wire [7:0] _T_1257; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@493.6]
  wire [15:0] _T_1258; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@494.6]
  wire [15:0] _GEN_46; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@491.4]
  wire  _T_1259; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@497.4]
  wire  _T_1260; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@498.4]
  wire  _T_1261; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@499.4]
  wire [7:0] _T_1262; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@501.6]
  wire [7:0] _T_1263; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@502.6]
  wire [15:0] _T_1264; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@503.6]
  wire [15:0] _GEN_47; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@500.4]
  wire  _T_1265; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@506.4]
  wire  _T_1266; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@507.4]
  wire  _T_1267; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@508.4]
  wire [7:0] _T_1268; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@510.6]
  wire [7:0] _T_1269; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@511.6]
  wire [15:0] _T_1270; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@512.6]
  wire [15:0] _GEN_48; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@509.4]
  wire  _T_1271; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@515.4]
  wire  _T_1272; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@516.4]
  wire  _T_1273; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@517.4]
  wire [7:0] _T_1274; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@519.6]
  wire [7:0] _T_1275; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@520.6]
  wire [15:0] _T_1276; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@521.6]
  wire [15:0] _GEN_49; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@518.4]
  wire  _T_1277; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@524.4]
  wire  _T_1278; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@525.4]
  wire  _T_1279; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@526.4]
  wire [7:0] _T_1280; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@528.6]
  wire [7:0] _T_1281; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@529.6]
  wire [15:0] _T_1282; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@530.6]
  wire [15:0] _GEN_50; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@527.4]
  wire  _T_1283; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@533.4]
  wire  _T_1284; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@534.4]
  wire  _T_1285; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@535.4]
  wire [7:0] _T_1286; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@537.6]
  wire [7:0] _T_1287; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@538.6]
  wire [15:0] _T_1288; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@539.6]
  wire [15:0] _GEN_51; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@536.4]
  wire  _T_1289; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@542.4]
  wire  _T_1290; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@543.4]
  wire  _T_1291; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@544.4]
  wire [7:0] _T_1292; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@546.6]
  wire [7:0] _T_1293; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@547.6]
  wire [15:0] _T_1294; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@548.6]
  wire [15:0] _GEN_52; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@545.4]
  wire  _T_1295; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@551.4]
  wire  _T_1296; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@552.4]
  wire  _T_1297; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@553.4]
  wire [7:0] _T_1298; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@555.6]
  wire [7:0] _T_1299; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@556.6]
  wire [15:0] _T_1300; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@557.6]
  wire [15:0] _GEN_53; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@554.4]
  wire  _T_1301; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@560.4]
  wire  _T_1302; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@561.4]
  wire  _T_1303; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@562.4]
  wire [7:0] _T_1304; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@564.6]
  wire [7:0] _T_1305; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@565.6]
  wire [15:0] _T_1306; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@566.6]
  wire [15:0] _GEN_54; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@563.4]
  wire  _T_1307; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@569.4]
  wire  _T_1308; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@570.4]
  wire  _T_1309; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@571.4]
  wire [7:0] _T_1310; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@573.6]
  wire [7:0] _T_1311; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@574.6]
  wire [15:0] _T_1312; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@575.6]
  wire [15:0] _GEN_55; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@572.4]
  wire  _T_1313; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@578.4]
  wire  _T_1314; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@579.4]
  wire  _T_1315; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@580.4]
  wire [7:0] _T_1316; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@582.6]
  wire [7:0] _T_1317; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@583.6]
  wire [15:0] _T_1318; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@584.6]
  wire [15:0] _GEN_56; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@581.4]
  wire  _T_1319; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@587.4]
  wire  _T_1320; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@588.4]
  wire  _T_1321; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@589.4]
  wire [7:0] _T_1322; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@591.6]
  wire [7:0] _T_1323; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@592.6]
  wire [15:0] _T_1324; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@593.6]
  wire [15:0] _GEN_57; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@590.4]
  wire  _T_1325; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@596.4]
  wire  _T_1326; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@597.4]
  wire  _T_1327; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@598.4]
  wire [7:0] _T_1328; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@600.6]
  wire [7:0] _T_1329; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@601.6]
  wire [15:0] _T_1330; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@602.6]
  wire [15:0] _GEN_58; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@599.4]
  wire  _T_1331; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@605.4]
  wire  _T_1332; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@606.4]
  wire  _T_1333; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@607.4]
  wire [7:0] _T_1334; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@609.6]
  wire [7:0] _T_1335; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@610.6]
  wire [15:0] _T_1336; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@611.6]
  wire [15:0] _GEN_59; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@608.4]
  wire  _T_1337; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@614.4]
  wire  _T_1338; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@615.4]
  wire  _T_1339; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@616.4]
  wire [7:0] _T_1340; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@618.6]
  wire [7:0] _T_1341; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@619.6]
  wire [15:0] _T_1342; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@620.6]
  wire [15:0] _GEN_60; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@617.4]
  wire  _T_1343; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@623.4]
  wire  _T_1344; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@624.4]
  wire  _T_1345; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@625.4]
  wire [7:0] _T_1346; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@627.6]
  wire [7:0] _T_1347; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@628.6]
  wire [15:0] _T_1348; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@629.6]
  wire [15:0] _GEN_61; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@626.4]
  wire  _T_1349; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@632.4]
  wire  _T_1350; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@633.4]
  wire  _T_1351; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@634.4]
  wire [7:0] _T_1352; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@636.6]
  wire [7:0] _T_1353; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@637.6]
  wire [15:0] _T_1354; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@638.6]
  wire [15:0] _GEN_62; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@635.4]
  wire  _T_1355; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@641.4]
  wire  _T_1356; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@642.4]
  wire  _T_1357; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@643.4]
  wire [7:0] _T_1358; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@645.6]
  wire [7:0] _T_1359; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@646.6]
  wire [15:0] _T_1360; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@647.6]
  wire [15:0] _GEN_63; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@644.4]
  wire [16:0] _T_1361; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@650.4]
  wire [16:0] _GEN_70; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@651.4]
  wire [17:0] _T_1362; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@651.4]
  wire [17:0] _GEN_71; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@652.4]
  wire [18:0] _T_1363; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@652.4]
  wire [18:0] _GEN_72; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@653.4]
  wire [19:0] _T_1364; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@653.4]
  wire [19:0] _GEN_73; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@654.4]
  wire [20:0] _T_1365; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@654.4]
  wire [20:0] _GEN_74; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@655.4]
  wire [21:0] _T_1366; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@655.4]
  wire [21:0] _GEN_75; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@656.4]
  wire [22:0] _T_1367; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@656.4]
  wire [22:0] _GEN_76; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@657.4]
  wire [23:0] _T_1368; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@657.4]
  wire [23:0] _GEN_77; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@658.4]
  wire [24:0] _T_1369; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@658.4]
  wire [24:0] _GEN_78; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@659.4]
  wire [25:0] _T_1370; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@659.4]
  wire [25:0] _GEN_79; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@660.4]
  wire [26:0] _T_1371; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@660.4]
  wire [26:0] _GEN_80; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@661.4]
  wire [27:0] _T_1372; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@661.4]
  wire [27:0] _GEN_81; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@662.4]
  wire [28:0] _T_1373; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@662.4]
  wire [28:0] _GEN_82; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@663.4]
  wire [29:0] _T_1374; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@663.4]
  wire [29:0] _GEN_83; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@664.4]
  wire [30:0] _T_1375; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@664.4]
  wire [30:0] _GEN_84; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@665.4]
  wire [31:0] _T_1376; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@665.4]
  wire [31:0] _GEN_85; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@666.4]
  wire [32:0] _T_1377; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@666.4]
  wire [32:0] _GEN_86; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@667.4]
  wire [33:0] _T_1378; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@667.4]
  wire [33:0] _GEN_87; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@668.4]
  wire [34:0] _T_1379; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@668.4]
  wire [34:0] _GEN_88; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@669.4]
  wire [35:0] _T_1380; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@669.4]
  wire [35:0] _GEN_89; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@670.4]
  wire [36:0] _T_1381; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@670.4]
  wire [36:0] _GEN_90; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@671.4]
  wire [37:0] _T_1382; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@671.4]
  wire [37:0] _GEN_91; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@672.4]
  wire [38:0] _T_1383; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@672.4]
  wire [38:0] _GEN_92; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@673.4]
  wire [39:0] _T_1384; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@673.4]
  wire [39:0] _GEN_93; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@674.4]
  wire [40:0] _T_1385; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@674.4]
  wire [40:0] _GEN_94; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@675.4]
  wire [41:0] _T_1386; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@675.4]
  wire [41:0] _GEN_95; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@676.4]
  wire [42:0] _T_1387; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@676.4]
  wire [42:0] _GEN_96; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@677.4]
  wire [43:0] _T_1388; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@677.4]
  wire [43:0] _GEN_97; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@678.4]
  wire [44:0] _T_1389; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@678.4]
  wire [44:0] _GEN_98; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@679.4]
  wire [45:0] _T_1390; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@679.4]
  wire [45:0] _GEN_99; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@680.4]
  wire [46:0] _T_1391; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@680.4]
  wire [46:0] _GEN_100; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@681.4]
  wire [47:0] _T_1392; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@681.4]
  wire [47:0] _GEN_101; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@682.4]
  wire [48:0] _T_1393; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@682.4]
  wire [48:0] _GEN_102; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@683.4]
  wire [49:0] _T_1394; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@683.4]
  wire [49:0] _GEN_103; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@684.4]
  wire [50:0] _T_1395; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@684.4]
  wire [50:0] _GEN_104; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@685.4]
  wire [51:0] _T_1396; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@685.4]
  wire [51:0] _GEN_105; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@686.4]
  wire [52:0] _T_1397; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@686.4]
  wire [52:0] _GEN_106; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@687.4]
  wire [53:0] _T_1398; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@687.4]
  wire [53:0] _GEN_107; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@688.4]
  wire [54:0] _T_1399; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@688.4]
  wire [54:0] _GEN_108; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@689.4]
  wire [55:0] _T_1400; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@689.4]
  wire [55:0] _GEN_109; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@690.4]
  wire [56:0] _T_1401; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@690.4]
  wire [56:0] _GEN_110; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@691.4]
  wire [57:0] _T_1402; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@691.4]
  wire [57:0] _GEN_111; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@692.4]
  wire [58:0] _T_1403; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@692.4]
  wire [58:0] _GEN_112; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@693.4]
  wire [59:0] _T_1404; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@693.4]
  wire [59:0] _GEN_113; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@694.4]
  wire [60:0] _T_1405; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@694.4]
  wire [60:0] _GEN_114; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@695.4]
  wire [61:0] _T_1406; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@695.4]
  wire [61:0] _GEN_115; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@696.4]
  wire [62:0] _T_1407; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@696.4]
  wire [62:0] _GEN_116; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@697.4]
  wire [63:0] _T_1408; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@697.4]
  wire [63:0] _GEN_117; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@698.4]
  wire [64:0] _T_1409; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@698.4]
  wire [64:0] _GEN_118; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@699.4]
  wire [65:0] _T_1410; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@699.4]
  wire [65:0] _GEN_119; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@700.4]
  wire [66:0] _T_1411; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@700.4]
  wire [66:0] _GEN_120; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@701.4]
  wire [67:0] _T_1412; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@701.4]
  wire [67:0] _GEN_121; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@702.4]
  wire [68:0] _T_1413; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@702.4]
  wire [68:0] _GEN_122; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@703.4]
  wire [69:0] _T_1414; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@703.4]
  wire [69:0] _GEN_123; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@704.4]
  wire [70:0] _T_1415; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@704.4]
  wire [70:0] _GEN_124; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@705.4]
  wire [71:0] _T_1416; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@705.4]
  wire [71:0] _GEN_125; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@706.4]
  wire [72:0] _T_1417; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@706.4]
  wire [72:0] _GEN_126; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@707.4]
  wire [73:0] _T_1418; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@707.4]
  wire [73:0] _GEN_127; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@708.4]
  wire [74:0] _T_1419; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@708.4]
  wire [74:0] _GEN_128; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@709.4]
  wire [75:0] _T_1420; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@709.4]
  wire [75:0] _GEN_129; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@710.4]
  wire [76:0] _T_1421; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@710.4]
  wire [76:0] _GEN_130; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@711.4]
  wire [77:0] _T_1422; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@711.4]
  wire [77:0] _GEN_131; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@712.4]
  wire [78:0] _T_1423; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@712.4]
  wire [78:0] _T_1424; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:37:@713.4]
  wire  _T_1425; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 59:42:@714.4]
  reg [78:0] _T_1427; // @[Reg.scala 11:16:@715.4]
  reg [95:0] _RAND_0;
  reg [78:0] _T_1429; // @[Reg.scala 11:16:@719.4]
  reg [95:0] _RAND_1;
  reg [78:0] _T_1431; // @[Reg.scala 11:16:@723.4]
  reg [95:0] _RAND_2;
  reg  _T_1433; // @[Reg.scala 11:16:@728.4]
  reg [31:0] _RAND_3;
  reg  _T_1435; // @[Reg.scala 11:16:@732.4]
  reg [31:0] _RAND_4;
  reg  _T_1437; // @[Reg.scala 11:16:@736.4]
  reg [31:0] _RAND_5;
  assign _T_977 = io_wt_actv_0_valid & io_wt_actv_0_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@74.4]
  assign _T_978 = _T_977 & io_dat_actv_0_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@75.4]
  assign _T_979 = _T_978 & io_dat_actv_0_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@76.4]
  assign _T_980 = $signed(io_wt_actv_0_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@78.6]
  assign _T_981 = $signed(io_dat_actv_0_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@79.6]
  assign _T_982 = $signed(_T_980) * $signed(_T_981); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@80.6]
  assign _GEN_0 = _T_979 ? $signed(_T_982) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@77.4]
  assign _T_983 = io_wt_actv_1_valid & io_wt_actv_1_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@83.4]
  assign _T_984 = _T_983 & io_dat_actv_1_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@84.4]
  assign _T_985 = _T_984 & io_dat_actv_1_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@85.4]
  assign _T_986 = $signed(io_wt_actv_1_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@87.6]
  assign _T_987 = $signed(io_dat_actv_1_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@88.6]
  assign _T_988 = $signed(_T_986) * $signed(_T_987); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@89.6]
  assign _GEN_1 = _T_985 ? $signed(_T_988) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@86.4]
  assign _T_989 = io_wt_actv_2_valid & io_wt_actv_2_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@92.4]
  assign _T_990 = _T_989 & io_dat_actv_2_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@93.4]
  assign _T_991 = _T_990 & io_dat_actv_2_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@94.4]
  assign _T_992 = $signed(io_wt_actv_2_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@96.6]
  assign _T_993 = $signed(io_dat_actv_2_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@97.6]
  assign _T_994 = $signed(_T_992) * $signed(_T_993); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@98.6]
  assign _GEN_2 = _T_991 ? $signed(_T_994) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@95.4]
  assign _T_995 = io_wt_actv_3_valid & io_wt_actv_3_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@101.4]
  assign _T_996 = _T_995 & io_dat_actv_3_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@102.4]
  assign _T_997 = _T_996 & io_dat_actv_3_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@103.4]
  assign _T_998 = $signed(io_wt_actv_3_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@105.6]
  assign _T_999 = $signed(io_dat_actv_3_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@106.6]
  assign _T_1000 = $signed(_T_998) * $signed(_T_999); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@107.6]
  assign _GEN_3 = _T_997 ? $signed(_T_1000) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@104.4]
  assign _T_1001 = io_wt_actv_4_valid & io_wt_actv_4_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@110.4]
  assign _T_1002 = _T_1001 & io_dat_actv_4_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@111.4]
  assign _T_1003 = _T_1002 & io_dat_actv_4_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@112.4]
  assign _T_1004 = $signed(io_wt_actv_4_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@114.6]
  assign _T_1005 = $signed(io_dat_actv_4_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@115.6]
  assign _T_1006 = $signed(_T_1004) * $signed(_T_1005); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@116.6]
  assign _GEN_4 = _T_1003 ? $signed(_T_1006) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@113.4]
  assign _T_1007 = io_wt_actv_5_valid & io_wt_actv_5_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@119.4]
  assign _T_1008 = _T_1007 & io_dat_actv_5_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@120.4]
  assign _T_1009 = _T_1008 & io_dat_actv_5_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@121.4]
  assign _T_1010 = $signed(io_wt_actv_5_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@123.6]
  assign _T_1011 = $signed(io_dat_actv_5_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@124.6]
  assign _T_1012 = $signed(_T_1010) * $signed(_T_1011); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@125.6]
  assign _GEN_5 = _T_1009 ? $signed(_T_1012) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@122.4]
  assign _T_1013 = io_wt_actv_6_valid & io_wt_actv_6_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@128.4]
  assign _T_1014 = _T_1013 & io_dat_actv_6_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@129.4]
  assign _T_1015 = _T_1014 & io_dat_actv_6_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@130.4]
  assign _T_1016 = $signed(io_wt_actv_6_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@132.6]
  assign _T_1017 = $signed(io_dat_actv_6_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@133.6]
  assign _T_1018 = $signed(_T_1016) * $signed(_T_1017); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@134.6]
  assign _GEN_6 = _T_1015 ? $signed(_T_1018) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@131.4]
  assign _T_1019 = io_wt_actv_7_valid & io_wt_actv_7_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@137.4]
  assign _T_1020 = _T_1019 & io_dat_actv_7_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@138.4]
  assign _T_1021 = _T_1020 & io_dat_actv_7_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@139.4]
  assign _T_1022 = $signed(io_wt_actv_7_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@141.6]
  assign _T_1023 = $signed(io_dat_actv_7_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@142.6]
  assign _T_1024 = $signed(_T_1022) * $signed(_T_1023); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@143.6]
  assign _GEN_7 = _T_1021 ? $signed(_T_1024) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@140.4]
  assign _T_1025 = io_wt_actv_8_valid & io_wt_actv_8_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@146.4]
  assign _T_1026 = _T_1025 & io_dat_actv_8_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@147.4]
  assign _T_1027 = _T_1026 & io_dat_actv_8_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@148.4]
  assign _T_1028 = $signed(io_wt_actv_8_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@150.6]
  assign _T_1029 = $signed(io_dat_actv_8_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@151.6]
  assign _T_1030 = $signed(_T_1028) * $signed(_T_1029); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@152.6]
  assign _GEN_8 = _T_1027 ? $signed(_T_1030) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@149.4]
  assign _T_1031 = io_wt_actv_9_valid & io_wt_actv_9_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@155.4]
  assign _T_1032 = _T_1031 & io_dat_actv_9_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@156.4]
  assign _T_1033 = _T_1032 & io_dat_actv_9_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@157.4]
  assign _T_1034 = $signed(io_wt_actv_9_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@159.6]
  assign _T_1035 = $signed(io_dat_actv_9_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@160.6]
  assign _T_1036 = $signed(_T_1034) * $signed(_T_1035); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@161.6]
  assign _GEN_9 = _T_1033 ? $signed(_T_1036) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@158.4]
  assign _T_1037 = io_wt_actv_10_valid & io_wt_actv_10_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@164.4]
  assign _T_1038 = _T_1037 & io_dat_actv_10_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@165.4]
  assign _T_1039 = _T_1038 & io_dat_actv_10_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@166.4]
  assign _T_1040 = $signed(io_wt_actv_10_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@168.6]
  assign _T_1041 = $signed(io_dat_actv_10_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@169.6]
  assign _T_1042 = $signed(_T_1040) * $signed(_T_1041); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@170.6]
  assign _GEN_10 = _T_1039 ? $signed(_T_1042) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@167.4]
  assign _T_1043 = io_wt_actv_11_valid & io_wt_actv_11_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@173.4]
  assign _T_1044 = _T_1043 & io_dat_actv_11_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@174.4]
  assign _T_1045 = _T_1044 & io_dat_actv_11_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@175.4]
  assign _T_1046 = $signed(io_wt_actv_11_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@177.6]
  assign _T_1047 = $signed(io_dat_actv_11_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@178.6]
  assign _T_1048 = $signed(_T_1046) * $signed(_T_1047); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@179.6]
  assign _GEN_11 = _T_1045 ? $signed(_T_1048) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@176.4]
  assign _T_1049 = io_wt_actv_12_valid & io_wt_actv_12_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@182.4]
  assign _T_1050 = _T_1049 & io_dat_actv_12_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@183.4]
  assign _T_1051 = _T_1050 & io_dat_actv_12_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@184.4]
  assign _T_1052 = $signed(io_wt_actv_12_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@186.6]
  assign _T_1053 = $signed(io_dat_actv_12_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@187.6]
  assign _T_1054 = $signed(_T_1052) * $signed(_T_1053); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@188.6]
  assign _GEN_12 = _T_1051 ? $signed(_T_1054) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@185.4]
  assign _T_1055 = io_wt_actv_13_valid & io_wt_actv_13_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@191.4]
  assign _T_1056 = _T_1055 & io_dat_actv_13_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@192.4]
  assign _T_1057 = _T_1056 & io_dat_actv_13_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@193.4]
  assign _T_1058 = $signed(io_wt_actv_13_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@195.6]
  assign _T_1059 = $signed(io_dat_actv_13_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@196.6]
  assign _T_1060 = $signed(_T_1058) * $signed(_T_1059); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@197.6]
  assign _GEN_13 = _T_1057 ? $signed(_T_1060) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@194.4]
  assign _T_1061 = io_wt_actv_14_valid & io_wt_actv_14_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@200.4]
  assign _T_1062 = _T_1061 & io_dat_actv_14_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@201.4]
  assign _T_1063 = _T_1062 & io_dat_actv_14_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@202.4]
  assign _T_1064 = $signed(io_wt_actv_14_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@204.6]
  assign _T_1065 = $signed(io_dat_actv_14_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@205.6]
  assign _T_1066 = $signed(_T_1064) * $signed(_T_1065); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@206.6]
  assign _GEN_14 = _T_1063 ? $signed(_T_1066) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@203.4]
  assign _T_1067 = io_wt_actv_15_valid & io_wt_actv_15_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@209.4]
  assign _T_1068 = _T_1067 & io_dat_actv_15_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@210.4]
  assign _T_1069 = _T_1068 & io_dat_actv_15_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@211.4]
  assign _T_1070 = $signed(io_wt_actv_15_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@213.6]
  assign _T_1071 = $signed(io_dat_actv_15_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@214.6]
  assign _T_1072 = $signed(_T_1070) * $signed(_T_1071); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@215.6]
  assign _GEN_15 = _T_1069 ? $signed(_T_1072) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@212.4]
  assign _T_1073 = io_wt_actv_16_valid & io_wt_actv_16_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@218.4]
  assign _T_1074 = _T_1073 & io_dat_actv_16_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@219.4]
  assign _T_1075 = _T_1074 & io_dat_actv_16_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@220.4]
  assign _T_1076 = $signed(io_wt_actv_16_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@222.6]
  assign _T_1077 = $signed(io_dat_actv_16_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@223.6]
  assign _T_1078 = $signed(_T_1076) * $signed(_T_1077); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@224.6]
  assign _GEN_16 = _T_1075 ? $signed(_T_1078) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@221.4]
  assign _T_1079 = io_wt_actv_17_valid & io_wt_actv_17_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@227.4]
  assign _T_1080 = _T_1079 & io_dat_actv_17_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@228.4]
  assign _T_1081 = _T_1080 & io_dat_actv_17_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@229.4]
  assign _T_1082 = $signed(io_wt_actv_17_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@231.6]
  assign _T_1083 = $signed(io_dat_actv_17_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@232.6]
  assign _T_1084 = $signed(_T_1082) * $signed(_T_1083); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@233.6]
  assign _GEN_17 = _T_1081 ? $signed(_T_1084) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@230.4]
  assign _T_1085 = io_wt_actv_18_valid & io_wt_actv_18_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@236.4]
  assign _T_1086 = _T_1085 & io_dat_actv_18_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@237.4]
  assign _T_1087 = _T_1086 & io_dat_actv_18_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@238.4]
  assign _T_1088 = $signed(io_wt_actv_18_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@240.6]
  assign _T_1089 = $signed(io_dat_actv_18_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@241.6]
  assign _T_1090 = $signed(_T_1088) * $signed(_T_1089); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@242.6]
  assign _GEN_18 = _T_1087 ? $signed(_T_1090) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@239.4]
  assign _T_1091 = io_wt_actv_19_valid & io_wt_actv_19_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@245.4]
  assign _T_1092 = _T_1091 & io_dat_actv_19_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@246.4]
  assign _T_1093 = _T_1092 & io_dat_actv_19_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@247.4]
  assign _T_1094 = $signed(io_wt_actv_19_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@249.6]
  assign _T_1095 = $signed(io_dat_actv_19_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@250.6]
  assign _T_1096 = $signed(_T_1094) * $signed(_T_1095); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@251.6]
  assign _GEN_19 = _T_1093 ? $signed(_T_1096) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@248.4]
  assign _T_1097 = io_wt_actv_20_valid & io_wt_actv_20_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@254.4]
  assign _T_1098 = _T_1097 & io_dat_actv_20_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@255.4]
  assign _T_1099 = _T_1098 & io_dat_actv_20_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@256.4]
  assign _T_1100 = $signed(io_wt_actv_20_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@258.6]
  assign _T_1101 = $signed(io_dat_actv_20_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@259.6]
  assign _T_1102 = $signed(_T_1100) * $signed(_T_1101); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@260.6]
  assign _GEN_20 = _T_1099 ? $signed(_T_1102) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@257.4]
  assign _T_1103 = io_wt_actv_21_valid & io_wt_actv_21_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@263.4]
  assign _T_1104 = _T_1103 & io_dat_actv_21_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@264.4]
  assign _T_1105 = _T_1104 & io_dat_actv_21_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@265.4]
  assign _T_1106 = $signed(io_wt_actv_21_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@267.6]
  assign _T_1107 = $signed(io_dat_actv_21_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@268.6]
  assign _T_1108 = $signed(_T_1106) * $signed(_T_1107); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@269.6]
  assign _GEN_21 = _T_1105 ? $signed(_T_1108) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@266.4]
  assign _T_1109 = io_wt_actv_22_valid & io_wt_actv_22_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@272.4]
  assign _T_1110 = _T_1109 & io_dat_actv_22_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@273.4]
  assign _T_1111 = _T_1110 & io_dat_actv_22_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@274.4]
  assign _T_1112 = $signed(io_wt_actv_22_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@276.6]
  assign _T_1113 = $signed(io_dat_actv_22_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@277.6]
  assign _T_1114 = $signed(_T_1112) * $signed(_T_1113); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@278.6]
  assign _GEN_22 = _T_1111 ? $signed(_T_1114) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@275.4]
  assign _T_1115 = io_wt_actv_23_valid & io_wt_actv_23_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@281.4]
  assign _T_1116 = _T_1115 & io_dat_actv_23_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@282.4]
  assign _T_1117 = _T_1116 & io_dat_actv_23_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@283.4]
  assign _T_1118 = $signed(io_wt_actv_23_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@285.6]
  assign _T_1119 = $signed(io_dat_actv_23_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@286.6]
  assign _T_1120 = $signed(_T_1118) * $signed(_T_1119); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@287.6]
  assign _GEN_23 = _T_1117 ? $signed(_T_1120) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@284.4]
  assign _T_1121 = io_wt_actv_24_valid & io_wt_actv_24_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@290.4]
  assign _T_1122 = _T_1121 & io_dat_actv_24_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@291.4]
  assign _T_1123 = _T_1122 & io_dat_actv_24_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@292.4]
  assign _T_1124 = $signed(io_wt_actv_24_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@294.6]
  assign _T_1125 = $signed(io_dat_actv_24_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@295.6]
  assign _T_1126 = $signed(_T_1124) * $signed(_T_1125); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@296.6]
  assign _GEN_24 = _T_1123 ? $signed(_T_1126) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@293.4]
  assign _T_1127 = io_wt_actv_25_valid & io_wt_actv_25_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@299.4]
  assign _T_1128 = _T_1127 & io_dat_actv_25_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@300.4]
  assign _T_1129 = _T_1128 & io_dat_actv_25_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@301.4]
  assign _T_1130 = $signed(io_wt_actv_25_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@303.6]
  assign _T_1131 = $signed(io_dat_actv_25_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@304.6]
  assign _T_1132 = $signed(_T_1130) * $signed(_T_1131); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@305.6]
  assign _GEN_25 = _T_1129 ? $signed(_T_1132) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@302.4]
  assign _T_1133 = io_wt_actv_26_valid & io_wt_actv_26_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@308.4]
  assign _T_1134 = _T_1133 & io_dat_actv_26_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@309.4]
  assign _T_1135 = _T_1134 & io_dat_actv_26_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@310.4]
  assign _T_1136 = $signed(io_wt_actv_26_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@312.6]
  assign _T_1137 = $signed(io_dat_actv_26_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@313.6]
  assign _T_1138 = $signed(_T_1136) * $signed(_T_1137); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@314.6]
  assign _GEN_26 = _T_1135 ? $signed(_T_1138) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@311.4]
  assign _T_1139 = io_wt_actv_27_valid & io_wt_actv_27_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@317.4]
  assign _T_1140 = _T_1139 & io_dat_actv_27_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@318.4]
  assign _T_1141 = _T_1140 & io_dat_actv_27_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@319.4]
  assign _T_1142 = $signed(io_wt_actv_27_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@321.6]
  assign _T_1143 = $signed(io_dat_actv_27_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@322.6]
  assign _T_1144 = $signed(_T_1142) * $signed(_T_1143); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@323.6]
  assign _GEN_27 = _T_1141 ? $signed(_T_1144) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@320.4]
  assign _T_1145 = io_wt_actv_28_valid & io_wt_actv_28_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@326.4]
  assign _T_1146 = _T_1145 & io_dat_actv_28_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@327.4]
  assign _T_1147 = _T_1146 & io_dat_actv_28_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@328.4]
  assign _T_1148 = $signed(io_wt_actv_28_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@330.6]
  assign _T_1149 = $signed(io_dat_actv_28_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@331.6]
  assign _T_1150 = $signed(_T_1148) * $signed(_T_1149); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@332.6]
  assign _GEN_28 = _T_1147 ? $signed(_T_1150) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@329.4]
  assign _T_1151 = io_wt_actv_29_valid & io_wt_actv_29_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@335.4]
  assign _T_1152 = _T_1151 & io_dat_actv_29_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@336.4]
  assign _T_1153 = _T_1152 & io_dat_actv_29_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@337.4]
  assign _T_1154 = $signed(io_wt_actv_29_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@339.6]
  assign _T_1155 = $signed(io_dat_actv_29_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@340.6]
  assign _T_1156 = $signed(_T_1154) * $signed(_T_1155); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@341.6]
  assign _GEN_29 = _T_1153 ? $signed(_T_1156) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@338.4]
  assign _T_1157 = io_wt_actv_30_valid & io_wt_actv_30_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@344.4]
  assign _T_1158 = _T_1157 & io_dat_actv_30_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@345.4]
  assign _T_1159 = _T_1158 & io_dat_actv_30_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@346.4]
  assign _T_1160 = $signed(io_wt_actv_30_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@348.6]
  assign _T_1161 = $signed(io_dat_actv_30_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@349.6]
  assign _T_1162 = $signed(_T_1160) * $signed(_T_1161); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@350.6]
  assign _GEN_30 = _T_1159 ? $signed(_T_1162) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@347.4]
  assign _T_1163 = io_wt_actv_31_valid & io_wt_actv_31_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@353.4]
  assign _T_1164 = _T_1163 & io_dat_actv_31_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@354.4]
  assign _T_1165 = _T_1164 & io_dat_actv_31_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@355.4]
  assign _T_1166 = $signed(io_wt_actv_31_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@357.6]
  assign _T_1167 = $signed(io_dat_actv_31_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@358.6]
  assign _T_1168 = $signed(_T_1166) * $signed(_T_1167); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@359.6]
  assign _GEN_31 = _T_1165 ? $signed(_T_1168) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@356.4]
  assign _T_1169 = io_wt_actv_32_valid & io_wt_actv_32_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@362.4]
  assign _T_1170 = _T_1169 & io_dat_actv_32_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@363.4]
  assign _T_1171 = _T_1170 & io_dat_actv_32_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@364.4]
  assign _T_1172 = $signed(io_wt_actv_32_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@366.6]
  assign _T_1173 = $signed(io_dat_actv_32_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@367.6]
  assign _T_1174 = $signed(_T_1172) * $signed(_T_1173); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@368.6]
  assign _GEN_32 = _T_1171 ? $signed(_T_1174) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@365.4]
  assign _T_1175 = io_wt_actv_33_valid & io_wt_actv_33_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@371.4]
  assign _T_1176 = _T_1175 & io_dat_actv_33_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@372.4]
  assign _T_1177 = _T_1176 & io_dat_actv_33_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@373.4]
  assign _T_1178 = $signed(io_wt_actv_33_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@375.6]
  assign _T_1179 = $signed(io_dat_actv_33_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@376.6]
  assign _T_1180 = $signed(_T_1178) * $signed(_T_1179); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@377.6]
  assign _GEN_33 = _T_1177 ? $signed(_T_1180) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@374.4]
  assign _T_1181 = io_wt_actv_34_valid & io_wt_actv_34_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@380.4]
  assign _T_1182 = _T_1181 & io_dat_actv_34_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@381.4]
  assign _T_1183 = _T_1182 & io_dat_actv_34_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@382.4]
  assign _T_1184 = $signed(io_wt_actv_34_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@384.6]
  assign _T_1185 = $signed(io_dat_actv_34_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@385.6]
  assign _T_1186 = $signed(_T_1184) * $signed(_T_1185); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@386.6]
  assign _GEN_34 = _T_1183 ? $signed(_T_1186) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@383.4]
  assign _T_1187 = io_wt_actv_35_valid & io_wt_actv_35_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@389.4]
  assign _T_1188 = _T_1187 & io_dat_actv_35_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@390.4]
  assign _T_1189 = _T_1188 & io_dat_actv_35_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@391.4]
  assign _T_1190 = $signed(io_wt_actv_35_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@393.6]
  assign _T_1191 = $signed(io_dat_actv_35_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@394.6]
  assign _T_1192 = $signed(_T_1190) * $signed(_T_1191); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@395.6]
  assign _GEN_35 = _T_1189 ? $signed(_T_1192) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@392.4]
  assign _T_1193 = io_wt_actv_36_valid & io_wt_actv_36_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@398.4]
  assign _T_1194 = _T_1193 & io_dat_actv_36_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@399.4]
  assign _T_1195 = _T_1194 & io_dat_actv_36_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@400.4]
  assign _T_1196 = $signed(io_wt_actv_36_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@402.6]
  assign _T_1197 = $signed(io_dat_actv_36_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@403.6]
  assign _T_1198 = $signed(_T_1196) * $signed(_T_1197); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@404.6]
  assign _GEN_36 = _T_1195 ? $signed(_T_1198) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@401.4]
  assign _T_1199 = io_wt_actv_37_valid & io_wt_actv_37_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@407.4]
  assign _T_1200 = _T_1199 & io_dat_actv_37_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@408.4]
  assign _T_1201 = _T_1200 & io_dat_actv_37_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@409.4]
  assign _T_1202 = $signed(io_wt_actv_37_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@411.6]
  assign _T_1203 = $signed(io_dat_actv_37_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@412.6]
  assign _T_1204 = $signed(_T_1202) * $signed(_T_1203); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@413.6]
  assign _GEN_37 = _T_1201 ? $signed(_T_1204) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@410.4]
  assign _T_1205 = io_wt_actv_38_valid & io_wt_actv_38_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@416.4]
  assign _T_1206 = _T_1205 & io_dat_actv_38_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@417.4]
  assign _T_1207 = _T_1206 & io_dat_actv_38_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@418.4]
  assign _T_1208 = $signed(io_wt_actv_38_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@420.6]
  assign _T_1209 = $signed(io_dat_actv_38_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@421.6]
  assign _T_1210 = $signed(_T_1208) * $signed(_T_1209); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@422.6]
  assign _GEN_38 = _T_1207 ? $signed(_T_1210) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@419.4]
  assign _T_1211 = io_wt_actv_39_valid & io_wt_actv_39_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@425.4]
  assign _T_1212 = _T_1211 & io_dat_actv_39_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@426.4]
  assign _T_1213 = _T_1212 & io_dat_actv_39_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@427.4]
  assign _T_1214 = $signed(io_wt_actv_39_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@429.6]
  assign _T_1215 = $signed(io_dat_actv_39_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@430.6]
  assign _T_1216 = $signed(_T_1214) * $signed(_T_1215); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@431.6]
  assign _GEN_39 = _T_1213 ? $signed(_T_1216) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@428.4]
  assign _T_1217 = io_wt_actv_40_valid & io_wt_actv_40_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@434.4]
  assign _T_1218 = _T_1217 & io_dat_actv_40_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@435.4]
  assign _T_1219 = _T_1218 & io_dat_actv_40_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@436.4]
  assign _T_1220 = $signed(io_wt_actv_40_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@438.6]
  assign _T_1221 = $signed(io_dat_actv_40_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@439.6]
  assign _T_1222 = $signed(_T_1220) * $signed(_T_1221); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@440.6]
  assign _GEN_40 = _T_1219 ? $signed(_T_1222) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@437.4]
  assign _T_1223 = io_wt_actv_41_valid & io_wt_actv_41_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@443.4]
  assign _T_1224 = _T_1223 & io_dat_actv_41_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@444.4]
  assign _T_1225 = _T_1224 & io_dat_actv_41_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@445.4]
  assign _T_1226 = $signed(io_wt_actv_41_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@447.6]
  assign _T_1227 = $signed(io_dat_actv_41_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@448.6]
  assign _T_1228 = $signed(_T_1226) * $signed(_T_1227); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@449.6]
  assign _GEN_41 = _T_1225 ? $signed(_T_1228) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@446.4]
  assign _T_1229 = io_wt_actv_42_valid & io_wt_actv_42_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@452.4]
  assign _T_1230 = _T_1229 & io_dat_actv_42_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@453.4]
  assign _T_1231 = _T_1230 & io_dat_actv_42_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@454.4]
  assign _T_1232 = $signed(io_wt_actv_42_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@456.6]
  assign _T_1233 = $signed(io_dat_actv_42_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@457.6]
  assign _T_1234 = $signed(_T_1232) * $signed(_T_1233); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@458.6]
  assign _GEN_42 = _T_1231 ? $signed(_T_1234) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@455.4]
  assign _T_1235 = io_wt_actv_43_valid & io_wt_actv_43_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@461.4]
  assign _T_1236 = _T_1235 & io_dat_actv_43_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@462.4]
  assign _T_1237 = _T_1236 & io_dat_actv_43_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@463.4]
  assign _T_1238 = $signed(io_wt_actv_43_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@465.6]
  assign _T_1239 = $signed(io_dat_actv_43_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@466.6]
  assign _T_1240 = $signed(_T_1238) * $signed(_T_1239); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@467.6]
  assign _GEN_43 = _T_1237 ? $signed(_T_1240) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@464.4]
  assign _T_1241 = io_wt_actv_44_valid & io_wt_actv_44_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@470.4]
  assign _T_1242 = _T_1241 & io_dat_actv_44_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@471.4]
  assign _T_1243 = _T_1242 & io_dat_actv_44_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@472.4]
  assign _T_1244 = $signed(io_wt_actv_44_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@474.6]
  assign _T_1245 = $signed(io_dat_actv_44_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@475.6]
  assign _T_1246 = $signed(_T_1244) * $signed(_T_1245); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@476.6]
  assign _GEN_44 = _T_1243 ? $signed(_T_1246) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@473.4]
  assign _T_1247 = io_wt_actv_45_valid & io_wt_actv_45_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@479.4]
  assign _T_1248 = _T_1247 & io_dat_actv_45_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@480.4]
  assign _T_1249 = _T_1248 & io_dat_actv_45_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@481.4]
  assign _T_1250 = $signed(io_wt_actv_45_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@483.6]
  assign _T_1251 = $signed(io_dat_actv_45_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@484.6]
  assign _T_1252 = $signed(_T_1250) * $signed(_T_1251); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@485.6]
  assign _GEN_45 = _T_1249 ? $signed(_T_1252) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@482.4]
  assign _T_1253 = io_wt_actv_46_valid & io_wt_actv_46_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@488.4]
  assign _T_1254 = _T_1253 & io_dat_actv_46_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@489.4]
  assign _T_1255 = _T_1254 & io_dat_actv_46_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@490.4]
  assign _T_1256 = $signed(io_wt_actv_46_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@492.6]
  assign _T_1257 = $signed(io_dat_actv_46_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@493.6]
  assign _T_1258 = $signed(_T_1256) * $signed(_T_1257); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@494.6]
  assign _GEN_46 = _T_1255 ? $signed(_T_1258) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@491.4]
  assign _T_1259 = io_wt_actv_47_valid & io_wt_actv_47_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@497.4]
  assign _T_1260 = _T_1259 & io_dat_actv_47_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@498.4]
  assign _T_1261 = _T_1260 & io_dat_actv_47_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@499.4]
  assign _T_1262 = $signed(io_wt_actv_47_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@501.6]
  assign _T_1263 = $signed(io_dat_actv_47_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@502.6]
  assign _T_1264 = $signed(_T_1262) * $signed(_T_1263); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@503.6]
  assign _GEN_47 = _T_1261 ? $signed(_T_1264) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@500.4]
  assign _T_1265 = io_wt_actv_48_valid & io_wt_actv_48_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@506.4]
  assign _T_1266 = _T_1265 & io_dat_actv_48_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@507.4]
  assign _T_1267 = _T_1266 & io_dat_actv_48_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@508.4]
  assign _T_1268 = $signed(io_wt_actv_48_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@510.6]
  assign _T_1269 = $signed(io_dat_actv_48_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@511.6]
  assign _T_1270 = $signed(_T_1268) * $signed(_T_1269); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@512.6]
  assign _GEN_48 = _T_1267 ? $signed(_T_1270) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@509.4]
  assign _T_1271 = io_wt_actv_49_valid & io_wt_actv_49_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@515.4]
  assign _T_1272 = _T_1271 & io_dat_actv_49_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@516.4]
  assign _T_1273 = _T_1272 & io_dat_actv_49_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@517.4]
  assign _T_1274 = $signed(io_wt_actv_49_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@519.6]
  assign _T_1275 = $signed(io_dat_actv_49_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@520.6]
  assign _T_1276 = $signed(_T_1274) * $signed(_T_1275); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@521.6]
  assign _GEN_49 = _T_1273 ? $signed(_T_1276) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@518.4]
  assign _T_1277 = io_wt_actv_50_valid & io_wt_actv_50_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@524.4]
  assign _T_1278 = _T_1277 & io_dat_actv_50_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@525.4]
  assign _T_1279 = _T_1278 & io_dat_actv_50_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@526.4]
  assign _T_1280 = $signed(io_wt_actv_50_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@528.6]
  assign _T_1281 = $signed(io_dat_actv_50_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@529.6]
  assign _T_1282 = $signed(_T_1280) * $signed(_T_1281); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@530.6]
  assign _GEN_50 = _T_1279 ? $signed(_T_1282) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@527.4]
  assign _T_1283 = io_wt_actv_51_valid & io_wt_actv_51_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@533.4]
  assign _T_1284 = _T_1283 & io_dat_actv_51_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@534.4]
  assign _T_1285 = _T_1284 & io_dat_actv_51_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@535.4]
  assign _T_1286 = $signed(io_wt_actv_51_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@537.6]
  assign _T_1287 = $signed(io_dat_actv_51_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@538.6]
  assign _T_1288 = $signed(_T_1286) * $signed(_T_1287); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@539.6]
  assign _GEN_51 = _T_1285 ? $signed(_T_1288) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@536.4]
  assign _T_1289 = io_wt_actv_52_valid & io_wt_actv_52_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@542.4]
  assign _T_1290 = _T_1289 & io_dat_actv_52_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@543.4]
  assign _T_1291 = _T_1290 & io_dat_actv_52_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@544.4]
  assign _T_1292 = $signed(io_wt_actv_52_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@546.6]
  assign _T_1293 = $signed(io_dat_actv_52_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@547.6]
  assign _T_1294 = $signed(_T_1292) * $signed(_T_1293); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@548.6]
  assign _GEN_52 = _T_1291 ? $signed(_T_1294) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@545.4]
  assign _T_1295 = io_wt_actv_53_valid & io_wt_actv_53_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@551.4]
  assign _T_1296 = _T_1295 & io_dat_actv_53_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@552.4]
  assign _T_1297 = _T_1296 & io_dat_actv_53_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@553.4]
  assign _T_1298 = $signed(io_wt_actv_53_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@555.6]
  assign _T_1299 = $signed(io_dat_actv_53_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@556.6]
  assign _T_1300 = $signed(_T_1298) * $signed(_T_1299); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@557.6]
  assign _GEN_53 = _T_1297 ? $signed(_T_1300) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@554.4]
  assign _T_1301 = io_wt_actv_54_valid & io_wt_actv_54_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@560.4]
  assign _T_1302 = _T_1301 & io_dat_actv_54_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@561.4]
  assign _T_1303 = _T_1302 & io_dat_actv_54_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@562.4]
  assign _T_1304 = $signed(io_wt_actv_54_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@564.6]
  assign _T_1305 = $signed(io_dat_actv_54_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@565.6]
  assign _T_1306 = $signed(_T_1304) * $signed(_T_1305); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@566.6]
  assign _GEN_54 = _T_1303 ? $signed(_T_1306) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@563.4]
  assign _T_1307 = io_wt_actv_55_valid & io_wt_actv_55_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@569.4]
  assign _T_1308 = _T_1307 & io_dat_actv_55_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@570.4]
  assign _T_1309 = _T_1308 & io_dat_actv_55_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@571.4]
  assign _T_1310 = $signed(io_wt_actv_55_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@573.6]
  assign _T_1311 = $signed(io_dat_actv_55_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@574.6]
  assign _T_1312 = $signed(_T_1310) * $signed(_T_1311); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@575.6]
  assign _GEN_55 = _T_1309 ? $signed(_T_1312) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@572.4]
  assign _T_1313 = io_wt_actv_56_valid & io_wt_actv_56_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@578.4]
  assign _T_1314 = _T_1313 & io_dat_actv_56_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@579.4]
  assign _T_1315 = _T_1314 & io_dat_actv_56_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@580.4]
  assign _T_1316 = $signed(io_wt_actv_56_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@582.6]
  assign _T_1317 = $signed(io_dat_actv_56_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@583.6]
  assign _T_1318 = $signed(_T_1316) * $signed(_T_1317); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@584.6]
  assign _GEN_56 = _T_1315 ? $signed(_T_1318) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@581.4]
  assign _T_1319 = io_wt_actv_57_valid & io_wt_actv_57_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@587.4]
  assign _T_1320 = _T_1319 & io_dat_actv_57_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@588.4]
  assign _T_1321 = _T_1320 & io_dat_actv_57_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@589.4]
  assign _T_1322 = $signed(io_wt_actv_57_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@591.6]
  assign _T_1323 = $signed(io_dat_actv_57_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@592.6]
  assign _T_1324 = $signed(_T_1322) * $signed(_T_1323); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@593.6]
  assign _GEN_57 = _T_1321 ? $signed(_T_1324) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@590.4]
  assign _T_1325 = io_wt_actv_58_valid & io_wt_actv_58_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@596.4]
  assign _T_1326 = _T_1325 & io_dat_actv_58_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@597.4]
  assign _T_1327 = _T_1326 & io_dat_actv_58_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@598.4]
  assign _T_1328 = $signed(io_wt_actv_58_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@600.6]
  assign _T_1329 = $signed(io_dat_actv_58_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@601.6]
  assign _T_1330 = $signed(_T_1328) * $signed(_T_1329); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@602.6]
  assign _GEN_58 = _T_1327 ? $signed(_T_1330) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@599.4]
  assign _T_1331 = io_wt_actv_59_valid & io_wt_actv_59_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@605.4]
  assign _T_1332 = _T_1331 & io_dat_actv_59_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@606.4]
  assign _T_1333 = _T_1332 & io_dat_actv_59_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@607.4]
  assign _T_1334 = $signed(io_wt_actv_59_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@609.6]
  assign _T_1335 = $signed(io_dat_actv_59_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@610.6]
  assign _T_1336 = $signed(_T_1334) * $signed(_T_1335); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@611.6]
  assign _GEN_59 = _T_1333 ? $signed(_T_1336) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@608.4]
  assign _T_1337 = io_wt_actv_60_valid & io_wt_actv_60_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@614.4]
  assign _T_1338 = _T_1337 & io_dat_actv_60_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@615.4]
  assign _T_1339 = _T_1338 & io_dat_actv_60_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@616.4]
  assign _T_1340 = $signed(io_wt_actv_60_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@618.6]
  assign _T_1341 = $signed(io_dat_actv_60_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@619.6]
  assign _T_1342 = $signed(_T_1340) * $signed(_T_1341); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@620.6]
  assign _GEN_60 = _T_1339 ? $signed(_T_1342) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@617.4]
  assign _T_1343 = io_wt_actv_61_valid & io_wt_actv_61_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@623.4]
  assign _T_1344 = _T_1343 & io_dat_actv_61_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@624.4]
  assign _T_1345 = _T_1344 & io_dat_actv_61_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@625.4]
  assign _T_1346 = $signed(io_wt_actv_61_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@627.6]
  assign _T_1347 = $signed(io_dat_actv_61_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@628.6]
  assign _T_1348 = $signed(_T_1346) * $signed(_T_1347); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@629.6]
  assign _GEN_61 = _T_1345 ? $signed(_T_1348) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@626.4]
  assign _T_1349 = io_wt_actv_62_valid & io_wt_actv_62_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@632.4]
  assign _T_1350 = _T_1349 & io_dat_actv_62_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@633.4]
  assign _T_1351 = _T_1350 & io_dat_actv_62_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@634.4]
  assign _T_1352 = $signed(io_wt_actv_62_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@636.6]
  assign _T_1353 = $signed(io_dat_actv_62_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@637.6]
  assign _T_1354 = $signed(_T_1352) * $signed(_T_1353); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@638.6]
  assign _GEN_62 = _T_1351 ? $signed(_T_1354) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@635.4]
  assign _T_1355 = io_wt_actv_63_valid & io_wt_actv_63_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:33:@641.4]
  assign _T_1356 = _T_1355 & io_dat_actv_63_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:55:@642.4]
  assign _T_1357 = _T_1356 & io_dat_actv_63_bits_nz; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:76:@643.4]
  assign _T_1358 = $signed(io_wt_actv_63_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:49:@645.6]
  assign _T_1359 = $signed(io_dat_actv_63_bits_data); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:81:@646.6]
  assign _T_1360 = $signed(_T_1358) * $signed(_T_1359); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 52:55:@647.6]
  assign _GEN_63 = _T_1357 ? $signed(_T_1360) : $signed(16'sh0); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 51:100:@644.4]
  assign _T_1361 = $signed(_GEN_0) + $signed(_GEN_1); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@650.4]
  assign _GEN_70 = {{1{_GEN_2[15]}},_GEN_2}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@651.4]
  assign _T_1362 = $signed(_T_1361) + $signed(_GEN_70); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@651.4]
  assign _GEN_71 = {{2{_GEN_3[15]}},_GEN_3}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@652.4]
  assign _T_1363 = $signed(_T_1362) + $signed(_GEN_71); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@652.4]
  assign _GEN_72 = {{3{_GEN_4[15]}},_GEN_4}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@653.4]
  assign _T_1364 = $signed(_T_1363) + $signed(_GEN_72); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@653.4]
  assign _GEN_73 = {{4{_GEN_5[15]}},_GEN_5}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@654.4]
  assign _T_1365 = $signed(_T_1364) + $signed(_GEN_73); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@654.4]
  assign _GEN_74 = {{5{_GEN_6[15]}},_GEN_6}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@655.4]
  assign _T_1366 = $signed(_T_1365) + $signed(_GEN_74); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@655.4]
  assign _GEN_75 = {{6{_GEN_7[15]}},_GEN_7}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@656.4]
  assign _T_1367 = $signed(_T_1366) + $signed(_GEN_75); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@656.4]
  assign _GEN_76 = {{7{_GEN_8[15]}},_GEN_8}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@657.4]
  assign _T_1368 = $signed(_T_1367) + $signed(_GEN_76); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@657.4]
  assign _GEN_77 = {{8{_GEN_9[15]}},_GEN_9}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@658.4]
  assign _T_1369 = $signed(_T_1368) + $signed(_GEN_77); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@658.4]
  assign _GEN_78 = {{9{_GEN_10[15]}},_GEN_10}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@659.4]
  assign _T_1370 = $signed(_T_1369) + $signed(_GEN_78); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@659.4]
  assign _GEN_79 = {{10{_GEN_11[15]}},_GEN_11}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@660.4]
  assign _T_1371 = $signed(_T_1370) + $signed(_GEN_79); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@660.4]
  assign _GEN_80 = {{11{_GEN_12[15]}},_GEN_12}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@661.4]
  assign _T_1372 = $signed(_T_1371) + $signed(_GEN_80); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@661.4]
  assign _GEN_81 = {{12{_GEN_13[15]}},_GEN_13}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@662.4]
  assign _T_1373 = $signed(_T_1372) + $signed(_GEN_81); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@662.4]
  assign _GEN_82 = {{13{_GEN_14[15]}},_GEN_14}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@663.4]
  assign _T_1374 = $signed(_T_1373) + $signed(_GEN_82); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@663.4]
  assign _GEN_83 = {{14{_GEN_15[15]}},_GEN_15}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@664.4]
  assign _T_1375 = $signed(_T_1374) + $signed(_GEN_83); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@664.4]
  assign _GEN_84 = {{15{_GEN_16[15]}},_GEN_16}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@665.4]
  assign _T_1376 = $signed(_T_1375) + $signed(_GEN_84); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@665.4]
  assign _GEN_85 = {{16{_GEN_17[15]}},_GEN_17}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@666.4]
  assign _T_1377 = $signed(_T_1376) + $signed(_GEN_85); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@666.4]
  assign _GEN_86 = {{17{_GEN_18[15]}},_GEN_18}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@667.4]
  assign _T_1378 = $signed(_T_1377) + $signed(_GEN_86); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@667.4]
  assign _GEN_87 = {{18{_GEN_19[15]}},_GEN_19}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@668.4]
  assign _T_1379 = $signed(_T_1378) + $signed(_GEN_87); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@668.4]
  assign _GEN_88 = {{19{_GEN_20[15]}},_GEN_20}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@669.4]
  assign _T_1380 = $signed(_T_1379) + $signed(_GEN_88); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@669.4]
  assign _GEN_89 = {{20{_GEN_21[15]}},_GEN_21}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@670.4]
  assign _T_1381 = $signed(_T_1380) + $signed(_GEN_89); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@670.4]
  assign _GEN_90 = {{21{_GEN_22[15]}},_GEN_22}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@671.4]
  assign _T_1382 = $signed(_T_1381) + $signed(_GEN_90); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@671.4]
  assign _GEN_91 = {{22{_GEN_23[15]}},_GEN_23}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@672.4]
  assign _T_1383 = $signed(_T_1382) + $signed(_GEN_91); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@672.4]
  assign _GEN_92 = {{23{_GEN_24[15]}},_GEN_24}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@673.4]
  assign _T_1384 = $signed(_T_1383) + $signed(_GEN_92); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@673.4]
  assign _GEN_93 = {{24{_GEN_25[15]}},_GEN_25}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@674.4]
  assign _T_1385 = $signed(_T_1384) + $signed(_GEN_93); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@674.4]
  assign _GEN_94 = {{25{_GEN_26[15]}},_GEN_26}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@675.4]
  assign _T_1386 = $signed(_T_1385) + $signed(_GEN_94); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@675.4]
  assign _GEN_95 = {{26{_GEN_27[15]}},_GEN_27}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@676.4]
  assign _T_1387 = $signed(_T_1386) + $signed(_GEN_95); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@676.4]
  assign _GEN_96 = {{27{_GEN_28[15]}},_GEN_28}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@677.4]
  assign _T_1388 = $signed(_T_1387) + $signed(_GEN_96); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@677.4]
  assign _GEN_97 = {{28{_GEN_29[15]}},_GEN_29}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@678.4]
  assign _T_1389 = $signed(_T_1388) + $signed(_GEN_97); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@678.4]
  assign _GEN_98 = {{29{_GEN_30[15]}},_GEN_30}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@679.4]
  assign _T_1390 = $signed(_T_1389) + $signed(_GEN_98); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@679.4]
  assign _GEN_99 = {{30{_GEN_31[15]}},_GEN_31}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@680.4]
  assign _T_1391 = $signed(_T_1390) + $signed(_GEN_99); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@680.4]
  assign _GEN_100 = {{31{_GEN_32[15]}},_GEN_32}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@681.4]
  assign _T_1392 = $signed(_T_1391) + $signed(_GEN_100); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@681.4]
  assign _GEN_101 = {{32{_GEN_33[15]}},_GEN_33}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@682.4]
  assign _T_1393 = $signed(_T_1392) + $signed(_GEN_101); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@682.4]
  assign _GEN_102 = {{33{_GEN_34[15]}},_GEN_34}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@683.4]
  assign _T_1394 = $signed(_T_1393) + $signed(_GEN_102); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@683.4]
  assign _GEN_103 = {{34{_GEN_35[15]}},_GEN_35}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@684.4]
  assign _T_1395 = $signed(_T_1394) + $signed(_GEN_103); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@684.4]
  assign _GEN_104 = {{35{_GEN_36[15]}},_GEN_36}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@685.4]
  assign _T_1396 = $signed(_T_1395) + $signed(_GEN_104); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@685.4]
  assign _GEN_105 = {{36{_GEN_37[15]}},_GEN_37}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@686.4]
  assign _T_1397 = $signed(_T_1396) + $signed(_GEN_105); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@686.4]
  assign _GEN_106 = {{37{_GEN_38[15]}},_GEN_38}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@687.4]
  assign _T_1398 = $signed(_T_1397) + $signed(_GEN_106); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@687.4]
  assign _GEN_107 = {{38{_GEN_39[15]}},_GEN_39}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@688.4]
  assign _T_1399 = $signed(_T_1398) + $signed(_GEN_107); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@688.4]
  assign _GEN_108 = {{39{_GEN_40[15]}},_GEN_40}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@689.4]
  assign _T_1400 = $signed(_T_1399) + $signed(_GEN_108); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@689.4]
  assign _GEN_109 = {{40{_GEN_41[15]}},_GEN_41}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@690.4]
  assign _T_1401 = $signed(_T_1400) + $signed(_GEN_109); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@690.4]
  assign _GEN_110 = {{41{_GEN_42[15]}},_GEN_42}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@691.4]
  assign _T_1402 = $signed(_T_1401) + $signed(_GEN_110); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@691.4]
  assign _GEN_111 = {{42{_GEN_43[15]}},_GEN_43}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@692.4]
  assign _T_1403 = $signed(_T_1402) + $signed(_GEN_111); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@692.4]
  assign _GEN_112 = {{43{_GEN_44[15]}},_GEN_44}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@693.4]
  assign _T_1404 = $signed(_T_1403) + $signed(_GEN_112); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@693.4]
  assign _GEN_113 = {{44{_GEN_45[15]}},_GEN_45}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@694.4]
  assign _T_1405 = $signed(_T_1404) + $signed(_GEN_113); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@694.4]
  assign _GEN_114 = {{45{_GEN_46[15]}},_GEN_46}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@695.4]
  assign _T_1406 = $signed(_T_1405) + $signed(_GEN_114); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@695.4]
  assign _GEN_115 = {{46{_GEN_47[15]}},_GEN_47}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@696.4]
  assign _T_1407 = $signed(_T_1406) + $signed(_GEN_115); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@696.4]
  assign _GEN_116 = {{47{_GEN_48[15]}},_GEN_48}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@697.4]
  assign _T_1408 = $signed(_T_1407) + $signed(_GEN_116); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@697.4]
  assign _GEN_117 = {{48{_GEN_49[15]}},_GEN_49}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@698.4]
  assign _T_1409 = $signed(_T_1408) + $signed(_GEN_117); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@698.4]
  assign _GEN_118 = {{49{_GEN_50[15]}},_GEN_50}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@699.4]
  assign _T_1410 = $signed(_T_1409) + $signed(_GEN_118); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@699.4]
  assign _GEN_119 = {{50{_GEN_51[15]}},_GEN_51}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@700.4]
  assign _T_1411 = $signed(_T_1410) + $signed(_GEN_119); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@700.4]
  assign _GEN_120 = {{51{_GEN_52[15]}},_GEN_52}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@701.4]
  assign _T_1412 = $signed(_T_1411) + $signed(_GEN_120); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@701.4]
  assign _GEN_121 = {{52{_GEN_53[15]}},_GEN_53}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@702.4]
  assign _T_1413 = $signed(_T_1412) + $signed(_GEN_121); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@702.4]
  assign _GEN_122 = {{53{_GEN_54[15]}},_GEN_54}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@703.4]
  assign _T_1414 = $signed(_T_1413) + $signed(_GEN_122); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@703.4]
  assign _GEN_123 = {{54{_GEN_55[15]}},_GEN_55}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@704.4]
  assign _T_1415 = $signed(_T_1414) + $signed(_GEN_123); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@704.4]
  assign _GEN_124 = {{55{_GEN_56[15]}},_GEN_56}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@705.4]
  assign _T_1416 = $signed(_T_1415) + $signed(_GEN_124); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@705.4]
  assign _GEN_125 = {{56{_GEN_57[15]}},_GEN_57}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@706.4]
  assign _T_1417 = $signed(_T_1416) + $signed(_GEN_125); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@706.4]
  assign _GEN_126 = {{57{_GEN_58[15]}},_GEN_58}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@707.4]
  assign _T_1418 = $signed(_T_1417) + $signed(_GEN_126); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@707.4]
  assign _GEN_127 = {{58{_GEN_59[15]}},_GEN_59}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@708.4]
  assign _T_1419 = $signed(_T_1418) + $signed(_GEN_127); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@708.4]
  assign _GEN_128 = {{59{_GEN_60[15]}},_GEN_60}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@709.4]
  assign _T_1420 = $signed(_T_1419) + $signed(_GEN_128); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@709.4]
  assign _GEN_129 = {{60{_GEN_61[15]}},_GEN_61}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@710.4]
  assign _T_1421 = $signed(_T_1420) + $signed(_GEN_129); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@710.4]
  assign _GEN_130 = {{61{_GEN_62[15]}},_GEN_62}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@711.4]
  assign _T_1422 = $signed(_T_1421) + $signed(_GEN_130); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@711.4]
  assign _GEN_131 = {{62{_GEN_63[15]}},_GEN_63}; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@712.4]
  assign _T_1423 = $signed(_T_1422) + $signed(_GEN_131); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:32:@712.4]
  assign _T_1424 = $unsigned(_T_1423); // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 56:37:@713.4]
  assign _T_1425 = io_dat_actv_0_valid & io_wt_actv_0_valid; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 59:42:@714.4]
  assign io_mac_out_valid = _T_1437; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 62:22:@740.4]
  assign io_mac_out_bits = _T_1431[21:0]; // @[NV_NVDLA_CMAC_CORE_mac_dft.scala 61:21:@727.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  _T_1427 = _RAND_0[78:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  _T_1429 = _RAND_1[78:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {3{`RANDOM}};
  _T_1431 = _RAND_2[78:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1433 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1435 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1437 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (_T_1425) begin
      _T_1427 <= _T_1424;
    end
    if (_T_1425) begin
      _T_1429 <= _T_1427;
    end
    if (_T_1425) begin
      _T_1431 <= _T_1429;
    end
    if (_T_1425) begin
      _T_1433 <= _T_1425;
    end
    if (_T_1425) begin
      _T_1435 <= _T_1433;
    end
    if (_T_1425) begin
      _T_1437 <= _T_1435;
    end
  end
endmodule
